* NGSPICE file created from tt_um_jimktrains_vslc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt tt_um_jimktrains_vslc VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XTAP_TAPCELL_ROW_77_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1444__138 _1313__7/A VGND VGND VPWR VPWR _1596_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ _1459_/Q _1280_/B VGND VGND VPWR VPWR _1270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0985_ hold7/X _0987_/A _0984_/Y VGND VGND VPWR VPWR _1543_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1468_ _1468_/CLK _1468_/D VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
X_1537_ _1537_/CLK _1537_/D VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ _1550_/Q _1588_/Q VGND VGND VPWR VPWR _0770_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1253_ _1287_/A1 _1252_/X _1251_/X _1287_/C1 VGND VGND VPWR VPWR _1253_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1184_ _1487_/Q _1131_/C _1123_/Y _1174_/X VGND VGND VPWR VPWR _1184_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_19_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0968_ hold23/A _0993_/A VGND VGND VPWR VPWR _0991_/A sky130_fd_sc_hd__and2_1
Xclkbuf_4_12_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1313__7/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0899_ _0899_/A1 _1571_/Q _0889_/Y _0889_/B _1063_/A1 VGND VGND VPWR VPWR _0900_/B
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_58_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0822_ _0867_/A _0822_/B VGND VGND VPWR VPWR _1590_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1236_ hold35/A _0864_/Y _1246_/B1 _1235_/X VGND VGND VPWR VPWR _1236_/X sky130_fd_sc_hd__o211a_1
X_1305_ _1459_/Q _1458_/Q _1457_/Q _1471_/Q hold43/A _1489_/Q VGND VGND VPWR VPWR
+ _1306_/B sky130_fd_sc_hd__mux4_1
X_1098_ _1525_/Q _1096_/X _1098_/S VGND VGND VPWR VPWR _1098_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1167_ _1523_/Q _1109_/A _1165_/X _1166_/X VGND VGND VPWR VPWR _1182_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ _1018_/A _1138_/A _1020_/X _1294_/A VGND VGND VPWR VPWR _1529_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0805_ _0867_/A _0805_/B VGND VGND VPWR VPWR _1598_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0736_ _0736_/A VGND VGND VPWR VPWR _1069_/B sky130_fd_sc_hd__inv_2
X_1219_ _1082_/B _1020_/A _1007_/A VGND VGND VPWR VPWR _1219_/X sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1570_ _1570_/CLK _1570_/D VGND VGND VPWR VPWR _1570_/Q sky130_fd_sc_hd__dfxtp_1
X_1004_ hold27/A _1004_/B VGND VGND VPWR VPWR _1533_/D sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_32_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ _1484_/CLK _1484_/D VGND VGND VPWR VPWR _1484_/Q sky130_fd_sc_hd__dfxtp_1
X_1553_ _1553_/CLK _1553_/D VGND VGND VPWR VPWR _1553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1375__69 _1483_/CLK VGND VGND VPWR VPWR _1527_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0984_ hold7/X _0987_/A _1004_/B VGND VGND VPWR VPWR _0984_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1536_ _1536_/CLK _1536_/D VGND VGND VPWR VPWR _1536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1467_ _1467_/CLK _1467_/D VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1411__105 clkload5/A VGND VGND VPWR VPWR _1563_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1252_ hold42/A _1463_/Q _1252_/S VGND VGND VPWR VPWR _1252_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1183_ _1072_/A _1182_/X _1168_/A VGND VGND VPWR VPWR _1183_/Y sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_19_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0967_ hold11/A _1538_/Q hold10/A _0967_/D VGND VGND VPWR VPWR _0993_/A sky130_fd_sc_hd__and4_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1519_ _1519_/CLK _1519_/D VGND VGND VPWR VPWR _1519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ _1105_/A _0898_/B VGND VGND VPWR VPWR _1572_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1345__39 clkload1/A VGND VGND VPWR VPWR _1497_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0821_ _0912_/A1 _1590_/Q _0813_/Y _0813_/B _1291_/D VGND VGND VPWR VPWR _0822_/B
+ sky130_fd_sc_hd__a32o_1
X_0752_ _1600_/Q VGND VGND VPWR VPWR _0752_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ hold40/A _1280_/B VGND VGND VPWR VPWR _1235_/X sky130_fd_sc_hd__or2_1
X_1304_ _1463_/Q _1462_/Q _1461_/Q _1460_/Q hold43/A _1489_/Q VGND VGND VPWR VPWR
+ _1304_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1166_ hold15/A hold21/A hold31/A hold24/A VGND VGND VPWR VPWR _1166_/X sky130_fd_sc_hd__or4_1
XFILLER_0_74_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1097_ uo_out[5] _1097_/B VGND VGND VPWR VPWR _1097_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1417__111 clkload3/A VGND VGND VPWR VPWR _1569_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_11_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1312__6/A sky130_fd_sc_hd__clkbuf_8
X_1020_ _1020_/A _1030_/B VGND VGND VPWR VPWR _1020_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0735_ _1075_/A VGND VGND VPWR VPWR _1072_/A sky130_fd_sc_hd__inv_2
X_0804_ _0912_/A1 _1598_/Q _0792_/Y _0792_/A _1291_/D VGND VGND VPWR VPWR _0805_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1218_ _1082_/B _1528_/Q _1007_/A VGND VGND VPWR VPWR _1218_/Y sky130_fd_sc_hd__a21oi_2
X_1149_ _1149_/A _1149_/B VGND VGND VPWR VPWR _1149_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_58_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ hold27/X _1534_/Q _1002_/Y VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1552_ _1552_/CLK hold13/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1483_ _1483_/CLK input9/X VGND VGND VPWR VPWR _1483_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ _0972_/B _0995_/B _0983_/C VGND VGND VPWR VPWR _1544_/D sky130_fd_sc_hd__and3b_1
X_1535_ _1535_/CLK _1535_/D VGND VGND VPWR VPWR _1535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1466_ _1466_/CLK _1466_/D VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1450__144 clkload6/A VGND VGND VPWR VPWR _1602_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1251_ hold42/A _0864_/Y _1285_/C1 _1250_/X VGND VGND VPWR VPWR _1251_/X sky130_fd_sc_hd__o211a_1
X_1182_ _1182_/A _1182_/B _1182_/C VGND VGND VPWR VPWR _1182_/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0966_ hold11/A _1538_/Q _0967_/D VGND VGND VPWR VPWR _0966_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0897_ _0899_/A1 _1572_/Q _0889_/Y _0889_/B _1207_/A VGND VGND VPWR VPWR _0898_/B
+ sky130_fd_sc_hd__a32o_1
X_1434__128 clkload12/A VGND VGND VPWR VPWR _1586_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1518_ _1518_/CLK _1518_/D VGND VGND VPWR VPWR _1518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0751_ _1597_/Q VGND VGND VPWR VPWR _0751_/Y sky130_fd_sc_hd__inv_2
X_0820_ hold46/X _0801_/X _0813_/Y _0813_/B _0800_/A VGND VGND VPWR VPWR _1591_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1303_ _1292_/B _1301_/Y _1302_/X _1294_/A VGND VGND VPWR VPWR _1452_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1234_ hold35/X _1288_/A2 _1233_/X _1009_/A VGND VGND VPWR VPWR _1468_/D sky130_fd_sc_hd__o211a_1
X_1096_ _1292_/B uo_out[5] _1096_/S VGND VGND VPWR VPWR _1096_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1165_ hold17/A hold37/A _1496_/Q hold25/A VGND VGND VPWR VPWR _1165_/X sky130_fd_sc_hd__or4_1
XFILLER_0_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0949_ _0946_/X _0949_/B _0953_/C VGND VGND VPWR VPWR _1556_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1405__99 clkload7/A VGND VGND VPWR VPWR _1557_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0734_ _1169_/B VGND VGND VPWR VPWR _1024_/A sky130_fd_sc_hd__inv_2
X_0803_ hold26/X _0792_/Y _0801_/X _0800_/A _0792_/A VGND VGND VPWR VPWR _1599_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1079_ _1074_/X _1076_/X _1078_/X _1100_/A VGND VGND VPWR VPWR _1207_/B sky130_fd_sc_hd__o22ai_1
X_1217_ _1471_/Q _1005_/Y _1214_/X _1216_/X _1307_/C1 VGND VGND VPWR VPWR _1471_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1148_ hold45/A hold47/A hold50/A _1512_/Q VGND VGND VPWR VPWR _1149_/B sky130_fd_sc_hd__or4_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_58_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1002_ hold27/A _1534_/Q _1004_/B VGND VGND VPWR VPWR _1002_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1315__9/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1482_ _1482_/CLK input8/X VGND VGND VPWR VPWR _1482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1551_ _1551_/CLK _1551_/D VGND VGND VPWR VPWR _1551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ hold30/A hold7/A _0989_/A _1544_/Q VGND VGND VPWR VPWR _0983_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_73_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1465_ _1465_/CLK _1465_/D VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfxtp_1
X_1534_ _1534_/CLK hold28/X VGND VGND VPWR VPWR _1534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380__74 _1312__6/A VGND VGND VPWR VPWR _1532_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1250_ _1463_/Q _1280_/B VGND VGND VPWR VPWR _1250_/X sky130_fd_sc_hd__or2_1
X_1181_ hold36/X _1126_/B _1180_/X _0867_/A VGND VGND VPWR VPWR _1485_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_62_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0965_ hold27/A _1534_/Q _1535_/Q _1536_/Q VGND VGND VPWR VPWR _0967_/D sky130_fd_sc_hd__and4_1
X_0896_ hold14/X _0801_/X _0889_/Y _0889_/B _0800_/A VGND VGND VPWR VPWR _1573_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1517_ _1517_/CLK _1517_/D VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_36_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0750_ _1593_/Q VGND VGND VPWR VPWR _0750_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1302_ _1301_/A _1301_/B uo_out[0] VGND VGND VPWR VPWR _1302_/X sky130_fd_sc_hd__a21o_1
X_1233_ _1098_/S _1232_/X _1231_/X _1219_/X VGND VGND VPWR VPWR _1233_/X sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_63_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1095_ _1100_/A _1298_/A VGND VGND VPWR VPWR _1096_/S sky130_fd_sc_hd__nand2_1
X_1164_ _1523_/Q _1109_/A _1153_/Y _1162_/X _1163_/X VGND VGND VPWR VPWR _1182_/A
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_72_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0948_ _1556_/Q _0951_/A VGND VGND VPWR VPWR _0949_/B sky130_fd_sc_hd__or2_1
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0879_ _0899_/A1 _1580_/Q _0871_/Y _0871_/B _1207_/A VGND VGND VPWR VPWR _0880_/B
+ sky130_fd_sc_hd__a32o_1
X_1350__44 clkload0/A VGND VGND VPWR VPWR _1502_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0802_ _0867_/A _1196_/B VGND VGND VPWR VPWR _0974_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0733_ _1553_/Q VGND VGND VPWR VPWR _0733_/Y sky130_fd_sc_hd__inv_2
X_1216_ _1285_/C1 _1215_/X _1007_/A VGND VGND VPWR VPWR _1216_/X sky130_fd_sc_hd__a21o_1
X_1078_ uo_out[3] _1069_/Y _1295_/A uo_out[2] _1077_/X VGND VGND VPWR VPWR _1078_/X
+ sky130_fd_sc_hd__a221o_1
X_1147_ hold54/A hold48/A _1509_/Q hold53/A VGND VGND VPWR VPWR _1149_/A sky130_fd_sc_hd__or4_1
XFILLER_0_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1001_ _1001_/A _1004_/B _1001_/C VGND VGND VPWR VPWR _1535_/D sky130_fd_sc_hd__and3_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1320__14 clkload8/A VGND VGND VPWR VPWR _1463_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_57_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1407__101 clkload5/A VGND VGND VPWR VPWR _1559_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1481_ _1482_/CLK input7/X VGND VGND VPWR VPWR _1481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1386__80 _1482_/CLK VGND VGND VPWR VPWR _1538_/CLK sky130_fd_sc_hd__inv_2
X_1550_ _1550_/CLK _1550_/D VGND VGND VPWR VPWR _1550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ _0981_/A _0981_/B VGND VGND VPWR VPWR _1545_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1602_ _1602_/CLK _1602_/D VGND VGND VPWR VPWR _1602_/Q sky130_fd_sc_hd__dfxtp_1
X_1464_ _1464_/CLK _1464_/D VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
X_1533_ _1533_/CLK _1533_/D VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1356__50 clkload2/A VGND VGND VPWR VPWR _1508_/CLK sky130_fd_sc_hd__inv_2
X_1180_ _1301_/A _1168_/X _1180_/A3 _1179_/X VGND VGND VPWR VPWR _1180_/X sky130_fd_sc_hd__a31o_1
X_0964_ hold27/A _1534_/Q _1535_/Q VGND VGND VPWR VPWR _1001_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_54_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1516_ _1516_/CLK _1516_/D VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_1
X_0895_ _1105_/A _0895_/B VGND VGND VPWR VPWR _1574_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1301_ _1301_/A _1301_/B VGND VGND VPWR VPWR _1301_/Y sky130_fd_sc_hd__nand2_1
X_1232_ hold33/A hold41/A _1282_/S VGND VGND VPWR VPWR _1232_/X sky130_fd_sc_hd__mux2_1
X_1094_ uo_out[6] _1097_/B _1092_/X _1093_/X _1009_/A VGND VGND VPWR VPWR _1505_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1163_ hold21/A hold44/A VGND VGND VPWR VPWR _1163_/X sky130_fd_sc_hd__and2b_1
X_1440__134 _1313__7/A VGND VGND VPWR VPWR _1592_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0947_ _1557_/Q _0946_/X _0953_/C _0920_/Y VGND VGND VPWR VPWR _1557_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0878_ hold20/X _0801_/X _0871_/Y _0871_/B _0800_/A VGND VGND VPWR VPWR _1581_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_7_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clkload0/A VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_12
X_1326__20 _1315__9/A VGND VGND VPWR VPWR _1469_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1424__118 clkload1/A VGND VGND VPWR VPWR _1576_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0801_ _0893_/A _0801_/B VGND VGND VPWR VPWR _0801_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0732_ _1556_/Q VGND VGND VPWR VPWR _0732_/Y sky130_fd_sc_hd__inv_2
X_1215_ _1291_/D _1169_/B _1525_/Q _1075_/B _1471_/Q _1457_/Q VGND VGND VPWR VPWR
+ _1215_/X sky130_fd_sc_hd__mux4_1
X_1146_ hold43/X _1139_/B _1145_/Y VGND VGND VPWR VPWR _1488_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1077_ uo_out[1] _1298_/A _1301_/A uo_out[0] VGND VGND VPWR VPWR _1077_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ hold27/A _1534_/Q _1535_/Q VGND VGND VPWR VPWR _1001_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1446__140 _1313__7/A VGND VGND VPWR VPWR _1598_/CLK sky130_fd_sc_hd__inv_2
X_1129_ hold36/X _1492_/Q _1130_/S VGND VGND VPWR VPWR _1492_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1480_ _1482_/CLK input6/X VGND VGND VPWR VPWR _1480_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0980_ hold29/X _0972_/B _0995_/B VGND VGND VPWR VPWR _0981_/B sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_74_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1532_ _1532_/CLK _1532_/D VGND VGND VPWR VPWR _1532_/Q sky130_fd_sc_hd__dfxtp_1
X_1601_ _1601_/CLK _1601_/D VGND VGND VPWR VPWR _1601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1463_ _1463_/CLK _1463_/D VGND VGND VPWR VPWR _1463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1371__65 clkload0/A VGND VGND VPWR VPWR _1523_/CLK sky130_fd_sc_hd__inv_2
X_0963_ _0960_/B _0963_/B _0963_/C VGND VGND VPWR VPWR _1549_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0894_ _0801_/B _1574_/Q _0889_/Y _0889_/B _1289_/A VGND VGND VPWR VPWR _0895_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1515_ _1515_/CLK _1515_/D VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1300_ _1292_/B _1298_/Y _1299_/X _1294_/A VGND VGND VPWR VPWR _1453_/D sky130_fd_sc_hd__o211a_1
X_1231_ hold33/A _0864_/Y _1246_/B1 _1230_/X VGND VGND VPWR VPWR _1231_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1162_ _1521_/Q _1112_/A _1160_/X _1161_/X VGND VGND VPWR VPWR _1162_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1093_ _1100_/A _1246_/B1 _1087_/Y VGND VGND VPWR VPWR _1093_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_59_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0946_ _1556_/Q hold51/A _0946_/C VGND VGND VPWR VPWR _0946_/X sky130_fd_sc_hd__and3_1
X_0877_ _0886_/A _0877_/B VGND VGND VPWR VPWR _1582_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clkload1/A VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_21_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1341__35 clkload3/A VGND VGND VPWR VPWR _1493_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0800_ _0800_/A VGND VGND VPWR VPWR _1289_/B sky130_fd_sc_hd__inv_2
X_0731_ _1557_/Q VGND VGND VPWR VPWR _0731_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1214_ _1457_/Q _1252_/S _1287_/A1 _1213_/X VGND VGND VPWR VPWR _1214_/X sky130_fd_sc_hd__o211a_1
X_1145_ _1145_/A _1145_/B VGND VGND VPWR VPWR _1145_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1076_ uo_out[6] _1295_/A _1301_/A uo_out[4] _1024_/A VGND VGND VPWR VPWR _1076_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0929_ _1564_/Q _0931_/B VGND VGND VPWR VPWR _0932_/A sky130_fd_sc_hd__or2_1
XFILLER_0_30_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_69_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1128_ _1486_/Q hold4/X _1130_/S VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__mux2_1
X_1059_ _1020_/A _1051_/X _1058_/X _1063_/C1 VGND VGND VPWR VPWR _1512_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1377__71 _1483_/CLK VGND VGND VPWR VPWR _1529_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1531_ _1531_/CLK _1531_/D VGND VGND VPWR VPWR _1531_/Q sky130_fd_sc_hd__dfxtp_1
X_1462_ _1462_/CLK _1462_/D VGND VGND VPWR VPWR _1462_/Q sky130_fd_sc_hd__dfxtp_1
X_1600_ _1600_/CLK _1600_/D VGND VGND VPWR VPWR _1600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0962_ _1549_/Q _0974_/A VGND VGND VPWR VPWR _0963_/C sky130_fd_sc_hd__or2_1
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0893_ _0893_/A _0893_/B VGND VGND VPWR VPWR _1575_/D sky130_fd_sc_hd__and2_1
X_1514_ _1514_/CLK _1514_/D VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1347__41 clkload0/A VGND VGND VPWR VPWR _1499_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1309__3 _1312__6/A VGND VGND VPWR VPWR _1452_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout60 _1196_/A VGND VGND VPWR VPWR _1294_/A sky130_fd_sc_hd__buf_2
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1092_ _1292_/B _1090_/Y _1091_/X _1098_/S VGND VGND VPWR VPWR _1092_/X sky130_fd_sc_hd__o211a_1
X_1230_ hold41/A _1245_/B VGND VGND VPWR VPWR _1230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1161_ _1521_/Q _1112_/A _0739_/Y _1520_/Q VGND VGND VPWR VPWR _1161_/X sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_32_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0876_ _0899_/A1 _1582_/Q _0871_/Y _0871_/B _1289_/A VGND VGND VPWR VPWR _0877_/B
+ sky130_fd_sc_hd__a32o_1
X_0945_ hold51/A _0946_/C VGND VGND VPWR VPWR _0951_/A sky130_fd_sc_hd__and2_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clkload2/A VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_12
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0730_ _1558_/Q VGND VGND VPWR VPWR _0730_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1213_ _1207_/Y _1210_/X _1212_/X _1291_/C VGND VGND VPWR VPWR _1213_/X sky130_fd_sc_hd__a31o_1
X_1317__11 clkload8/A VGND VGND VPWR VPWR _1460_/CLK sky130_fd_sc_hd__inv_2
X_1075_ _1075_/A _1075_/B VGND VGND VPWR VPWR _1301_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1144_ _1144_/A _1144_/B VGND VGND VPWR VPWR _1489_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0859_ _1016_/A _1071_/B _0906_/C VGND VGND VPWR VPWR _0859_/X sky130_fd_sc_hd__or3_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ _1563_/Q hold49/A _0928_/C VGND VGND VPWR VPWR _0931_/B sky130_fd_sc_hd__and3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1401__95 clkload7/A VGND VGND VPWR VPWR _1553_/CLK sky130_fd_sc_hd__inv_2
X_1430__124 clkload4/A VGND VGND VPWR VPWR _1582_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1127_ _1178_/A hold3/X _1130_/S VGND VGND VPWR VPWR _1494_/D sky130_fd_sc_hd__mux2_1
X_1058_ _1512_/Q _1066_/B VGND VGND VPWR VPWR _1058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1414__108 _1483_/CLK VGND VGND VPWR VPWR _1566_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1392__86 _1482_/CLK VGND VGND VPWR VPWR _1544_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1530_ _1530_/CLK _1530_/D VGND VGND VPWR VPWR _1530_/Q sky130_fd_sc_hd__dfxtp_1
X_1436__130 clkload9/A VGND VGND VPWR VPWR _1588_/CLK sky130_fd_sc_hd__inv_2
X_1461_ _1461_/CLK _1461_/D VGND VGND VPWR VPWR _1461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0961_ _0958_/B _0961_/B _0963_/B VGND VGND VPWR VPWR _1550_/D sky130_fd_sc_hd__and3b_1
X_0892_ _0899_/A1 _1575_/Q _0889_/Y _0889_/B _1016_/A VGND VGND VPWR VPWR _0893_/B
+ sky130_fd_sc_hd__a32o_1
X_1513_ _1513_/CLK _1513_/D VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfxtp_1
X_1362__56 clkload2/A VGND VGND VPWR VPWR _1514_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout61 _1196_/A VGND VGND VPWR VPWR _0915_/A sky130_fd_sc_hd__buf_1
Xfanout50 _1487_/Q VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1091_ _1100_/A _1295_/A uo_out[6] VGND VGND VPWR VPWR _1091_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1160_ _1157_/X _1158_/X _1159_/X VGND VGND VPWR VPWR _1160_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0944_ _1554_/Q _0960_/B _0944_/C VGND VGND VPWR VPWR _0946_/C sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_15_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0886_/A _0875_/B VGND VGND VPWR VPWR _1583_/D sky130_fd_sc_hd__and2_1
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1311__5 _1312__6/A VGND VGND VPWR VPWR _1454_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_65_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1289_ _1289_/A _1289_/B _1289_/C _1289_/D VGND VGND VPWR VPWR _1290_/S sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload3 clkload3/A VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_12
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1212_ _1477_/Q _1298_/A _1206_/X _1211_/X VGND VGND VPWR VPWR _1212_/X sky130_fd_sc_hd__a211o_1
X_1332__26 clkload9/A VGND VGND VPWR VPWR _1484_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1074_ uo_out[7] _1069_/Y _1298_/A uo_out[5] VGND VGND VPWR VPWR _1074_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1143_ _1489_/Q _1145_/B _1068_/A VGND VGND VPWR VPWR _1144_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ hold49/X _0928_/C VGND VGND VPWR VPWR _0927_/Y sky130_fd_sc_hd__nand2_1
X_0858_ _1071_/A _1082_/B _0906_/C VGND VGND VPWR VPWR _1291_/C sky130_fd_sc_hd__nor3_2
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0789_ hold39/A _0789_/B _0789_/C _0789_/D VGND VGND VPWR VPWR _0789_/X sky130_fd_sc_hd__and4_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1398__92 clkload12/A VGND VGND VPWR VPWR _1550_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1126_ _1145_/A _1126_/B VGND VGND VPWR VPWR _1130_/S sky130_fd_sc_hd__nand2_1
X_1057_ _1289_/A _1051_/X _1056_/X _1063_/C1 VGND VGND VPWR VPWR _1513_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _1109_/A _1111_/A VGND VGND VPWR VPWR _1502_/D sky130_fd_sc_hd__xnor2_1
X_1368__62 clkload3/A VGND VGND VPWR VPWR _1520_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ _1460_/CLK _1460_/D VGND VGND VPWR VPWR _1460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1589_ _1589_/CLK _1589_/D VGND VGND VPWR VPWR _1589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ _1550_/Q _0960_/B VGND VGND VPWR VPWR _0961_/B sky130_fd_sc_hd__or2_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1512_ _1512_/CLK _1512_/D VGND VGND VPWR VPWR _1512_/Q sky130_fd_sc_hd__dfxtp_1
X_0891_ _1105_/A _0891_/B VGND VGND VPWR VPWR _1576_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1338__32 clkload2/A VGND VGND VPWR VPWR _1490_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_76_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout62 input1/X VGND VGND VPWR VPWR _1196_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout40 _1529_/Q VGND VGND VPWR VPWR _1289_/A sky130_fd_sc_hd__buf_2
Xfanout51 _1145_/A VGND VGND VPWR VPWR _1063_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ _1100_/A _1295_/A VGND VGND VPWR VPWR _1090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload10 _1312__6/A VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_8
X_0943_ _0960_/B _0944_/C VGND VGND VPWR VPWR _0952_/B sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_15_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0874_ _0899_/A1 _1583_/Q _0871_/Y _0871_/B _1016_/A VGND VGND VPWR VPWR _0875_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1288_ _1457_/Q _1288_/A2 _1287_/X _1288_/C1 VGND VGND VPWR VPWR _1457_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_38_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload4 clkload4/A VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_12
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ _1478_/Q _1295_/A _1207_/A _1169_/B VGND VGND VPWR VPWR _1211_/X sky130_fd_sc_hd__a211o_1
X_1142_ _1490_/Q _1144_/A _1141_/Y VGND VGND VPWR VPWR _1490_/D sky130_fd_sc_hd__a21o_1
X_1073_ _1525_/Q _1075_/B VGND VGND VPWR VPWR _1298_/A sky130_fd_sc_hd__and2b_2
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0857_ _1018_/A _1020_/A VGND VGND VPWR VPWR _0906_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ _0928_/C VGND VGND VPWR VPWR _0926_/Y sky130_fd_sc_hd__inv_2
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0788_ _1553_/Q _0749_/Y _0751_/Y _1559_/Q _0773_/X VGND VGND VPWR VPWR _0790_/C
+ sky130_fd_sc_hd__a221o_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ _1126_/B VGND VGND VPWR VPWR _1125_/Y sky130_fd_sc_hd__inv_2
X_1056_ hold50/X _1066_/B VGND VGND VPWR VPWR _1056_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0909_ _1294_/A _0909_/B VGND VGND VPWR VPWR _1568_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1039_ _1289_/A _1033_/X _1038_/X _1063_/C1 VGND VGND VPWR VPWR _1521_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ hold21/A hold31/A _1114_/A VGND VGND VPWR VPWR _1111_/A sky130_fd_sc_hd__and3_1
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1420__114 clkload4/A VGND VGND VPWR VPWR _1572_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1383__77 clkload12/A VGND VGND VPWR VPWR _1535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_66_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1588_ _1588_/CLK _1588_/D VGND VGND VPWR VPWR _1588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0899_/A1 _1576_/Q _0889_/Y _0889_/B _1071_/B VGND VGND VPWR VPWR _0891_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1511_ _1511_/CLK _1511_/D VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1353__47 _1315__9/A VGND VGND VPWR VPWR _1505_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout41 _1528_/Q VGND VGND VPWR VPWR _1020_/A sky130_fd_sc_hd__buf_2
Xfanout30 _1245_/B VGND VGND VPWR VPWR _1280_/B sky130_fd_sc_hd__clkbuf_2
Xfanout52 _0886_/A VGND VGND VPWR VPWR _1105_/A sky130_fd_sc_hd__clkbuf_2
X_1426__120 clkload5/A VGND VGND VPWR VPWR _1578_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload11 _1313__7/A VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_8
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0942_ _1551_/Q _1550_/Q _0960_/B VGND VGND VPWR VPWR _0942_/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_15_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0873_ _0886_/A _0873_/B VGND VGND VPWR VPWR _1584_/D sky130_fd_sc_hd__and2_1
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1287_ _1287_/A1 _1286_/X _1285_/X _1287_/C1 VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_38_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload5 clkload5/A VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_8
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ _1483_/Q _1069_/Y _1208_/X _1209_/X VGND VGND VPWR VPWR _1210_/X sky130_fd_sc_hd__a211o_1
X_1072_ _1072_/A _1075_/B VGND VGND VPWR VPWR _1295_/A sky130_fd_sc_hd__nor2_2
X_1141_ _1490_/Q _1144_/A _1145_/A VGND VGND VPWR VPWR _1141_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0856_ _1071_/A _1082_/B _1471_/Q _1018_/A VGND VGND VPWR VPWR _0856_/X sky130_fd_sc_hd__or4b_1
X_0787_ _0769_/X _0770_/Y _0771_/X _0772_/Y _0768_/X VGND VGND VPWR VPWR _0790_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0925_ _1561_/Q _1560_/Q _1559_/Q _0925_/D VGND VGND VPWR VPWR _0928_/C sky130_fd_sc_hd__and4_1
X_1323__17 _1315__9/A VGND VGND VPWR VPWR _1466_/CLK sky130_fd_sc_hd__inv_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1389__83 _1482_/CLK VGND VGND VPWR VPWR _1541_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1124_ _1490_/Q _1489_/Q hold43/A _1123_/A VGND VGND VPWR VPWR _1126_/B sky130_fd_sc_hd__o31ai_4
X_1055_ _1016_/A _1051_/X _1054_/X _1063_/C1 VGND VGND VPWR VPWR _1514_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0908_ _1196_/B _1568_/Q _0907_/Y _0907_/B _1291_/D VGND VGND VPWR VPWR _0909_/B
+ sky130_fd_sc_hd__a32o_1
X_0839_ _0732_/Y _1576_/Q _1550_/Q _0744_/Y VGND VGND VPWR VPWR _0841_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1038_ _1521_/Q _1048_/B VGND VGND VPWR VPWR _1038_/X sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1107_ hold24/A _1116_/A VGND VGND VPWR VPWR _1114_/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1359__53 clkload3/A VGND VGND VPWR VPWR _1511_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1443__137 clkload6/A VGND VGND VPWR VPWR _1595_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_75_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1587_ _1587_/CLK _1587_/D VGND VGND VPWR VPWR _1587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1510_ _1510_/CLK _1510_/D VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout42 _1207_/A VGND VGND VPWR VPWR _1291_/D sky130_fd_sc_hd__buf_2
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout53 _0893_/A VGND VGND VPWR VPWR _0886_/A sky130_fd_sc_hd__clkbuf_2
Xfanout31 _0801_/B VGND VGND VPWR VPWR _0899_/A1 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1329__23 _1315__9/A VGND VGND VPWR VPWR _1472_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ _1550_/Q _0960_/B VGND VGND VPWR VPWR _0958_/B sky130_fd_sc_hd__and2_1
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload12 clkload12/A VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_8
XFILLER_0_42_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0872_ _0899_/A1 _1584_/Q _0871_/Y _0871_/B _1071_/B VGND VGND VPWR VPWR _0873_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1286_ _1471_/Q _1458_/Q _1291_/C VGND VGND VPWR VPWR _1286_/X sky130_fd_sc_hd__mux2_1
X_1449__143 clkload6/A VGND VGND VPWR VPWR _1601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload6 clkload6/A VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_8
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1071_ _1071_/A _1071_/B _1018_/A _1020_/A VGND VGND VPWR VPWR _1071_/X sky130_fd_sc_hd__or4bb_1
X_1140_ _1489_/Q _1145_/B VGND VGND VPWR VPWR _1144_/A sky130_fd_sc_hd__or2_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0924_ _0937_/A _0937_/B VGND VGND VPWR VPWR _0924_/Y sky130_fd_sc_hd__nor2_1
X_0786_ hold51/A _0750_/Y _0778_/X _0784_/X _0785_/Y VGND VGND VPWR VPWR _0790_/A
+ sky130_fd_sc_hd__a2111o_1
X_0855_ _0888_/A _1492_/Q _1491_/Q VGND VGND VPWR VPWR _1289_/C sky130_fd_sc_hd__or3b_2
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1269_ _1461_/Q _1288_/A2 _1268_/X _1307_/C1 VGND VGND VPWR VPWR _1461_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1123_ _1123_/A VGND VGND VPWR VPWR _1123_/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1054_ hold47/X _1066_/B VGND VGND VPWR VPWR _1054_/X sky130_fd_sc_hd__or2_1
X_0907_ _0907_/A _0907_/B VGND VGND VPWR VPWR _0907_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0769_ _1550_/Q _1588_/Q VGND VGND VPWR VPWR _0769_/X sky130_fd_sc_hd__or2_1
X_0838_ _1549_/Q _0743_/Y _0745_/Y _1551_/Q VGND VGND VPWR VPWR _0841_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_54_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1106_ hold17/A hold37/A _1117_/B VGND VGND VPWR VPWR _1116_/A sky130_fd_sc_hd__and3_1
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1037_ _1016_/A _1033_/X _1036_/X _1063_/C1 VGND VGND VPWR VPWR _1522_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1374__68 _1483_/CLK VGND VGND VPWR VPWR _1526_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1586_ _1586_/CLK _1586_/D VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1314__8 clkload8/A VGND VGND VPWR VPWR _1457_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1410__104 clkload5/A VGND VGND VPWR VPWR _1562_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1569_ _1569_/CLK _1569_/D VGND VGND VPWR VPWR _1569_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout21 _1105_/D VGND VGND VPWR VPWR _1138_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout43 _1527_/Q VGND VGND VPWR VPWR _1207_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout54 _1145_/A VGND VGND VPWR VPWR _0893_/A sky130_fd_sc_hd__clkbuf_2
Xfanout32 _1585_/Q VGND VGND VPWR VPWR _0801_/B sky130_fd_sc_hd__buf_2
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1344__38 clkload4/A VGND VGND VPWR VPWR _1496_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ _1558_/Q _0920_/A _0922_/Y _0963_/B VGND VGND VPWR VPWR _1558_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload13 _1483_/CLK VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_6
X_0871_ _0907_/A _0871_/B VGND VGND VPWR VPWR _0871_/Y sky130_fd_sc_hd__nor2_2
X_1285_ _1458_/Q _1285_/A2 _0867_/C _1285_/C1 VGND VGND VPWR VPWR _1285_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload7 clkload7/A VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_16
XTAP_TAPCELL_ROW_6_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _1075_/A _1075_/B VGND VGND VPWR VPWR _1292_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0854_ _0854_/A hold3/A hold4/A VGND VGND VPWR VPWR _0888_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0923_ _1559_/Q _0925_/D VGND VGND VPWR VPWR _0937_/B sky130_fd_sc_hd__nand2_1
X_1416__110 clkload12/A VGND VGND VPWR VPWR _1568_/CLK sky130_fd_sc_hd__inv_2
X_0785_ _0730_/Y _1596_/Q _0767_/Y _0776_/Y _0777_/Y VGND VGND VPWR VPWR _0785_/Y
+ sky130_fd_sc_hd__o2111ai_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ _1287_/A1 _1267_/X _1266_/X _1287_/C1 VGND VGND VPWR VPWR _1268_/X sky130_fd_sc_hd__a211o_1
X_1199_ _1490_/Q _1201_/A _1199_/C VGND VGND VPWR VPWR _1199_/Y sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ _1178_/A _1486_/Q _1122_/C VGND VGND VPWR VPWR _1123_/A sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_48_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1053_ _1071_/B _1051_/X _1052_/X _1063_/C1 VGND VGND VPWR VPWR _1515_/D sky130_fd_sc_hd__o211a_1
X_0906_ _1071_/B _1289_/C _0906_/C _1071_/A VGND VGND VPWR VPWR _0907_/B sky130_fd_sc_hd__and4bb_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0837_ _0729_/Y _1579_/Q _1580_/Q _0937_/A _0831_/X VGND VGND VPWR VPWR _0841_/A
+ sky130_fd_sc_hd__a221o_1
X_0768_ hold12/A _1590_/Q VGND VGND VPWR VPWR _0768_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ _1105_/A _1496_/Q hold25/A _1105_/D VGND VGND VPWR VPWR _1117_/B sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_51_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1036_ hold44/X _1048_/B VGND VGND VPWR VPWR _1036_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1585_ _1585_/CLK _1585_/D VGND VGND VPWR VPWR _1585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _1071_/A _1105_/D _1018_/X _0915_/A VGND VGND VPWR VPWR _1530_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1568_ _1568_/CLK _1568_/D VGND VGND VPWR VPWR _1568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1499_ _1499_/CLK _1499_/D VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
Xfanout44 _1169_/B VGND VGND VPWR VPWR _1100_/A sky130_fd_sc_hd__buf_2
XFILLER_0_68_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout22 _1015_/X VGND VGND VPWR VPWR _1105_/D sky130_fd_sc_hd__clkbuf_2
Xfanout33 _1585_/Q VGND VGND VPWR VPWR _0912_/A1 sky130_fd_sc_hd__buf_2
Xfanout55 input1/X VGND VGND VPWR VPWR _1145_/A sky130_fd_sc_hd__buf_2
Xfanout11 _0963_/B VGND VGND VPWR VPWR _0953_/C sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1433__127 clkload9/A VGND VGND VPWR VPWR _1585_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ _0888_/A _1033_/B VGND VGND VPWR VPWR _0871_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload14 _1482_/CLK VGND VGND VPWR VPWR clkload14/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1284_ _1458_/Q _1288_/A2 _1283_/X _1307_/C1 VGND VGND VPWR VPWR _1458_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_73_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ _0967_/D _1004_/B _0999_/C VGND VGND VPWR VPWR _1536_/D sky130_fd_sc_hd__and3b_1
Xclkload8 clkload8/A VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1404__98 clkload5/A VGND VGND VPWR VPWR _1556_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0753__1 _1315__9/A VGND VGND VPWR VPWR _1451_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0853_ hold39/X _0930_/B _0852_/Y VGND VGND VPWR VPWR _1586_/D sky130_fd_sc_hd__o21a_1
X_0922_ _0925_/D VGND VGND VPWR VPWR _0922_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0784_ _1549_/Q _0747_/Y _0765_/X _0774_/X _0775_/X VGND VGND VPWR VPWR _0784_/X
+ sky130_fd_sc_hd__a2111o_1
Xinput1 rst_n VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1267_ _1462_/Q _1460_/Q _1282_/S VGND VGND VPWR VPWR _1267_/X sky130_fd_sc_hd__mux2_1
X_1198_ _1512_/Q hold50/A hold47/A hold45/A hold43/A _1489_/Q VGND VGND VPWR VPWR
+ _1199_/C sky130_fd_sc_hd__mux4_1
XFILLER_0_61_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1439__133 clkload6/A VGND VGND VPWR VPWR _1591_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1121_ _1484_/Q hold36/A VGND VGND VPWR VPWR _1122_/C sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_48_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1052_ hold45/X _1066_/B VGND VGND VPWR VPWR _1052_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0905_ _1082_/B _1071_/A VGND VGND VPWR VPWR _1289_/D sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0767_ _1554_/Q _1592_/Q VGND VGND VPWR VPWR _0767_/Y sky130_fd_sc_hd__nand2b_1
X_0836_ _0733_/Y hold14/A _0829_/Y _0835_/X hold39/A VGND VGND VPWR VPWR _0850_/A
+ sky130_fd_sc_hd__a2111o_1
X_1395__89 _1482_/CLK VGND VGND VPWR VPWR _1547_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1104_ uo_out[4] _1097_/B _1103_/X _1288_/C1 VGND VGND VPWR VPWR _1503_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1035_ _1071_/B _1033_/X _1034_/X _1063_/C1 VGND VGND VPWR VPWR _1523_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_75_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0819_ _0867_/A _0819_/B VGND VGND VPWR VPWR _1592_/D sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_26_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1584_ _1584_/CLK _1584_/D VGND VGND VPWR VPWR _1584_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_53_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1365__59 clkload1/A VGND VGND VPWR VPWR _1517_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1018_ _1018_/A _1030_/B VGND VGND VPWR VPWR _1018_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_62_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_80_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1567_ _1567_/CLK _1567_/D VGND VGND VPWR VPWR _1567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1498_ _1498_/CLK _1498_/D VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout45 _1063_/A1 VGND VGND VPWR VPWR _1169_/B sky130_fd_sc_hd__buf_2
Xfanout56 _1288_/C1 VGND VGND VPWR VPWR _1307_/C1 sky130_fd_sc_hd__buf_2
Xfanout23 _1252_/S VGND VGND VPWR VPWR _1282_/S sky130_fd_sc_hd__clkbuf_4
Xfanout34 _1585_/Q VGND VGND VPWR VPWR _1196_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout12 _0930_/Y VGND VGND VPWR VPWR _0963_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1283_ _1287_/A1 _1282_/X _1281_/X _1287_/C1 VGND VGND VPWR VPWR _1283_/X sky130_fd_sc_hd__a211o_1
X_1335__29 clkload9/A VGND VGND VPWR VPWR _1487_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0998_ hold27/A _1534_/Q _1535_/Q _1536_/Q VGND VGND VPWR VPWR _0999_/C sky130_fd_sc_hd__a31o_1
Xclkload9 clkload9/A VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_16
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0753__2 _1315__9/A VGND VGND VPWR VPWR _1308_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0921_ _1558_/Q _0960_/B _0944_/C _0921_/D VGND VGND VPWR VPWR _0925_/D sky130_fd_sc_hd__and4_1
X_0852_ hold39/A _0930_/B _0974_/B VGND VGND VPWR VPWR _0852_/Y sky130_fd_sc_hd__a21oi_1
X_0783_ _0732_/Y _1594_/Q _1595_/Q _0731_/Y _0766_/X VGND VGND VPWR VPWR _0789_/D
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 ui_in[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
X_1266_ _1462_/Q _1285_/A2 _1285_/C1 _1265_/X VGND VGND VPWR VPWR _1266_/X sky130_fd_sc_hd__o211a_1
X_1197_ hold48/A hold54/A hold43/A VGND VGND VPWR VPWR _1201_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1051_ _1051_/A _1051_/B VGND VGND VPWR VPWR _1051_/X sky130_fd_sc_hd__or2_2
X_1120_ hold25/X _1120_/B VGND VGND VPWR VPWR _1495_/D sky130_fd_sc_hd__xnor2_1
X_0904_ _1145_/A _0904_/B VGND VGND VPWR VPWR _1569_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0766_ hold26/A _1561_/Q VGND VGND VPWR VPWR _0766_/X sky130_fd_sc_hd__and2b_1
X_0835_ _0727_/Y hold20/A _1582_/Q _0726_/Y _0834_/X VGND VGND VPWR VPWR _0835_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1249_ hold42/X _1218_/Y _1248_/X _1009_/A VGND VGND VPWR VPWR _1465_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap20 _1182_/C VGND VGND VPWR VPWR _1180_/A3 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_45_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1406__100 clkload7/A VGND VGND VPWR VPWR _1558_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1103_ _0736_/A _1246_/B1 _1087_/Y _1102_/X VGND VGND VPWR VPWR _1103_/X sky130_fd_sc_hd__a211o_1
X_1034_ _1523_/Q _1048_/B VGND VGND VPWR VPWR _1034_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0818_ _0912_/A1 _1592_/Q _0813_/Y _0813_/B _1018_/A VGND VGND VPWR VPWR _0819_/B
+ sky130_fd_sc_hd__a32o_1
X_0749_ hold46/A VGND VGND VPWR VPWR _0749_/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1583_ _1583_/CLK _1583_/D VGND VGND VPWR VPWR _1583_/Q sky130_fd_sc_hd__dfxtp_1
X_1017_ _1082_/B _1138_/A _1016_/X _1294_/A VGND VGND VPWR VPWR _1531_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_64_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1566_ _1566_/CLK _1566_/D VGND VGND VPWR VPWR _1566_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_18_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1497_ _1497_/CLK _1497_/D VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
Xfanout57 _1288_/C1 VGND VGND VPWR VPWR _1009_/A sky130_fd_sc_hd__buf_2
XFILLER_0_76_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout46 _1526_/Q VGND VGND VPWR VPWR _1063_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout35 _1071_/B VGND VGND VPWR VPWR _1082_/B sky130_fd_sc_hd__clkbuf_4
Xfanout24 _0859_/X VGND VGND VPWR VPWR _1252_/S sky130_fd_sc_hd__clkbuf_2
Xfanout13 _1219_/X VGND VGND VPWR VPWR _1287_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1282_ _1459_/Q _1457_/Q _1282_/S VGND VGND VPWR VPWR _1282_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1618_ _1618_/A VGND VGND VPWR VPWR uio_out[7] sky130_fd_sc_hd__clkbuf_4
X_0997_ hold11/X _0967_/D _0996_/Y VGND VGND VPWR VPWR _1537_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1549_ _1549_/CLK _1549_/D VGND VGND VPWR VPWR _1549_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0920_ _0920_/A VGND VGND VPWR VPWR _0920_/Y sky130_fd_sc_hd__inv_2
X_0851_ wire17/X _0850_/Y _0974_/A VGND VGND VPWR VPWR _0930_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0782_ _1549_/Q _0747_/Y _1594_/Q _0732_/Y _0781_/Y VGND VGND VPWR VPWR _0789_/C
+ sky130_fd_sc_hd__o221a_1
X_1265_ _1460_/Q _1280_/B VGND VGND VPWR VPWR _1265_/X sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 ui_in[1] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
X_1196_ _1196_/A _1196_/B _1196_/C VGND VGND VPWR VPWR _1473_/D sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1423__117 clkload4/A VGND VGND VPWR VPWR _1575_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1050_ _1051_/A _1051_/B VGND VGND VPWR VPWR _1066_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0903_ _1585_/Q _0743_/Y _0889_/Y _0889_/B _1069_/B VGND VGND VPWR VPWR _0904_/B
+ sky130_fd_sc_hd__a32o_1
X_0834_ _1564_/Q _1584_/Q VGND VGND VPWR VPWR _0834_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0765_ _1592_/Q _1554_/Q VGND VGND VPWR VPWR _0765_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1248_ _1098_/S _1247_/X _1246_/X _1219_/X VGND VGND VPWR VPWR _1248_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1179_ _1152_/A _1122_/C _1125_/Y _1150_/X _1178_/Y VGND VGND VPWR VPWR _1179_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1102_ _1292_/B _1100_/Y _1101_/X _1098_/S VGND VGND VPWR VPWR _1102_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_76_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1033_ _1051_/A _1033_/B VGND VGND VPWR VPWR _1033_/X sky130_fd_sc_hd__or2_2
X_0817_ _0867_/A _0817_/B VGND VGND VPWR VPWR _1593_/D sky130_fd_sc_hd__and2_1
XFILLER_0_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0748_ _1588_/Q VGND VGND VPWR VPWR _0748_/Y sky130_fd_sc_hd__inv_2
X_1429__123 clkload6/A VGND VGND VPWR VPWR _1581_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1582_ _1582_/CLK _1582_/D VGND VGND VPWR VPWR _1582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1016_ _1016_/A _1030_/B VGND VGND VPWR VPWR _1016_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1370__64 clkload0/A VGND VGND VPWR VPWR _1522_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1565_ _1565_/CLK _1565_/D VGND VGND VPWR VPWR _1565_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1496_ _1496_/CLK _1496_/D VGND VGND VPWR VPWR _1496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout58 input1/X VGND VGND VPWR VPWR _1288_/C1 sky130_fd_sc_hd__clkbuf_2
Xfanout47 _1525_/Q VGND VGND VPWR VPWR _1075_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout36 _1531_/Q VGND VGND VPWR VPWR _1071_/B sky130_fd_sc_hd__clkbuf_4
Xfanout25 _1082_/Y VGND VGND VPWR VPWR _1287_/A1 sky130_fd_sc_hd__buf_2
Xfanout14 _1218_/Y VGND VGND VPWR VPWR _1288_/A2 sky130_fd_sc_hd__buf_2
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ _1459_/Q _1285_/A2 _1285_/C1 _1280_/X VGND VGND VPWR VPWR _1281_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_58_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0996_ hold11/X _0967_/D _1004_/B VGND VGND VPWR VPWR _0996_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1617_ _1617_/A VGND VGND VPWR VPWR uio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ _1482_/CLK input5/X VGND VGND VPWR VPWR _1479_/Q sky130_fd_sc_hd__dfxtp_1
X_1548_ _1548_/CLK _1548_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_59_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1340__34 clkload9/A VGND VGND VPWR VPWR _1492_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0850_ _0850_/A _0850_/B _0850_/C VGND VGND VPWR VPWR _0850_/Y sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_11_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0781_ _1564_/Q _1602_/Q VGND VGND VPWR VPWR _0781_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 ui_in[2] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
X_1264_ _1462_/Q _1288_/A2 _1263_/X _1307_/C1 VGND VGND VPWR VPWR _1462_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1195_ _1618_/A _1194_/Y _1195_/S VGND VGND VPWR VPWR _1196_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0979_ hold6/X _0981_/A _0978_/Y VGND VGND VPWR VPWR _1546_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0833_ _1551_/Q _1571_/Q VGND VGND VPWR VPWR _0833_/X sky130_fd_sc_hd__and2b_1
X_0902_ _1105_/A _0902_/B VGND VGND VPWR VPWR _1570_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0764_ _0758_/X _0760_/X _0763_/X _1568_/Q VGND VGND VPWR VPWR _0974_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1247_ hold40/A hold34/A _1282_/S VGND VGND VPWR VPWR _1247_/X sky130_fd_sc_hd__mux2_1
X_1178_ _1178_/A _1486_/Q _1152_/B VGND VGND VPWR VPWR _1178_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ _1100_/A _1301_/A uo_out[4] VGND VGND VPWR VPWR _1101_/X sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_76_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1032_ _1051_/A _1033_/B VGND VGND VPWR VPWR _1048_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0747_ _1587_/Q VGND VGND VPWR VPWR _0747_/Y sky130_fd_sc_hd__inv_2
X_0816_ _0912_/A1 _1593_/Q _0813_/Y _0813_/B _1016_/A VGND VGND VPWR VPWR _0817_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376__70 clkload9/A VGND VGND VPWR VPWR _1528_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1581_ _1581_/CLK _1581_/D VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1015_ _1173_/B _1152_/A _1173_/A VGND VGND VPWR VPWR _1015_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1564_ _1564_/CLK _1564_/D VGND VGND VPWR VPWR _1564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1346__40 clkload1/A VGND VGND VPWR VPWR _1498_/CLK sky130_fd_sc_hd__inv_2
X_1495_ _1495_/CLK _1495_/D VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfxtp_1
Xfanout15 _1004_/B VGND VGND VPWR VPWR _0995_/B sky130_fd_sc_hd__clkbuf_2
Xfanout26 _1082_/Y VGND VGND VPWR VPWR _1098_/S sky130_fd_sc_hd__buf_2
Xfanout37 _1016_/A VGND VGND VPWR VPWR _1071_/A sky130_fd_sc_hd__buf_2
Xfanout48 _0736_/A VGND VGND VPWR VPWR _1075_/B sky130_fd_sc_hd__clkbuf_4
Xfanout59 _1196_/A VGND VGND VPWR VPWR _0867_/A sky130_fd_sc_hd__buf_2
XFILLER_0_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1280_ _1457_/Q _1280_/B VGND VGND VPWR VPWR _1280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ _0966_/X _0995_/B _0995_/C VGND VGND VPWR VPWR _1538_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1616_ hold2/A VGND VGND VPWR VPWR uio_out[2] sky130_fd_sc_hd__clkbuf_4
X_1547_ _1547_/CLK _1547_/D VGND VGND VPWR VPWR _1547_/Q sky130_fd_sc_hd__dfxtp_1
X_1478_ _1482_/CLK input4/X VGND VGND VPWR VPWR _1478_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ _0731_/Y _1595_/Q _0752_/Y hold49/A _0779_/Y VGND VGND VPWR VPWR _0789_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_11_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 ui_in[3] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
X_1194_ hold19/A wire17/X _1618_/A VGND VGND VPWR VPWR _1194_/Y sky130_fd_sc_hd__a21oi_1
X_1263_ _1287_/A1 _1262_/X _1261_/X _1287_/C1 VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__a211o_1
X_1316__10 clkload8/A VGND VGND VPWR VPWR _1459_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0978_ hold6/X _0981_/A _0995_/B VGND VGND VPWR VPWR _0978_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1400__94 clkload7/A VGND VGND VPWR VPWR _1552_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_78_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0763_ _0761_/X _0762_/X _1567_/Q VGND VGND VPWR VPWR _0763_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0901_ _0801_/B _1570_/Q _0889_/Y _0889_/B _1075_/A VGND VGND VPWR VPWR _0902_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0832_ _1556_/Q _1576_/Q VGND VGND VPWR VPWR _0832_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1246_ hold40/A _1285_/A2 _1246_/B1 _1245_/X VGND VGND VPWR VPWR _1246_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1177_ _1486_/Q _1126_/B _1176_/X _1307_/C1 VGND VGND VPWR VPWR _1486_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1413__107 _1483_/CLK VGND VGND VPWR VPWR _1565_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload9/A sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_76_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1100_ _1100_/A _1301_/A VGND VGND VPWR VPWR _1100_/Y sky130_fd_sc_hd__nand2_1
X_1031_ _1075_/B _1138_/A _1030_/X _0915_/A VGND VGND VPWR VPWR _1524_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0815_ _0893_/A _0815_/B VGND VGND VPWR VPWR _1594_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0746_ _1583_/Q VGND VGND VPWR VPWR _0829_/B sky130_fd_sc_hd__inv_2
X_1391__85 _1482_/CLK VGND VGND VPWR VPWR _1543_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ hold33/X _1288_/A2 _1228_/X _1009_/A VGND VGND VPWR VPWR _1469_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_50_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1580_ _1580_/CLK _1580_/D VGND VGND VPWR VPWR _1580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1014_ _1173_/B _1152_/A _1173_/A VGND VGND VPWR VPWR _1030_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ _1559_/Q VGND VGND VPWR VPWR _0729_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1494_ _1494_/CLK _1494_/D VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfxtp_1
X_1419__113 clkload3/A VGND VGND VPWR VPWR _1571_/CLK sky130_fd_sc_hd__inv_2
X_1563_ _1563_/CLK _1563_/D VGND VGND VPWR VPWR _1563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1361__55 clkload2/A VGND VGND VPWR VPWR _1513_/CLK sky130_fd_sc_hd__inv_2
Xfanout49 _1524_/Q VGND VGND VPWR VPWR _0736_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout38 _1530_/Q VGND VGND VPWR VPWR _1016_/A sky130_fd_sc_hd__clkbuf_4
Xfanout16 _0974_/Y VGND VGND VPWR VPWR _1004_/B sky130_fd_sc_hd__clkbuf_2
Xfanout27 _1081_/X VGND VGND VPWR VPWR _1285_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ hold11/A _0967_/D _1538_/Q VGND VGND VPWR VPWR _0995_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1615_ hold9/A VGND VGND VPWR VPWR uio_out[1] sky130_fd_sc_hd__clkbuf_4
X_1477_ _1482_/CLK input3/X VGND VGND VPWR VPWR _1477_/Q sky130_fd_sc_hd__dfxtp_1
X_1546_ _1546_/CLK _1546_/D VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 ui_in[4] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1331__25 _1315__9/A VGND VGND VPWR VPWR _1474_/CLK sky130_fd_sc_hd__inv_2
X_1193_ hold19/A _1587_/Q _1187_/X _1192_/Y _0930_/B VGND VGND VPWR VPWR _1195_/S
+ sky130_fd_sc_hd__o41a_1
X_1262_ _1463_/Q _1461_/Q _1282_/S VGND VGND VPWR VPWR _1262_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ _0973_/X _0995_/B _0977_/C VGND VGND VPWR VPWR _1547_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1529_ _1529_/CLK _1529_/D VGND VGND VPWR VPWR _1529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1397__91 clkload12/A VGND VGND VPWR VPWR _1549_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_60_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _1105_/A _0900_/B VGND VGND VPWR VPWR _1571_/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0762_ hold11/A _1538_/Q hold10/A hold23/A _1565_/Q _1566_/Q VGND VGND VPWR VPWR
+ _0762_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_36_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ hold51/A _1575_/Q VGND VGND VPWR VPWR _0831_/X sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1245_ hold34/A _1245_/B VGND VGND VPWR VPWR _1245_/X sky130_fd_sc_hd__or2_1
X_1176_ _1168_/X _1170_/Y _1174_/X _1175_/X _1137_/B VGND VGND VPWR VPWR _1176_/X
+ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1030_ _1475_/Q _1030_/B VGND VGND VPWR VPWR _1030_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0814_ _0801_/B _1594_/Q _0813_/Y _0813_/B _1071_/B VGND VGND VPWR VPWR _0815_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0745_ _1571_/Q VGND VGND VPWR VPWR _0745_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ _1098_/S _1227_/X _1226_/X _1287_/C1 VGND VGND VPWR VPWR _1228_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1159_ _1520_/Q _0739_/Y _0740_/Y _1519_/Q VGND VGND VPWR VPWR _1159_/X sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1367__61 clkload0/A VGND VGND VPWR VPWR _1519_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_73_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1013_ _1178_/A _1486_/Q VGND VGND VPWR VPWR _1152_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0728_ _1560_/Q VGND VGND VPWR VPWR _0937_/A sky130_fd_sc_hd__inv_2
XFILLER_0_79_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload8/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1493_ _1493_/CLK hold5/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfxtp_1
X_1562_ _1562_/CLK _1562_/D VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfxtp_2
Xfanout28 _1081_/X VGND VGND VPWR VPWR _1246_/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout39 _1289_/A VGND VGND VPWR VPWR _1018_/A sky130_fd_sc_hd__buf_2
XFILLER_0_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1337__31 clkload8/A VGND VGND VPWR VPWR _1489_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0993_ _0993_/A _0993_/B VGND VGND VPWR VPWR _1539_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1614_ _1614_/A VGND VGND VPWR VPWR uio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1476_ _1482_/CLK input2/X VGND VGND VPWR VPWR _1476_/Q sky130_fd_sc_hd__dfxtp_1
X_1545_ _1545_/CLK _1545_/D VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1261_ _1463_/Q _1285_/A2 _1285_/C1 _1260_/X VGND VGND VPWR VPWR _1261_/X sky130_fd_sc_hd__o211a_1
Xinput7 ui_in[5] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
X_1192_ wire17/X _1192_/B VGND VGND VPWR VPWR _1192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0976_ hold29/A hold6/A _0972_/B _1547_/Q VGND VGND VPWR VPWR _0977_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1459_ _1459_/CLK _1459_/D VGND VGND VPWR VPWR _1459_/Q sky130_fd_sc_hd__dfxtp_1
X_1528_ _1528_/CLK _1528_/D VGND VGND VPWR VPWR _1528_/Q sky130_fd_sc_hd__dfxtp_1
X_0830_ _1557_/Q _1577_/Q VGND VGND VPWR VPWR _0830_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0761_ hold27/A _1534_/Q _1535_/Q _1536_/Q _1565_/Q _1566_/Q VGND VGND VPWR VPWR
+ _0761_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1244_ hold40/X _1288_/A2 _1243_/X _1009_/A VGND VGND VPWR VPWR _1466_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1175_ _1149_/Y _1201_/A VGND VGND VPWR VPWR _1175_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ _0942_/X _0959_/B _0963_/B VGND VGND VPWR VPWR _1551_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 uio_in[3] VGND VGND VPWR VPWR _1475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0813_ _0907_/A _0813_/B VGND VGND VPWR VPWR _0813_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0744_ _1570_/Q VGND VGND VPWR VPWR _0744_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1227_ hold32/A hold35/A _1252_/S VGND VGND VPWR VPWR _1227_/X sky130_fd_sc_hd__mux2_1
X_1158_ _1519_/Q _0740_/Y _1117_/A _1518_/Q VGND VGND VPWR VPWR _1158_/X sky130_fd_sc_hd__o22a_1
X_1089_ uo_out[7] _1097_/B _1088_/X _1009_/A VGND VGND VPWR VPWR _1506_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1382__76 clkload12/A VGND VGND VPWR VPWR _1534_/CLK sky130_fd_sc_hd__inv_2
X_1012_ hold36/A _1484_/Q VGND VGND VPWR VPWR _1173_/B sky130_fd_sc_hd__or2_1
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0727_ _1561_/Q VGND VGND VPWR VPWR _0727_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1492_ _1492_/CLK _1492_/D VGND VGND VPWR VPWR _1492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ _1561_/CLK _1561_/D VGND VGND VPWR VPWR _1561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout29 _0864_/Y VGND VGND VPWR VPWR _1285_/A2 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1352__46 _1312__6/A VGND VGND VPWR VPWR _1504_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_13_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ hold10/X _0966_/X _0995_/B VGND VGND VPWR VPWR _0993_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1613_ hold16/A VGND VGND VPWR VPWR uio_oe[7] sky130_fd_sc_hd__buf_2
X_1544_ _1544_/CLK _1544_/D VGND VGND VPWR VPWR _1544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1475_ _1483_/CLK _1475_/D VGND VGND VPWR VPWR _1475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_7_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload7/A sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_80_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1409__103 clkload5/A VGND VGND VPWR VPWR _1561_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 ui_in[6] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
X_1260_ _1461_/Q _1280_/B VGND VGND VPWR VPWR _1260_/X sky130_fd_sc_hd__or2_1
X_1191_ _1191_/A _1191_/B _1191_/C VGND VGND VPWR VPWR _1192_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ hold1/X _0973_/X _0995_/B VGND VGND VPWR VPWR _1548_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1527_ _1527_/CLK _1527_/D VGND VGND VPWR VPWR _1527_/Q sky130_fd_sc_hd__dfxtp_1
X_1322__16 _1315__9/A VGND VGND VPWR VPWR _1465_/CLK sky130_fd_sc_hd__inv_2
X_1458_ _1458_/CLK _1458_/D VGND VGND VPWR VPWR _1458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ _1567_/Q _0759_/X _1568_/Q VGND VGND VPWR VPWR _0760_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1388__82 _1482_/CLK VGND VGND VPWR VPWR _1540_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1243_ _1098_/S _1242_/X _1241_/X _1287_/C1 VGND VGND VPWR VPWR _1243_/X sky130_fd_sc_hd__a211o_1
X_1174_ hold36/A _1152_/A _1125_/Y _1173_/X VGND VGND VPWR VPWR _1174_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0958_ _1551_/Q _0958_/B VGND VGND VPWR VPWR _0959_/B sky130_fd_sc_hd__or2_1
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0889_ _0907_/A _0889_/B VGND VGND VPWR VPWR _0889_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0812_ _1051_/A _1492_/Q _1491_/Q VGND VGND VPWR VPWR _0813_/B sky130_fd_sc_hd__nor3b_4
X_0743_ _1569_/Q VGND VGND VPWR VPWR _0743_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1226_ hold32/A _1285_/A2 _1246_/B1 _1225_/X VGND VGND VPWR VPWR _1226_/X sky130_fd_sc_hd__o211a_1
X_1157_ _1518_/Q _1117_/A _1154_/Y _1156_/Y _1155_/X VGND VGND VPWR VPWR _1157_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1088_ _1291_/D _1246_/B1 _1084_/X _1087_/Y VGND VGND VPWR VPWR _1088_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_50_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1358__52 clkload2/A VGND VGND VPWR VPWR _1510_/CLK sky130_fd_sc_hd__inv_2
X_1011_ hold36/A _1484_/Q VGND VGND VPWR VPWR _1131_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0726_ hold49/A VGND VGND VPWR VPWR _0726_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1209_ _1482_/Q _1295_/A _1298_/A _1481_/Q VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__a22o_1
X_1442__136 clkload6/A VGND VGND VPWR VPWR _1594_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1560_ _1560_/CLK _1560_/D VGND VGND VPWR VPWR _1560_/Q sky130_fd_sc_hd__dfxtp_1
X_1491_ _1491_/CLK _1491_/D VGND VGND VPWR VPWR _1491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328__22 _1312__6/A VGND VGND VPWR VPWR _1471_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ _0991_/A _0991_/B VGND VGND VPWR VPWR _1540_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1612_ hold16/A VGND VGND VPWR VPWR uio_oe[6] sky130_fd_sc_hd__buf_2
X_1474_ _1474_/CLK _1474_/D VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
X_1543_ _1543_/CLK _1543_/D VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1448__142 clkload6/A VGND VGND VPWR VPWR _1600_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 ui_in[7] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
X_1190_ _1592_/Q _1593_/Q _1594_/Q _1595_/Q VGND VGND VPWR VPWR _1191_/C sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_59_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ _0974_/A _0974_/B VGND VGND VPWR VPWR _0974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1526_ _1526_/CLK _1526_/D VGND VGND VPWR VPWR _1526_/Q sky130_fd_sc_hd__dfxtp_1
X_1457_ _1457_/CLK _1457_/D VGND VGND VPWR VPWR _1457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1312__6 _1312__6/A VGND VGND VPWR VPWR _1455_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload6/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1242_ hold41/A hold42/A _1282_/S VGND VGND VPWR VPWR _1242_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1173_ _1173_/A _1173_/B _1173_/C VGND VGND VPWR VPWR _1173_/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ hold12/X _0942_/X _0956_/Y VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0888_ _0888_/A _1051_/B VGND VGND VPWR VPWR _0889_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1509_ _1509_/CLK _1509_/D VGND VGND VPWR VPWR _1509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0742_ _1490_/Q VGND VGND VPWR VPWR _1306_/A sky130_fd_sc_hd__inv_2
X_0811_ _0893_/A _0811_/B VGND VGND VPWR VPWR _1595_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1225_ hold35/A _1245_/B VGND VGND VPWR VPWR _1225_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1087_ _1082_/B _1085_/X _1005_/Y VGND VGND VPWR VPWR _1087_/Y sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_67_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1156_ hold38/A hold25/A VGND VGND VPWR VPWR _1156_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1373__67 _1483_/CLK VGND VGND VPWR VPWR _1525_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ _1486_/Q _1178_/A VGND VGND VPWR VPWR _1173_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_29_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0725_ _1009_/A VGND VGND VPWR VPWR _1068_/A sky130_fd_sc_hd__inv_2
X_1208_ _1480_/Q _1301_/A _1207_/A _1024_/A VGND VGND VPWR VPWR _1208_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1139_ hold43/A _1139_/B VGND VGND VPWR VPWR _1145_/B sky130_fd_sc_hd__or2_1
XFILLER_0_62_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1490_ _1490_/CLK _1490_/D VGND VGND VPWR VPWR _1490_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1343__37 clkload1/A VGND VGND VPWR VPWR _1495_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1611_ hold16/A VGND VGND VPWR VPWR uio_oe[2] sky130_fd_sc_hd__buf_2
X_0990_ hold23/X _0993_/A _0995_/B VGND VGND VPWR VPWR _0991_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1542_ _1542_/CLK _1542_/D VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__dfxtp_1
X_1473_ _1473_/CLK _1473_/D VGND VGND VPWR VPWR _1618_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ hold6/A _1547_/Q _0981_/A VGND VGND VPWR VPWR _0973_/X sky130_fd_sc_hd__and3_1
X_1525_ _1525_/CLK _1525_/D VGND VGND VPWR VPWR _1525_/Q sky130_fd_sc_hd__dfxtp_1
X_1456_ _1456_/CLK _1456_/D VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1241_ hold41/A _1285_/A2 _1246_/B1 _1240_/X VGND VGND VPWR VPWR _1241_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _1178_/A _1126_/B _1171_/X _1307_/C1 VGND VGND VPWR VPWR _1487_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ hold12/A _0942_/X _0963_/B VGND VGND VPWR VPWR _0956_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1379__73 _1483_/CLK VGND VGND VPWR VPWR _1531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0887_ _1492_/Q _1491_/Q VGND VGND VPWR VPWR _1051_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1508_ _1508_/CLK _1508_/D VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0810_ _0801_/B _1595_/Q _0792_/Y _0792_/A _0736_/A VGND VGND VPWR VPWR _0811_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0741_ hold37/X VGND VGND VPWR VPWR _1117_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1224_ hold32/X _1218_/Y _1223_/X _1288_/C1 VGND VGND VPWR VPWR _1470_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1086_ _1082_/B _1085_/X _1005_/Y VGND VGND VPWR VPWR _1097_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1155_ _1496_/Q hold52/A VGND VGND VPWR VPWR _1155_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0939_ _1559_/Q _0925_/D _0937_/B _0953_/C VGND VGND VPWR VPWR _1559_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload5/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1349__43 clkload0/A VGND VGND VPWR VPWR _1501_/CLK sky130_fd_sc_hd__inv_2
X_1207_ _1207_/A _1207_/B VGND VGND VPWR VPWR _1207_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1138_ _1138_/A _1138_/B VGND VGND VPWR VPWR _1139_/B sky130_fd_sc_hd__nor2_1
X_1069_ _1072_/A _1069_/B VGND VGND VPWR VPWR _1069_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1610_ hold16/A VGND VGND VPWR VPWR uio_oe[1] sky130_fd_sc_hd__buf_2
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1472_ _1472_/CLK _1472_/D VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfxtp_1
X_1541_ _1541_/CLK _1541_/D VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
X_1319__13 clkload8/A VGND VGND VPWR VPWR _1462_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1432__126 clkload4/A VGND VGND VPWR VPWR _1584_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1403__97 clkload5/A VGND VGND VPWR VPWR _1555_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ hold29/A _0972_/B VGND VGND VPWR VPWR _0981_/A sky130_fd_sc_hd__and2_1
XFILLER_0_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1524_ _1524_/CLK _1524_/D VGND VGND VPWR VPWR _1524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1455_ _1455_/CLK _1455_/D VGND VGND VPWR VPWR uo_out[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1240_ hold42/A _1280_/B VGND VGND VPWR VPWR _1240_/X sky130_fd_sc_hd__or2_1
X_1171_ _1298_/A _1168_/X _1170_/B _1151_/X VGND VGND VPWR VPWR _1171_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0955_ _0952_/B _0955_/B _0963_/B VGND VGND VPWR VPWR _1553_/D sky130_fd_sc_hd__and3b_1
X_0886_ _0886_/A _0886_/B VGND VGND VPWR VPWR _1577_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1507_ _1507_/CLK _1507_/D VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
X_1394__88 _1482_/CLK VGND VGND VPWR VPWR _1546_/CLK sky130_fd_sc_hd__inv_2
X_1438__132 _1313__7/A VGND VGND VPWR VPWR _1590_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap18 _1178_/Y VGND VGND VPWR VPWR _1186_/B1 sky130_fd_sc_hd__buf_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtt_um_jimktrains_vslc_63 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_63/HI uio_oe[3]
+ sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_61_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ hold17/A VGND VGND VPWR VPWR _0740_/Y sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_70_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1223_ _1098_/S _1222_/X _1221_/X _1219_/X VGND VGND VPWR VPWR _1223_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_67_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1154_ hold52/A _1496_/Q VGND VGND VPWR VPWR _1154_/Y sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_75_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1085_ _1018_/A _1020_/A _1291_/D VGND VGND VPWR VPWR _1085_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_47_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0869_ _1491_/Q _1492_/Q VGND VGND VPWR VPWR _1033_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0938_ _0924_/Y _0953_/C _0938_/C VGND VGND VPWR VPWR _1560_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1364__58 clkload3/A VGND VGND VPWR VPWR _1516_/CLK sky130_fd_sc_hd__inv_2
X_1206_ _1479_/Q _1069_/Y _1301_/A _1476_/Q VGND VGND VPWR VPWR _1206_/X sky130_fd_sc_hd__a22o_1
X_1137_ _1201_/A _1137_/B VGND VGND VPWR VPWR _1138_/B sky130_fd_sc_hd__or2_1
X_1068_ _1068_/A hold16/X VGND VGND VPWR VPWR _1507_/D sky130_fd_sc_hd__or2_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload4/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ _1540_/CLK _1540_/D VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ _1471_/CLK _1471_/D VGND VGND VPWR VPWR _1471_/Q sky130_fd_sc_hd__dfxtp_1
X_1334__28 clkload8/A VGND VGND VPWR VPWR _1486_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0971_ hold7/A _1544_/Q _0987_/A VGND VGND VPWR VPWR _0972_/B sky130_fd_sc_hd__and3_1
XFILLER_0_39_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1454_ _1454_/CLK _1454_/D VGND VGND VPWR VPWR uo_out[2] sky130_fd_sc_hd__dfxtp_4
X_1523_ _1523_/CLK _1523_/D VGND VGND VPWR VPWR _1523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _1298_/A _1170_/B VGND VGND VPWR VPWR _1170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0954_ hold12/A _0942_/X _1553_/Q VGND VGND VPWR VPWR _0955_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0885_ _0801_/B _1577_/Q _0871_/Y _0871_/B _0736_/A VGND VGND VPWR VPWR _0886_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1506_ _1506_/CLK _1506_/D VGND VGND VPWR VPWR uo_out[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1299_ _1298_/A _1301_/B uo_out[1] VGND VGND VPWR VPWR _1299_/X sky130_fd_sc_hd__a21o_1
Xmax_cap19 _1180_/A3 VGND VGND VPWR VPWR _1170_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_jimktrains_vslc_64 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_64/HI uio_oe[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1084_ _1024_/A _1292_/A _1292_/B _1287_/A1 _1083_/X VGND VGND VPWR VPWR _1084_/X
+ sky130_fd_sc_hd__o311a_1
X_1222_ _1532_/Q hold33/A _1252_/S VGND VGND VPWR VPWR _1222_/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1153_ hold44/A hold21/A VGND VGND VPWR VPWR _1153_/Y sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_75_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0868_ _0860_/X _0867_/Y _0862_/X VGND VGND VPWR VPWR _1585_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0799_ _0893_/A _1528_/Q VGND VGND VPWR VPWR _0800_/A sky130_fd_sc_hd__and2_2
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0937_ _0937_/A _0937_/B VGND VGND VPWR VPWR _0938_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1205_ hold2/X _1138_/B _1204_/X VGND VGND VPWR VPWR _1472_/D sky130_fd_sc_hd__o21ba_1
X_1136_ _1178_/A _1486_/Q _1152_/B _1135_/X VGND VGND VPWR VPWR _1137_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1067_ _0736_/A _1051_/X _1066_/X _1145_/A VGND VGND VPWR VPWR _1508_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1315__9 _1315__9/A VGND VGND VPWR VPWR _1458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _1117_/B _1119_/B VGND VGND VPWR VPWR _1496_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1470_ _1470_/CLK _1470_/D VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1599_ _1599_/CLK _1599_/D VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_3_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload3/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0970_ hold30/A _0989_/A VGND VGND VPWR VPWR _0987_/A sky130_fd_sc_hd__and2_1
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ _1453_/CLK _1453_/D VGND VGND VPWR VPWR uo_out[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1522_ _1522_/CLK _1522_/D VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1422__116 clkload1/A VGND VGND VPWR VPWR _1574_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0953_ _0946_/C _0953_/B _0953_/C VGND VGND VPWR VPWR _1554_/D sky130_fd_sc_hd__and3b_1
X_0884_ _0886_/A _0884_/B VGND VGND VPWR VPWR _1578_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1505_ _1505_/CLK _1505_/D VGND VGND VPWR VPWR uo_out[6] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ _1298_/A _1301_/B VGND VGND VPWR VPWR _1298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_jimktrains_vslc_65 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_65/HI uio_oe[5]
+ sky130_fd_sc_hd__conb_1
X_1385__79 clkload12/A VGND VGND VPWR VPWR _1537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1221_ _1532_/Q _0864_/Y _1285_/C1 _1220_/X VGND VGND VPWR VPWR _1221_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1083_ _1100_/A _1525_/Q _1075_/B uo_out[7] VGND VGND VPWR VPWR _1083_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_59_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1152_ _1152_/A _1152_/B VGND VGND VPWR VPWR _1168_/A sky130_fd_sc_hd__and2_1
XFILLER_0_74_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0936_ _1561_/Q _0924_/Y _0926_/Y _0953_/C VGND VGND VPWR VPWR _1561_/D sky130_fd_sc_hd__o211a_1
X_0867_ _0867_/A _1291_/C _0867_/C _1169_/C VGND VGND VPWR VPWR _0867_/Y sky130_fd_sc_hd__nand4_1
X_0798_ _0893_/A _0798_/B VGND VGND VPWR VPWR _1600_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1428__122 clkload4/A VGND VGND VPWR VPWR _1580_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ _1138_/B _1199_/Y _1203_/X _1068_/A VGND VGND VPWR VPWR _1204_/X sky130_fd_sc_hd__a31o_1
X_1135_ _1178_/A _1486_/Q hold36/A _1484_/Q VGND VGND VPWR VPWR _1135_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1066_ hold53/X _1066_/B VGND VGND VPWR VPWR _1066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0919_ _0960_/B _0944_/C _0921_/D VGND VGND VPWR VPWR _0920_/A sky130_fd_sc_hd__and3_1
XFILLER_0_35_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1355__49 _1315__9/A VGND VGND VPWR VPWR _1507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1049_ _0736_/A _1033_/X _1048_/X _0886_/A VGND VGND VPWR VPWR _1516_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1118_ _1105_/A hold25/A _1105_/D _1496_/Q VGND VGND VPWR VPWR _1119_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1325__19 _1315__9/A VGND VGND VPWR VPWR _1468_/CLK sky130_fd_sc_hd__inv_2
X_1598_ _1598_/CLK _1598_/D VGND VGND VPWR VPWR _1598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1452_ _1452_/CLK _1452_/D VGND VGND VPWR VPWR uo_out[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1521_ _1521_/CLK _1521_/D VGND VGND VPWR VPWR _1521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ _1554_/Q _0952_/B VGND VGND VPWR VPWR _0953_/B sky130_fd_sc_hd__or2_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1504_ _1504_/CLK _1504_/D VGND VGND VPWR VPWR uo_out[5] sky130_fd_sc_hd__dfxtp_4
X_0883_ _0899_/A1 _1578_/Q _0871_/Y _0871_/B _1075_/A VGND VGND VPWR VPWR _0884_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1297_ _1292_/B _1295_/Y _1296_/X _1294_/A VGND VGND VPWR VPWR _1454_/D sky130_fd_sc_hd__o211a_1
X_1445__139 _1313__7/A VGND VGND VPWR VPWR _1597_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload2/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_jimktrains_vslc_66 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_66/HI uio_out[3]
+ sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_21_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ hold33/A _1245_/B VGND VGND VPWR VPWR _1220_/X sky130_fd_sc_hd__or2_1
X_1151_ _1173_/A _1131_/C _1125_/Y _1137_/B _1150_/X VGND VGND VPWR VPWR _1151_/X
+ sky130_fd_sc_hd__a2111o_1
X_1082_ _1071_/A _1082_/B VGND VGND VPWR VPWR _1082_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0866_ _1018_/A _1020_/A VGND VGND VPWR VPWR _1169_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ hold49/A _0928_/C _0927_/Y _0953_/C VGND VGND VPWR VPWR _1562_/D sky130_fd_sc_hd__o211a_1
X_0797_ _0801_/B _1600_/Q _0792_/Y _0792_/A _1289_/A VGND VGND VPWR VPWR _0798_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1134_ hold36/A _1484_/Q VGND VGND VPWR VPWR _1152_/B sky130_fd_sc_hd__and2b_1
X_1203_ _1489_/Q _1201_/Y _1202_/Y _1201_/A _1490_/Q VGND VGND VPWR VPWR _1203_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1065_ _1075_/A _1051_/X _1064_/X _1145_/A VGND VGND VPWR VPWR _1509_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0918_ _1557_/Q _1556_/Q hold51/A _1554_/Q VGND VGND VPWR VPWR _0921_/D sky130_fd_sc_hd__and4_1
X_0849_ _0849_/A _0849_/B _0849_/C _0849_/D VGND VGND VPWR VPWR _0850_/C sky130_fd_sc_hd__nand4_1
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ _1117_/A _1117_/B VGND VGND VPWR VPWR _1497_/D sky130_fd_sc_hd__xnor2_1
X_1048_ hold38/X _1048_/B VGND VGND VPWR VPWR _1048_/X sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1597_ _1597_/CLK _1597_/D VGND VGND VPWR VPWR _1597_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_77_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1520_ _1520_/CLK _1520_/D VGND VGND VPWR VPWR _1520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1451_ _1451_/CLK _1451_/D VGND VGND VPWR VPWR _1617_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0951_ _0951_/A _0951_/B VGND VGND VPWR VPWR _1555_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0882_ _0886_/A _0882_/B VGND VGND VPWR VPWR _1579_/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_30_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1503_ _1503_/CLK _1503_/D VGND VGND VPWR VPWR uo_out[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1296_ _1295_/A _1301_/B uo_out[2] VGND VGND VPWR VPWR _1296_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtt_um_jimktrains_vslc_67 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_67/HI uio_out[4]
+ sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ _1178_/A _1133_/Y _1149_/Y _1201_/A VGND VGND VPWR VPWR _1150_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1081_ _1071_/A _1082_/B VGND VGND VPWR VPWR _1081_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_59_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0865_ _1471_/Q _1280_/B VGND VGND VPWR VPWR _0867_/C sky130_fd_sc_hd__or2_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ _0931_/B _0953_/C _0934_/C VGND VGND VPWR VPWR _1563_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0796_ _0893_/A _0796_/B VGND VGND VPWR VPWR _1601_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1412__106 clkload5/A VGND VGND VPWR VPWR _1564_/CLK sky130_fd_sc_hd__inv_2
X_1390__84 _1482_/CLK VGND VGND VPWR VPWR _1542_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1279_ _1459_/Q _1288_/A2 _1278_/X _1307_/C1 VGND VGND VPWR VPWR _1459_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_21_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1133_ _1486_/Q _1173_/C VGND VGND VPWR VPWR _1133_/Y sky130_fd_sc_hd__nor2_1
X_1202_ _1489_/Q _1202_/B VGND VGND VPWR VPWR _1202_/Y sky130_fd_sc_hd__nor2_1
X_1064_ _1509_/Q _1066_/B VGND VGND VPWR VPWR _1064_/X sky130_fd_sc_hd__or2_1
Xclkbuf_4_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload1/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0779_ _1563_/Q _1601_/Q VGND VGND VPWR VPWR _0779_/Y sky130_fd_sc_hd__xnor2_1
X_0917_ _1553_/Q hold12/A _1551_/Q _1550_/Q VGND VGND VPWR VPWR _0944_/C sky130_fd_sc_hd__and4_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0848_ _0729_/Y _1579_/Q _1580_/Q _0937_/A _0832_/Y VGND VGND VPWR VPWR _0849_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1360__54 clkload2/A VGND VGND VPWR VPWR _1512_/CLK sky130_fd_sc_hd__inv_2
X_1047_ _1075_/A _1033_/X _1046_/X _0886_/A VGND VGND VPWR VPWR _1517_/D sky130_fd_sc_hd__o211a_1
X_1116_ _1116_/A hold18/X VGND VGND VPWR VPWR _1498_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_75_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1418__112 clkload4/A VGND VGND VPWR VPWR _1570_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ _1596_/CLK _1596_/D VGND VGND VPWR VPWR _1596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1330__24 _1313__7/A VGND VGND VPWR VPWR _1473_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1579_ _1579_/CLK _1579_/D VGND VGND VPWR VPWR _1579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1396__90 _1483_/CLK VGND VGND VPWR VPWR _1548_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ hold51/X _0946_/C _0953_/C VGND VGND VPWR VPWR _0951_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0881_ _0899_/A1 _1579_/Q _0871_/Y _0871_/B _1063_/A1 VGND VGND VPWR VPWR _0882_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_30_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1502_ _1502_/CLK _1502_/D VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
X_1295_ _1295_/A _1301_/B VGND VGND VPWR VPWR _1295_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtt_um_jimktrains_vslc_68 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_68/HI uio_out[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ _0856_/X _1207_/B _1071_/X _1471_/Q VGND VGND VPWR VPWR _1292_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_67_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0864_ _1020_/A _1018_/A VGND VGND VPWR VPWR _0864_/Y sky130_fd_sc_hd__nand2b_2
X_0795_ _0801_/B _1601_/Q _0792_/Y _0792_/A _1016_/A VGND VGND VPWR VPWR _0796_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0933_ hold49/A _0928_/C _1563_/Q VGND VGND VPWR VPWR _0934_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1278_ _1287_/A1 _1277_/X _1276_/X _1287_/C1 VGND VGND VPWR VPWR _1278_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1366__60 clkload1/A VGND VGND VPWR VPWR _1518_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1435__129 _1313__7/A VGND VGND VPWR VPWR _1587_/CLK sky130_fd_sc_hd__inv_2
X_1201_ _1201_/A _1201_/B VGND VGND VPWR VPWR _1201_/Y sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_0_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1132_ hold36/A _1484_/Q VGND VGND VPWR VPWR _1173_/C sky130_fd_sc_hd__nand2_1
X_1063_ _1063_/A1 _1051_/X _1062_/X _1063_/C1 VGND VGND VPWR VPWR _1510_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ _0758_/X _0760_/X _0763_/X _1568_/Q _1549_/Q VGND VGND VPWR VPWR _0960_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0778_ hold51/A _0750_/Y _1596_/Q _0730_/Y VGND VGND VPWR VPWR _0778_/X sky130_fd_sc_hd__a2bb2o_1
X_0847_ _0733_/Y hold14/A hold20/A _0727_/Y _0830_/Y VGND VGND VPWR VPWR _0849_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1046_ hold52/X _1048_/B VGND VGND VPWR VPWR _1046_/X sky130_fd_sc_hd__or2_1
X_1115_ hold37/A _1117_/B hold17/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1336__30 clkload8/A VGND VGND VPWR VPWR _1488_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload0/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _1595_/CLK _1595_/D VGND VGND VPWR VPWR _1595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1029_ _1075_/A _1138_/A _1028_/Y _0915_/A VGND VGND VPWR VPWR _1525_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1578_ _1578_/CLK _1578_/D VGND VGND VPWR VPWR _1578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ _0886_/A _0880_/B VGND VGND VPWR VPWR _1580_/D sky130_fd_sc_hd__and2_1
X_1501_ _1501_/CLK _1501_/D VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1294_ _1294_/A _1294_/B _1294_/C VGND VGND VPWR VPWR _1455_/D sky130_fd_sc_hd__and3_1
XFILLER_0_41_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0932_ _0932_/A _0953_/C _0932_/C VGND VGND VPWR VPWR _1564_/D sky130_fd_sc_hd__and3_1
X_0863_ _1020_/A _1018_/A VGND VGND VPWR VPWR _1245_/B sky130_fd_sc_hd__and2b_1
X_0794_ _0893_/A _0794_/B VGND VGND VPWR VPWR _1602_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1277_ _1460_/Q _1458_/Q _1282_/S VGND VGND VPWR VPWR _1277_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1381__75 clkload12/A VGND VGND VPWR VPWR _1533_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1200_ hold53/A _1509_/Q hold43/A VGND VGND VPWR VPWR _1202_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1131_ _1178_/A _1486_/Q _1131_/C VGND VGND VPWR VPWR _1201_/A sky130_fd_sc_hd__and3_1
X_1062_ hold48/X _1066_/B VGND VGND VPWR VPWR _1062_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ _0915_/A _0915_/B VGND VGND VPWR VPWR _1565_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0777_ _1589_/Q _1551_/Q VGND VGND VPWR VPWR _0777_/Y sky130_fd_sc_hd__nand2b_1
X_0846_ _0846_/A _0846_/B VGND VGND VPWR VPWR _0849_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1114_ _1114_/A _1114_/B VGND VGND VPWR VPWR _1499_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ _1063_/A1 _1033_/X _1044_/X _1105_/A VGND VGND VPWR VPWR _1518_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_43_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0829_ _1563_/Q _0829_/B VGND VGND VPWR VPWR _0829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1351__45 _1315__9/A VGND VGND VPWR VPWR _1503_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1594_ _1594_/CLK _1594_/D VGND VGND VPWR VPWR _1594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_37_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1028_ _1069_/B _1138_/A VGND VGND VPWR VPWR _1028_/Y sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_46_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1408__102 clkload5/A VGND VGND VPWR VPWR _1560_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1577_ _1577_/CLK _1577_/D VGND VGND VPWR VPWR _1577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1321__15 _1315__9/A VGND VGND VPWR VPWR _1464_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1500_ _1500_/CLK _1500_/D VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfxtp_1
X_1293_ _1069_/Y _1301_/B uo_out[3] VGND VGND VPWR VPWR _1294_/C sky130_fd_sc_hd__a21o_1
X_1387__81 _1482_/CLK VGND VGND VPWR VPWR _1539_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0862_ _0862_/A _0974_/B _0860_/X VGND VGND VPWR VPWR _0862_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_55_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0931_ _1564_/Q _0931_/B VGND VGND VPWR VPWR _0932_/C sky130_fd_sc_hd__nand2_1
X_0793_ _0801_/B _1602_/Q _0792_/Y _0792_/A _1071_/B VGND VGND VPWR VPWR _0794_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_66_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1276_ _1460_/Q _1285_/A2 _1285_/C1 _1275_/X VGND VGND VPWR VPWR _1276_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1357__51 clkload2/A VGND VGND VPWR VPWR _1509_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1130_ _1484_/Q _1491_/Q _1130_/S VGND VGND VPWR VPWR _1491_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1061_ _1207_/A _1051_/X _1060_/X _1063_/C1 VGND VGND VPWR VPWR _1511_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ _1196_/B _1565_/Q _0907_/Y _0907_/B _1075_/B VGND VGND VPWR VPWR _0915_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0845_ _1558_/Q _1578_/Q VGND VGND VPWR VPWR _0846_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0776_ _1551_/Q _1589_/Q VGND VGND VPWR VPWR _0776_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1259_ _1463_/Q _1288_/A2 _1258_/X _1307_/C1 VGND VGND VPWR VPWR _1463_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1310__4 _1312__6/A VGND VGND VPWR VPWR _1453_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1441__135 _1313__7/A VGND VGND VPWR VPWR _1593_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_52_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ hold24/X _1116_/A VGND VGND VPWR VPWR _1114_/B sky130_fd_sc_hd__nor2_1
X_1044_ _1518_/Q _1048_/B VGND VGND VPWR VPWR _1044_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0759_ hold29/A hold6/A _1547_/Q hold1/A _1565_/Q _1566_/Q VGND VGND VPWR VPWR _0759_/X
+ sky130_fd_sc_hd__mux4_1
X_0828_ _1196_/A _0828_/B VGND VGND VPWR VPWR _1587_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1425__119 clkload6/A VGND VGND VPWR VPWR _1577_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1327__21 _1312__6/A VGND VGND VPWR VPWR _1470_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_57_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1593_ _1593_/CLK _1593_/D VGND VGND VPWR VPWR _1593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ _1169_/B _1138_/A _1026_/Y _1294_/A VGND VGND VPWR VPWR _1526_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1447__141 clkload6/A VGND VGND VPWR VPWR _1599_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1576_ _1576_/CLK _1576_/D VGND VGND VPWR VPWR _1576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ _1292_/A _1292_/B _1301_/B VGND VGND VPWR VPWR _1294_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1559_ _1559_/CLK _1559_/D VGND VGND VPWR VPWR _1559_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ _0974_/B _0930_/B VGND VGND VPWR VPWR _0930_/Y sky130_fd_sc_hd__nor2_1
X_0861_ _1291_/D _1289_/C _0856_/X _0907_/A VGND VGND VPWR VPWR _0862_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_55_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0792_ _0792_/A _0907_/A VGND VGND VPWR VPWR _0792_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1275_ _1458_/Q _1280_/B VGND VGND VPWR VPWR _1275_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1372__66 _1483_/CLK VGND VGND VPWR VPWR _1524_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ hold54/X _1066_/B VGND VGND VPWR VPWR _1060_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0913_ _1294_/A _0913_/B VGND VGND VPWR VPWR _1566_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0775_ _1559_/Q _1597_/Q VGND VGND VPWR VPWR _0775_/X sky130_fd_sc_hd__and2b_1
X_0844_ hold12/A _1572_/Q VGND VGND VPWR VPWR _0846_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1258_ _1287_/A1 _1257_/X _1256_/X _1287_/C1 VGND VGND VPWR VPWR _1258_/X sky130_fd_sc_hd__a211o_1
X_1189_ _1596_/Q _1597_/Q _1598_/Q hold26/A VGND VGND VPWR VPWR _1191_/B sky130_fd_sc_hd__or4_1
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1043_ _1207_/A _1033_/X _1042_/X _1105_/A VGND VGND VPWR VPWR _1519_/D sky130_fd_sc_hd__o211a_1
X_1112_ _1112_/A _1114_/A VGND VGND VPWR VPWR _1500_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0758_ _1567_/Q _0758_/B VGND VGND VPWR VPWR _0758_/X sky130_fd_sc_hd__and2b_1
X_0827_ _1196_/B _1587_/Q _0813_/Y _0813_/B _1075_/B VGND VGND VPWR VPWR _0828_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1342__36 clkload3/A VGND VGND VPWR VPWR _1494_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1592_ _1592_/CLK _1592_/D VGND VGND VPWR VPWR _1592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1026_ _1072_/A _1138_/A VGND VGND VPWR VPWR _1026_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1575_ _1575_/CLK _1575_/D VGND VGND VPWR VPWR _1575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ _1009_/A _1009_/B _1009_/C VGND VGND VPWR VPWR _1532_/D sky130_fd_sc_hd__and3_1
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1291_ _1100_/A _1289_/C _1291_/C _1291_/D VGND VGND VPWR VPWR _1301_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1378__72 _1483_/CLK VGND VGND VPWR VPWR _1530_/CLK sky130_fd_sc_hd__inv_2
X_1489_ _1489_/CLK _1489_/D VGND VGND VPWR VPWR _1489_/Q sky130_fd_sc_hd__dfxtp_2
X_1558_ _1558_/CLK _1558_/D VGND VGND VPWR VPWR _1558_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ _1291_/D _1289_/C _1252_/S _0856_/X VGND VGND VPWR VPWR _0860_/X sky130_fd_sc_hd__or4b_1
X_0791_ hold19/A _0974_/A wire17/X VGND VGND VPWR VPWR _0907_/A sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_79_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1274_ _1460_/Q _1288_/A2 _1273_/X _1307_/C1 VGND VGND VPWR VPWR _1460_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0989_/A _0989_/B VGND VGND VPWR VPWR _1541_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ _0912_/A1 _1566_/Q _0907_/Y _0907_/B _1075_/A VGND VGND VPWR VPWR _0913_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0774_ _1553_/Q hold46/A VGND VGND VPWR VPWR _0774_/X sky130_fd_sc_hd__and2b_1
X_0843_ _1550_/Q _0744_/Y _1582_/Q _0726_/Y _0842_/Y VGND VGND VPWR VPWR _0849_/A
+ sky130_fd_sc_hd__o221a_1
X_1348__42 clkload0/A VGND VGND VPWR VPWR _1500_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1257_ hold34/A _1462_/Q _1282_/S VGND VGND VPWR VPWR _1257_/X sky130_fd_sc_hd__mux2_1
X_1188_ _1600_/Q _1601_/Q _1602_/Q VGND VGND VPWR VPWR _1191_/A sky130_fd_sc_hd__or3_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1111_ _1111_/A hold22/X VGND VGND VPWR VPWR _1501_/D sky130_fd_sc_hd__nor2_1
X_1042_ _1519_/Q _1048_/B VGND VGND VPWR VPWR _1042_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0757_ hold8/A hold30/A hold7/A _1544_/Q _1565_/Q _1566_/Q VGND VGND VPWR VPWR _0758_/B
+ sky130_fd_sc_hd__mux4_1
X_0826_ _0867_/A _0826_/B VGND VGND VPWR VPWR _1588_/D sky130_fd_sc_hd__nand2_1
Xclkbuf_4_15_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1482_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1318__12 clkload8/A VGND VGND VPWR VPWR _1461_/CLK sky130_fd_sc_hd__inv_2
X_1591_ _1591_/CLK _1591_/D VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1025_ _1207_/A _1138_/A _1024_/Y _0915_/A VGND VGND VPWR VPWR _1527_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_72_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0809_ _0867_/A _0809_/B VGND VGND VPWR VPWR _1596_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1431__125 clkload4/A VGND VGND VPWR VPWR _1583_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_24_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1402__96 clkload7/A VGND VGND VPWR VPWR _1554_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_42_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1415__109 _1482_/CLK VGND VGND VPWR VPWR _1567_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_60_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1574_ _1574_/CLK _1574_/D VGND VGND VPWR VPWR _1574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1008_ _0906_/C _1005_/Y _1532_/Q VGND VGND VPWR VPWR _1009_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1290_ _1075_/B hold19/X _1290_/S VGND VGND VPWR VPWR _1456_/D sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1393__87 _1482_/CLK VGND VGND VPWR VPWR _1545_/CLK sky130_fd_sc_hd__inv_2
X_1488_ _1488_/CLK _1488_/D VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_4
X_1557_ _1557_/CLK _1557_/D VGND VGND VPWR VPWR _1557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1437__131 _1313__7/A VGND VGND VPWR VPWR _1589_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0790_ _0790_/A _0790_/B _0790_/C _0789_/X VGND VGND VPWR VPWR wire17/A sky130_fd_sc_hd__nor4b_1
XFILLER_0_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1273_ _1287_/A1 _1272_/X _1271_/X _1287_/C1 VGND VGND VPWR VPWR _1273_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ hold8/X _0991_/A _0995_/B VGND VGND VPWR VPWR _0989_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1609_ hold16/A VGND VGND VPWR VPWR uio_oe[0] sky130_fd_sc_hd__buf_2
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0911_ _1294_/A _0911_/B VGND VGND VPWR VPWR _1567_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0842_ _1554_/Q _1574_/Q VGND VGND VPWR VPWR _0842_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0773_ _0727_/Y hold26/A _0752_/Y hold49/A VGND VGND VPWR VPWR _0773_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1256_ hold34/A _1285_/A2 _1285_/C1 _1255_/X VGND VGND VPWR VPWR _1256_/X sky130_fd_sc_hd__o211a_1
X_1363__57 clkload2/A VGND VGND VPWR VPWR _1515_/CLK sky130_fd_sc_hd__inv_2
X_1187_ _1588_/Q _1589_/Q _1590_/Q hold46/A VGND VGND VPWR VPWR _1187_/X sky130_fd_sc_hd__or4_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ hold31/A _1114_/A hold21/X VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _1020_/A _1033_/X _1040_/X _1063_/C1 VGND VGND VPWR VPWR _1520_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0825_ _0912_/A1 _0748_/Y _0813_/Y _0813_/B _1072_/A VGND VGND VPWR VPWR _0826_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0756_ _1492_/Q _1491_/Q _1051_/A VGND VGND VPWR VPWR _0792_/A sky130_fd_sc_hd__nor3_4
X_1308_ hold9/A _1308_/B VGND VGND VPWR VPWR _1614_/A sky130_fd_sc_hd__nor2_2
X_1239_ hold41/X _1218_/Y _1238_/X _1009_/A VGND VGND VPWR VPWR _1467_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ _1590_/CLK _1590_/D VGND VGND VPWR VPWR _1590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ _1024_/A _1138_/A VGND VGND VPWR VPWR _1024_/Y sky130_fd_sc_hd__nand2_1
X_1333__27 clkload9/A VGND VGND VPWR VPWR _1485_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0808_ _0912_/A1 _1596_/Q _0792_/Y _0792_/A _1075_/A VGND VGND VPWR VPWR _0809_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0739_ hold24/A VGND VGND VPWR VPWR _0739_/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1399__93 clkload12/A VGND VGND VPWR VPWR _1551_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1483_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1573_ _1573_/CLK _1573_/D VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1007_ _1007_/A hold32/A _0906_/C VGND VGND VPWR VPWR _1009_/B sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_49_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1556_ _1556_/CLK _1556_/D VGND VGND VPWR VPWR _1556_/Q sky130_fd_sc_hd__dfxtp_1
X_1487_ _1487_/CLK _1487_/D VGND VGND VPWR VPWR _1487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1313__7 _1313__7/A VGND VGND VPWR VPWR _1456_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1369__63 clkload0/A VGND VGND VPWR VPWR _1521_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1272_ _1461_/Q _1459_/Q _1282_/S VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0987_ _0987_/A _0987_/B VGND VGND VPWR VPWR _1542_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1539_ _1539_/CLK _1539_/D VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0910_ _0912_/A1 _1567_/Q _0907_/Y _0907_/B _1100_/A VGND VGND VPWR VPWR _0911_/B
+ sky130_fd_sc_hd__a32o_1
X_0772_ _1560_/Q _1598_/Q VGND VGND VPWR VPWR _0772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0841_ _0841_/A _0841_/B _0841_/C _0841_/D VGND VGND VPWR VPWR _0850_/B sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1186_ hold9/X _1139_/B _1186_/B1 _1068_/A VGND VGND VPWR VPWR _1474_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1255_ _1462_/Q _1280_/B VGND VGND VPWR VPWR _1255_/X sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1339__33 clkload3/A VGND VGND VPWR VPWR _1491_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ _1520_/Q _1048_/B VGND VGND VPWR VPWR _1040_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0824_ _1196_/A _0824_/B VGND VGND VPWR VPWR _1589_/D sky130_fd_sc_hd__and2_1
X_0755_ hold4/A _0854_/A hold3/A VGND VGND VPWR VPWR _1051_/A sky130_fd_sc_hd__or3b_4
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1238_ _1098_/S _1237_/X _1236_/X _1219_/X VGND VGND VPWR VPWR _1238_/X sky130_fd_sc_hd__a211o_1
X_1169_ _1291_/D _1169_/B _1169_/C _1289_/D VGND VGND VPWR VPWR _1182_/C sky130_fd_sc_hd__nor4_1
X_1307_ _1490_/Q _1304_/X _1306_/X _1307_/C1 VGND VGND VPWR VPWR _1451_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ _1207_/A _1030_/B _1120_/B _1289_/B VGND VGND VPWR VPWR _1528_/D sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_56_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0807_ _0893_/A _0807_/B VGND VGND VPWR VPWR _1597_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0738_ hold31/X VGND VGND VPWR VPWR _1112_/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1572_ _1572_/CLK _1572_/D VGND VGND VPWR VPWR _1572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ _1071_/A _1289_/C VGND VGND VPWR VPWR _1007_/A sky130_fd_sc_hd__or2_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1421__115 clkload6/A VGND VGND VPWR VPWR _1573_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1555_ _1555_/CLK _1555_/D VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_77_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _1486_/CLK _1486_/D VGND VGND VPWR VPWR _1486_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1384__78 clkload12/A VGND VGND VPWR VPWR _1536_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_4_13_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload12/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire17 wire17/A VGND VGND VPWR VPWR wire17/X sky130_fd_sc_hd__buf_1
X_1271_ _1461_/Q _1285_/A2 _1285_/C1 _1270_/X VGND VGND VPWR VPWR _1271_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ hold30/X _0989_/A _0995_/B VGND VGND VPWR VPWR _0987_/B sky130_fd_sc_hd__o21ai_1
X_1469_ _1469_/CLK _1469_/D VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dfxtp_1
X_1538_ _1538_/CLK _1538_/D VGND VGND VPWR VPWR _1538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0771_ _1560_/Q _1598_/Q VGND VGND VPWR VPWR _0771_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0840_ _1549_/Q _0743_/Y _0829_/B _1563_/Q _0833_/X VGND VGND VPWR VPWR _0841_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1254_ hold34/X _1218_/Y _1253_/X _1009_/A VGND VGND VPWR VPWR _1464_/D sky130_fd_sc_hd__o211a_1
X_1185_ _1484_/Q _1126_/B _1183_/Y _1184_/X _0867_/A VGND VGND VPWR VPWR _1484_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_19_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1427__121 clkload5/A VGND VGND VPWR VPWR _1579_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ hold23/A hold8/A _0993_/A VGND VGND VPWR VPWR _0989_/A sky130_fd_sc_hd__and3_1
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1354__48 _1312__6/A VGND VGND VPWR VPWR _1506_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0823_ _0912_/A1 _1589_/Q _0813_/Y _0813_/B _1169_/B VGND VGND VPWR VPWR _0824_/B
+ sky130_fd_sc_hd__a32o_1
X_0754_ _1490_/Q _1489_/Q hold43/A VGND VGND VPWR VPWR _0854_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1306_ _1306_/A _1306_/B VGND VGND VPWR VPWR _1306_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1237_ hold35/A hold40/A _1282_/S VGND VGND VPWR VPWR _1237_/X sky130_fd_sc_hd__mux2_1
X_1099_ _1087_/Y _1098_/X _1097_/X _1288_/C1 VGND VGND VPWR VPWR _1504_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1168_ _1168_/A _1182_/A _1182_/B VGND VGND VPWR VPWR _1168_/X sky130_fd_sc_hd__and3_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _1105_/A _1105_/D VGND VGND VPWR VPWR _1120_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0806_ _0912_/A1 _1597_/Q _0792_/Y _0792_/A _1063_/A1 VGND VGND VPWR VPWR _0807_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0737_ hold15/X VGND VGND VPWR VPWR _1109_/A sky130_fd_sc_hd__inv_2
XFILLER_0_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1324__18 _1315__9/A VGND VGND VPWR VPWR _1467_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1571_ _1571_/CLK _1571_/D VGND VGND VPWR VPWR _1571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1005_ _1071_/A _1289_/C VGND VGND VPWR VPWR _1005_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1485_ _1485_/CLK _1485_/D VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfxtp_2
X_1554_ _1554_/CLK _1554_/D VGND VGND VPWR VPWR _1554_/Q sky130_fd_sc_hd__dfxtp_1
.ends

