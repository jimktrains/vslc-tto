VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.720 BY 13.720 ;
  OBS
      LAYER met1 ;
        RECT 0.000 13.440 13.720 13.720 ;
        RECT 0.000 12.880 1.680 13.440 ;
      LAYER met1 ;
        RECT 1.680 12.880 3.080 13.440 ;
      LAYER met1 ;
        RECT 3.080 12.880 4.480 13.440 ;
      LAYER met1 ;
        RECT 4.480 12.880 5.320 13.440 ;
      LAYER met1 ;
        RECT 5.320 12.880 6.720 13.440 ;
      LAYER met1 ;
        RECT 6.720 12.880 8.120 13.440 ;
      LAYER met1 ;
        RECT 8.120 12.880 8.960 13.440 ;
        RECT 0.000 12.320 1.400 12.880 ;
      LAYER met1 ;
        RECT 1.400 12.600 3.360 12.880 ;
        RECT 1.400 12.320 1.960 12.600 ;
      LAYER met1 ;
        RECT 1.960 12.320 2.520 12.600 ;
        RECT 0.000 11.760 2.520 12.320 ;
      LAYER met1 ;
        RECT 2.520 11.760 3.360 12.600 ;
      LAYER met1 ;
        RECT 3.360 12.320 4.200 12.880 ;
      LAYER met1 ;
        RECT 4.200 12.600 5.600 12.880 ;
      LAYER met1 ;
        RECT 5.600 12.600 6.440 12.880 ;
      LAYER met1 ;
        RECT 6.440 12.600 8.400 12.880 ;
        RECT 4.200 12.320 4.760 12.600 ;
      LAYER met1 ;
        RECT 3.360 11.760 3.920 12.320 ;
        RECT 0.000 11.480 2.240 11.760 ;
      LAYER met1 ;
        RECT 2.240 11.480 3.080 11.760 ;
      LAYER met1 ;
        RECT 0.000 10.920 1.960 11.480 ;
      LAYER met1 ;
        RECT 1.960 11.200 3.080 11.480 ;
      LAYER met1 ;
        RECT 3.080 11.200 3.920 11.760 ;
      LAYER met1 ;
        RECT 1.960 10.920 2.800 11.200 ;
      LAYER met1 ;
        RECT 2.800 10.920 3.920 11.200 ;
      LAYER met1 ;
        RECT 3.920 10.920 4.760 12.320 ;
      LAYER met1 ;
        RECT 0.000 10.360 1.680 10.920 ;
      LAYER met1 ;
        RECT 1.680 10.360 2.520 10.920 ;
      LAYER met1 ;
        RECT 2.520 10.640 4.200 10.920 ;
      LAYER met1 ;
        RECT 4.200 10.640 4.760 10.920 ;
      LAYER met1 ;
        RECT 4.760 10.640 5.040 12.600 ;
      LAYER met1 ;
        RECT 5.040 10.640 5.880 12.600 ;
      LAYER met1 ;
        RECT 5.880 12.320 6.440 12.600 ;
      LAYER met1 ;
        RECT 6.440 12.320 7.000 12.600 ;
      LAYER met1 ;
        RECT 7.000 12.320 7.560 12.600 ;
        RECT 5.880 11.760 7.560 12.320 ;
      LAYER met1 ;
        RECT 7.560 11.760 8.400 12.600 ;
      LAYER met1 ;
        RECT 8.400 11.760 8.960 12.880 ;
      LAYER met1 ;
        RECT 8.960 12.600 10.920 13.440 ;
      LAYER met1 ;
        RECT 10.920 12.600 13.720 13.440 ;
      LAYER met1 ;
        RECT 8.960 12.320 9.800 12.600 ;
      LAYER met1 ;
        RECT 9.800 12.320 13.720 12.600 ;
      LAYER met1 ;
        RECT 8.960 12.040 10.640 12.320 ;
      LAYER met1 ;
        RECT 10.640 12.040 13.720 12.320 ;
        RECT 5.880 11.480 7.280 11.760 ;
      LAYER met1 ;
        RECT 7.280 11.480 8.120 11.760 ;
      LAYER met1 ;
        RECT 5.880 10.920 7.000 11.480 ;
      LAYER met1 ;
        RECT 7.000 11.200 8.120 11.480 ;
      LAYER met1 ;
        RECT 8.120 11.200 8.960 11.760 ;
      LAYER met1 ;
        RECT 8.960 11.480 10.920 12.040 ;
        RECT 8.960 11.200 9.800 11.480 ;
      LAYER met1 ;
        RECT 9.800 11.200 10.080 11.480 ;
      LAYER met1 ;
        RECT 10.080 11.200 10.920 11.480 ;
        RECT 7.000 10.920 7.840 11.200 ;
      LAYER met1 ;
        RECT 7.840 10.920 10.360 11.200 ;
      LAYER met1 ;
        RECT 10.360 10.920 10.920 11.200 ;
      LAYER met1 ;
        RECT 5.880 10.640 6.720 10.920 ;
        RECT 2.520 10.360 2.800 10.640 ;
      LAYER met1 ;
        RECT 2.800 10.360 3.360 10.640 ;
      LAYER met1 ;
        RECT 3.360 10.360 4.200 10.640 ;
      LAYER met1 ;
        RECT 4.200 10.360 5.600 10.640 ;
      LAYER met1 ;
        RECT 5.600 10.360 6.720 10.640 ;
      LAYER met1 ;
        RECT 6.720 10.360 7.560 10.920 ;
      LAYER met1 ;
        RECT 7.560 10.640 8.960 10.920 ;
      LAYER met1 ;
        RECT 8.960 10.640 9.520 10.920 ;
      LAYER met1 ;
        RECT 9.520 10.640 10.080 10.920 ;
        RECT 7.560 10.360 7.840 10.640 ;
      LAYER met1 ;
        RECT 7.840 10.360 8.400 10.640 ;
      LAYER met1 ;
        RECT 8.400 10.360 8.960 10.640 ;
      LAYER met1 ;
        RECT 8.960 10.360 9.800 10.640 ;
      LAYER met1 ;
        RECT 9.800 10.360 10.080 10.640 ;
      LAYER met1 ;
        RECT 10.080 10.360 10.920 10.920 ;
      LAYER met1 ;
        RECT 10.920 10.360 13.720 12.040 ;
        RECT 0.000 9.800 1.400 10.360 ;
      LAYER met1 ;
        RECT 1.400 9.800 3.360 10.360 ;
      LAYER met1 ;
        RECT 3.360 9.800 4.480 10.360 ;
      LAYER met1 ;
        RECT 4.480 10.080 5.600 10.360 ;
      LAYER met1 ;
        RECT 5.600 10.080 6.440 10.360 ;
      LAYER met1 ;
        RECT 4.480 9.800 5.320 10.080 ;
      LAYER met1 ;
        RECT 5.320 9.800 6.440 10.080 ;
      LAYER met1 ;
        RECT 6.440 9.800 8.400 10.360 ;
      LAYER met1 ;
        RECT 8.400 9.800 9.240 10.360 ;
      LAYER met1 ;
        RECT 9.240 9.800 10.640 10.360 ;
      LAYER met1 ;
        RECT 10.640 9.800 13.720 10.360 ;
        RECT 0.000 9.520 13.720 9.800 ;
        RECT 0.000 8.680 1.120 9.520 ;
      LAYER met1 ;
        RECT 1.120 8.680 3.360 9.520 ;
      LAYER met1 ;
        RECT 3.360 9.240 4.480 9.520 ;
      LAYER met1 ;
        RECT 4.480 9.240 7.000 9.520 ;
      LAYER met1 ;
        RECT 3.360 8.680 4.200 9.240 ;
      LAYER met1 ;
        RECT 4.200 8.680 7.000 9.240 ;
      LAYER met1 ;
        RECT 7.000 8.680 7.560 9.520 ;
        RECT 0.000 8.400 1.400 8.680 ;
      LAYER met1 ;
        RECT 1.400 8.400 3.360 8.680 ;
      LAYER met1 ;
        RECT 3.360 8.400 3.920 8.680 ;
      LAYER met1 ;
        RECT 3.920 8.400 5.320 8.680 ;
      LAYER met1 ;
        RECT 5.320 8.400 6.160 8.680 ;
        RECT 0.000 5.880 1.680 8.400 ;
        RECT 0.000 5.040 0.280 5.880 ;
      LAYER met1 ;
        RECT 0.280 5.320 1.400 5.880 ;
      LAYER met1 ;
        RECT 1.400 5.320 1.680 5.880 ;
      LAYER met1 ;
        RECT 1.680 5.320 2.800 8.400 ;
      LAYER met1 ;
        RECT 2.800 7.280 3.920 8.400 ;
      LAYER met1 ;
        RECT 3.920 7.560 5.040 8.400 ;
      LAYER met1 ;
        RECT 5.040 7.840 6.160 8.400 ;
      LAYER met1 ;
        RECT 6.160 7.840 7.280 8.680 ;
      LAYER met1 ;
        RECT 7.280 7.840 7.560 8.680 ;
        RECT 5.040 7.560 7.560 7.840 ;
      LAYER met1 ;
        RECT 3.920 7.280 5.320 7.560 ;
      LAYER met1 ;
        RECT 5.320 7.280 6.160 7.560 ;
      LAYER met1 ;
        RECT 6.160 7.280 6.720 7.560 ;
      LAYER met1 ;
        RECT 6.720 7.280 7.560 7.560 ;
      LAYER met1 ;
        RECT 7.560 7.280 8.680 9.520 ;
      LAYER met1 ;
        RECT 8.680 8.960 9.800 9.520 ;
      LAYER met1 ;
        RECT 9.800 8.960 10.920 9.520 ;
      LAYER met1 ;
        RECT 8.680 8.120 9.520 8.960 ;
      LAYER met1 ;
        RECT 9.520 8.680 10.920 8.960 ;
      LAYER met1 ;
        RECT 10.920 8.680 13.720 9.520 ;
      LAYER met1 ;
        RECT 9.520 8.120 10.640 8.680 ;
      LAYER met1 ;
        RECT 8.680 7.280 8.960 8.120 ;
      LAYER met1 ;
        RECT 8.960 7.840 10.640 8.120 ;
      LAYER met1 ;
        RECT 10.640 7.840 13.720 8.680 ;
      LAYER met1 ;
        RECT 8.960 7.280 10.080 7.840 ;
      LAYER met1 ;
        RECT 2.800 6.720 4.200 7.280 ;
      LAYER met1 ;
        RECT 4.200 6.720 7.000 7.280 ;
      LAYER met1 ;
        RECT 7.000 6.720 7.560 7.280 ;
      LAYER met1 ;
        RECT 7.560 7.000 10.080 7.280 ;
      LAYER met1 ;
        RECT 10.080 7.000 13.720 7.840 ;
      LAYER met1 ;
        RECT 7.560 6.720 9.520 7.000 ;
      LAYER met1 ;
        RECT 9.520 6.720 13.720 7.000 ;
        RECT 2.800 6.440 4.480 6.720 ;
      LAYER met1 ;
        RECT 4.480 6.440 7.280 6.720 ;
      LAYER met1 ;
        RECT 2.800 5.880 6.160 6.440 ;
      LAYER met1 ;
        RECT 0.280 5.040 2.800 5.320 ;
      LAYER met1 ;
        RECT 2.800 5.040 3.920 5.880 ;
      LAYER met1 ;
        RECT 3.920 5.320 5.040 5.880 ;
      LAYER met1 ;
        RECT 5.040 5.320 6.160 5.880 ;
      LAYER met1 ;
        RECT 6.160 5.320 7.280 6.440 ;
        RECT 3.920 5.040 7.280 5.320 ;
      LAYER met1 ;
        RECT 7.280 5.040 7.560 6.720 ;
      LAYER met1 ;
        RECT 7.560 6.440 10.080 6.720 ;
      LAYER met1 ;
        RECT 0.000 4.480 0.560 5.040 ;
      LAYER met1 ;
        RECT 0.560 4.480 2.520 5.040 ;
      LAYER met1 ;
        RECT 2.520 4.480 4.200 5.040 ;
      LAYER met1 ;
        RECT 4.200 4.480 7.000 5.040 ;
      LAYER met1 ;
        RECT 0.000 4.200 0.840 4.480 ;
      LAYER met1 ;
        RECT 0.840 4.200 2.520 4.480 ;
      LAYER met1 ;
        RECT 2.520 4.200 4.480 4.480 ;
      LAYER met1 ;
        RECT 4.480 4.200 7.000 4.480 ;
      LAYER met1 ;
        RECT 7.000 4.200 7.560 5.040 ;
      LAYER met1 ;
        RECT 7.560 4.200 8.680 6.440 ;
      LAYER met1 ;
        RECT 8.680 5.600 8.960 6.440 ;
      LAYER met1 ;
        RECT 8.960 5.880 10.080 6.440 ;
      LAYER met1 ;
        RECT 10.080 5.880 13.720 6.720 ;
      LAYER met1 ;
        RECT 8.960 5.600 10.640 5.880 ;
      LAYER met1 ;
        RECT 8.680 5.040 9.520 5.600 ;
      LAYER met1 ;
        RECT 9.520 5.320 10.640 5.600 ;
      LAYER met1 ;
        RECT 10.640 5.320 13.720 5.880 ;
      LAYER met1 ;
        RECT 9.520 5.040 10.920 5.320 ;
      LAYER met1 ;
        RECT 8.680 4.200 9.800 5.040 ;
      LAYER met1 ;
        RECT 9.800 4.200 10.920 5.040 ;
      LAYER met1 ;
        RECT 10.920 4.200 13.720 5.320 ;
        RECT 0.000 3.920 13.720 4.200 ;
        RECT 0.000 3.080 1.120 3.920 ;
      LAYER met1 ;
        RECT 1.120 3.640 3.080 3.920 ;
      LAYER met1 ;
        RECT 3.080 3.640 3.640 3.920 ;
      LAYER met1 ;
        RECT 3.640 3.640 5.600 3.920 ;
      LAYER met1 ;
        RECT 5.600 3.640 7.000 3.920 ;
      LAYER met1 ;
        RECT 7.000 3.640 7.560 3.920 ;
        RECT 1.120 3.360 3.360 3.640 ;
      LAYER met1 ;
        RECT 3.360 3.360 3.640 3.640 ;
      LAYER met1 ;
        RECT 3.640 3.360 5.880 3.640 ;
      LAYER met1 ;
        RECT 5.880 3.360 6.720 3.640 ;
      LAYER met1 ;
        RECT 6.720 3.360 7.560 3.640 ;
      LAYER met1 ;
        RECT 7.560 3.360 9.240 3.920 ;
      LAYER met1 ;
        RECT 9.240 3.360 10.080 3.920 ;
      LAYER met1 ;
        RECT 10.080 3.360 13.720 3.920 ;
      LAYER met1 ;
        RECT 1.120 3.080 3.080 3.360 ;
      LAYER met1 ;
        RECT 3.080 3.080 3.640 3.360 ;
      LAYER met1 ;
        RECT 3.640 3.080 5.600 3.360 ;
      LAYER met1 ;
        RECT 5.600 3.080 6.440 3.360 ;
        RECT 0.000 0.280 1.680 3.080 ;
      LAYER met1 ;
        RECT 1.680 0.280 2.520 3.080 ;
      LAYER met1 ;
        RECT 2.520 0.280 4.200 3.080 ;
      LAYER met1 ;
        RECT 4.200 0.280 5.040 3.080 ;
      LAYER met1 ;
        RECT 5.040 2.800 6.440 3.080 ;
      LAYER met1 ;
        RECT 6.440 2.800 7.560 3.360 ;
      LAYER met1 ;
        RECT 7.560 2.800 8.960 3.360 ;
      LAYER met1 ;
        RECT 8.960 3.080 10.360 3.360 ;
      LAYER met1 ;
        RECT 10.360 3.080 13.720 3.360 ;
      LAYER met1 ;
        RECT 8.960 2.800 9.520 3.080 ;
      LAYER met1 ;
        RECT 5.040 1.120 6.720 2.800 ;
      LAYER met1 ;
        RECT 6.720 1.120 7.560 2.800 ;
      LAYER met1 ;
        RECT 7.560 1.400 8.680 2.800 ;
      LAYER met1 ;
        RECT 8.680 1.400 9.520 2.800 ;
      LAYER met1 ;
        RECT 7.560 1.120 8.960 1.400 ;
      LAYER met1 ;
        RECT 8.960 1.120 9.520 1.400 ;
      LAYER met1 ;
        RECT 9.520 1.120 9.800 3.080 ;
      LAYER met1 ;
        RECT 9.800 1.120 10.640 3.080 ;
      LAYER met1 ;
        RECT 10.640 1.120 13.720 3.080 ;
        RECT 5.040 0.280 6.440 1.120 ;
      LAYER met1 ;
        RECT 6.440 0.840 7.840 1.120 ;
      LAYER met1 ;
        RECT 7.840 0.840 8.960 1.120 ;
      LAYER met1 ;
        RECT 8.960 0.840 10.360 1.120 ;
        RECT 6.440 0.280 8.120 0.840 ;
      LAYER met1 ;
        RECT 8.120 0.280 9.240 0.840 ;
      LAYER met1 ;
        RECT 9.240 0.560 10.360 0.840 ;
      LAYER met1 ;
        RECT 10.360 0.560 13.720 1.120 ;
      LAYER met1 ;
        RECT 9.240 0.280 10.080 0.560 ;
      LAYER met1 ;
        RECT 10.080 0.280 13.720 0.560 ;
        RECT 0.000 0.000 13.720 0.280 ;
      LAYER met2 ;
        RECT 0.000 13.440 13.720 13.720 ;
        RECT 0.000 12.880 1.680 13.440 ;
      LAYER met2 ;
        RECT 1.680 12.880 3.080 13.440 ;
      LAYER met2 ;
        RECT 3.080 12.880 4.480 13.440 ;
      LAYER met2 ;
        RECT 4.480 12.880 5.320 13.440 ;
      LAYER met2 ;
        RECT 5.320 12.880 6.720 13.440 ;
      LAYER met2 ;
        RECT 6.720 12.880 8.120 13.440 ;
      LAYER met2 ;
        RECT 8.120 12.880 8.960 13.440 ;
        RECT 0.000 12.320 1.400 12.880 ;
      LAYER met2 ;
        RECT 1.400 12.600 3.360 12.880 ;
        RECT 1.400 12.320 1.960 12.600 ;
      LAYER met2 ;
        RECT 1.960 12.320 2.520 12.600 ;
        RECT 0.000 11.760 2.520 12.320 ;
      LAYER met2 ;
        RECT 2.520 11.760 3.360 12.600 ;
      LAYER met2 ;
        RECT 3.360 12.320 4.200 12.880 ;
      LAYER met2 ;
        RECT 4.200 12.600 5.600 12.880 ;
      LAYER met2 ;
        RECT 5.600 12.600 6.440 12.880 ;
      LAYER met2 ;
        RECT 6.440 12.600 8.400 12.880 ;
        RECT 4.200 12.320 4.760 12.600 ;
      LAYER met2 ;
        RECT 3.360 11.760 3.920 12.320 ;
        RECT 0.000 11.480 2.240 11.760 ;
      LAYER met2 ;
        RECT 2.240 11.480 3.080 11.760 ;
      LAYER met2 ;
        RECT 0.000 10.920 1.960 11.480 ;
      LAYER met2 ;
        RECT 1.960 11.200 3.080 11.480 ;
      LAYER met2 ;
        RECT 3.080 11.200 3.920 11.760 ;
      LAYER met2 ;
        RECT 1.960 10.920 2.800 11.200 ;
      LAYER met2 ;
        RECT 2.800 10.920 3.920 11.200 ;
      LAYER met2 ;
        RECT 3.920 10.920 4.760 12.320 ;
      LAYER met2 ;
        RECT 0.000 10.360 1.680 10.920 ;
      LAYER met2 ;
        RECT 1.680 10.360 2.520 10.920 ;
      LAYER met2 ;
        RECT 2.520 10.640 4.200 10.920 ;
      LAYER met2 ;
        RECT 4.200 10.640 4.760 10.920 ;
      LAYER met2 ;
        RECT 4.760 10.640 5.040 12.600 ;
      LAYER met2 ;
        RECT 5.040 10.640 5.880 12.600 ;
      LAYER met2 ;
        RECT 5.880 12.320 6.440 12.600 ;
      LAYER met2 ;
        RECT 6.440 12.320 7.000 12.600 ;
      LAYER met2 ;
        RECT 7.000 12.320 7.560 12.600 ;
        RECT 5.880 11.760 7.560 12.320 ;
      LAYER met2 ;
        RECT 7.560 11.760 8.400 12.600 ;
      LAYER met2 ;
        RECT 8.400 11.760 8.960 12.880 ;
      LAYER met2 ;
        RECT 8.960 12.600 10.920 13.440 ;
      LAYER met2 ;
        RECT 10.920 12.600 13.720 13.440 ;
      LAYER met2 ;
        RECT 8.960 12.320 9.800 12.600 ;
      LAYER met2 ;
        RECT 9.800 12.320 13.720 12.600 ;
      LAYER met2 ;
        RECT 8.960 12.040 10.640 12.320 ;
      LAYER met2 ;
        RECT 10.640 12.040 13.720 12.320 ;
        RECT 5.880 11.480 7.280 11.760 ;
      LAYER met2 ;
        RECT 7.280 11.480 8.120 11.760 ;
      LAYER met2 ;
        RECT 5.880 10.920 7.000 11.480 ;
      LAYER met2 ;
        RECT 7.000 11.200 8.120 11.480 ;
      LAYER met2 ;
        RECT 8.120 11.200 8.960 11.760 ;
      LAYER met2 ;
        RECT 8.960 11.480 10.920 12.040 ;
        RECT 8.960 11.200 9.800 11.480 ;
      LAYER met2 ;
        RECT 9.800 11.200 10.080 11.480 ;
      LAYER met2 ;
        RECT 10.080 11.200 10.920 11.480 ;
        RECT 7.000 10.920 7.840 11.200 ;
      LAYER met2 ;
        RECT 7.840 10.920 10.360 11.200 ;
      LAYER met2 ;
        RECT 10.360 10.920 10.920 11.200 ;
      LAYER met2 ;
        RECT 5.880 10.640 6.720 10.920 ;
        RECT 2.520 10.360 2.800 10.640 ;
      LAYER met2 ;
        RECT 2.800 10.360 3.360 10.640 ;
      LAYER met2 ;
        RECT 3.360 10.360 4.200 10.640 ;
      LAYER met2 ;
        RECT 4.200 10.360 5.600 10.640 ;
      LAYER met2 ;
        RECT 5.600 10.360 6.720 10.640 ;
      LAYER met2 ;
        RECT 6.720 10.360 7.560 10.920 ;
      LAYER met2 ;
        RECT 7.560 10.640 8.960 10.920 ;
      LAYER met2 ;
        RECT 8.960 10.640 9.520 10.920 ;
      LAYER met2 ;
        RECT 9.520 10.640 10.080 10.920 ;
        RECT 7.560 10.360 7.840 10.640 ;
      LAYER met2 ;
        RECT 7.840 10.360 8.400 10.640 ;
      LAYER met2 ;
        RECT 8.400 10.360 8.960 10.640 ;
      LAYER met2 ;
        RECT 8.960 10.360 9.800 10.640 ;
      LAYER met2 ;
        RECT 9.800 10.360 10.080 10.640 ;
      LAYER met2 ;
        RECT 10.080 10.360 10.920 10.920 ;
      LAYER met2 ;
        RECT 10.920 10.360 13.720 12.040 ;
        RECT 0.000 9.800 1.400 10.360 ;
      LAYER met2 ;
        RECT 1.400 9.800 3.360 10.360 ;
      LAYER met2 ;
        RECT 3.360 9.800 4.480 10.360 ;
      LAYER met2 ;
        RECT 4.480 10.080 5.600 10.360 ;
      LAYER met2 ;
        RECT 5.600 10.080 6.440 10.360 ;
      LAYER met2 ;
        RECT 4.480 9.800 5.320 10.080 ;
      LAYER met2 ;
        RECT 5.320 9.800 6.440 10.080 ;
      LAYER met2 ;
        RECT 6.440 9.800 8.400 10.360 ;
      LAYER met2 ;
        RECT 8.400 9.800 9.240 10.360 ;
      LAYER met2 ;
        RECT 9.240 9.800 10.640 10.360 ;
      LAYER met2 ;
        RECT 10.640 9.800 13.720 10.360 ;
        RECT 0.000 9.520 13.720 9.800 ;
        RECT 0.000 8.680 1.120 9.520 ;
      LAYER met2 ;
        RECT 1.120 8.680 3.360 9.520 ;
      LAYER met2 ;
        RECT 3.360 9.240 4.480 9.520 ;
      LAYER met2 ;
        RECT 4.480 9.240 7.000 9.520 ;
      LAYER met2 ;
        RECT 3.360 8.680 4.200 9.240 ;
      LAYER met2 ;
        RECT 4.200 8.680 7.000 9.240 ;
      LAYER met2 ;
        RECT 7.000 8.680 7.560 9.520 ;
        RECT 0.000 8.400 1.400 8.680 ;
      LAYER met2 ;
        RECT 1.400 8.400 3.360 8.680 ;
      LAYER met2 ;
        RECT 3.360 8.400 3.920 8.680 ;
      LAYER met2 ;
        RECT 3.920 8.400 5.320 8.680 ;
      LAYER met2 ;
        RECT 5.320 8.400 6.160 8.680 ;
        RECT 0.000 5.880 1.680 8.400 ;
        RECT 0.000 5.040 0.280 5.880 ;
      LAYER met2 ;
        RECT 0.280 5.320 1.400 5.880 ;
      LAYER met2 ;
        RECT 1.400 5.320 1.680 5.880 ;
      LAYER met2 ;
        RECT 1.680 5.320 2.800 8.400 ;
      LAYER met2 ;
        RECT 2.800 7.280 3.920 8.400 ;
      LAYER met2 ;
        RECT 3.920 7.560 5.040 8.400 ;
      LAYER met2 ;
        RECT 5.040 7.840 6.160 8.400 ;
      LAYER met2 ;
        RECT 6.160 7.840 7.280 8.680 ;
      LAYER met2 ;
        RECT 7.280 7.840 7.560 8.680 ;
        RECT 5.040 7.560 7.560 7.840 ;
      LAYER met2 ;
        RECT 3.920 7.280 5.320 7.560 ;
      LAYER met2 ;
        RECT 5.320 7.280 6.160 7.560 ;
      LAYER met2 ;
        RECT 6.160 7.280 6.720 7.560 ;
      LAYER met2 ;
        RECT 6.720 7.280 7.560 7.560 ;
      LAYER met2 ;
        RECT 7.560 7.280 8.680 9.520 ;
      LAYER met2 ;
        RECT 8.680 8.960 9.800 9.520 ;
      LAYER met2 ;
        RECT 9.800 8.960 10.920 9.520 ;
      LAYER met2 ;
        RECT 8.680 8.120 9.520 8.960 ;
      LAYER met2 ;
        RECT 9.520 8.680 10.920 8.960 ;
      LAYER met2 ;
        RECT 10.920 8.680 13.720 9.520 ;
      LAYER met2 ;
        RECT 9.520 8.120 10.640 8.680 ;
      LAYER met2 ;
        RECT 8.680 7.280 8.960 8.120 ;
      LAYER met2 ;
        RECT 8.960 7.840 10.640 8.120 ;
      LAYER met2 ;
        RECT 10.640 7.840 13.720 8.680 ;
      LAYER met2 ;
        RECT 8.960 7.280 10.080 7.840 ;
      LAYER met2 ;
        RECT 2.800 6.720 4.200 7.280 ;
      LAYER met2 ;
        RECT 4.200 6.720 7.000 7.280 ;
      LAYER met2 ;
        RECT 7.000 6.720 7.560 7.280 ;
      LAYER met2 ;
        RECT 7.560 7.000 10.080 7.280 ;
      LAYER met2 ;
        RECT 10.080 7.000 13.720 7.840 ;
      LAYER met2 ;
        RECT 7.560 6.720 9.520 7.000 ;
      LAYER met2 ;
        RECT 9.520 6.720 13.720 7.000 ;
        RECT 2.800 6.440 4.480 6.720 ;
      LAYER met2 ;
        RECT 4.480 6.440 7.280 6.720 ;
      LAYER met2 ;
        RECT 2.800 5.880 6.160 6.440 ;
      LAYER met2 ;
        RECT 0.280 5.040 2.800 5.320 ;
      LAYER met2 ;
        RECT 2.800 5.040 3.920 5.880 ;
      LAYER met2 ;
        RECT 3.920 5.320 5.040 5.880 ;
      LAYER met2 ;
        RECT 5.040 5.320 6.160 5.880 ;
      LAYER met2 ;
        RECT 6.160 5.320 7.280 6.440 ;
        RECT 3.920 5.040 7.280 5.320 ;
      LAYER met2 ;
        RECT 7.280 5.040 7.560 6.720 ;
      LAYER met2 ;
        RECT 7.560 6.440 10.080 6.720 ;
      LAYER met2 ;
        RECT 0.000 4.480 0.560 5.040 ;
      LAYER met2 ;
        RECT 0.560 4.480 2.520 5.040 ;
      LAYER met2 ;
        RECT 2.520 4.480 4.200 5.040 ;
      LAYER met2 ;
        RECT 4.200 4.480 7.000 5.040 ;
      LAYER met2 ;
        RECT 0.000 4.200 0.840 4.480 ;
      LAYER met2 ;
        RECT 0.840 4.200 2.520 4.480 ;
      LAYER met2 ;
        RECT 2.520 4.200 4.480 4.480 ;
      LAYER met2 ;
        RECT 4.480 4.200 7.000 4.480 ;
      LAYER met2 ;
        RECT 7.000 4.200 7.560 5.040 ;
      LAYER met2 ;
        RECT 7.560 4.200 8.680 6.440 ;
      LAYER met2 ;
        RECT 8.680 5.600 8.960 6.440 ;
      LAYER met2 ;
        RECT 8.960 5.880 10.080 6.440 ;
      LAYER met2 ;
        RECT 10.080 5.880 13.720 6.720 ;
      LAYER met2 ;
        RECT 8.960 5.600 10.640 5.880 ;
      LAYER met2 ;
        RECT 8.680 5.040 9.520 5.600 ;
      LAYER met2 ;
        RECT 9.520 5.320 10.640 5.600 ;
      LAYER met2 ;
        RECT 10.640 5.320 13.720 5.880 ;
      LAYER met2 ;
        RECT 9.520 5.040 10.920 5.320 ;
      LAYER met2 ;
        RECT 8.680 4.200 9.800 5.040 ;
      LAYER met2 ;
        RECT 9.800 4.200 10.920 5.040 ;
      LAYER met2 ;
        RECT 10.920 4.200 13.720 5.320 ;
        RECT 0.000 3.920 13.720 4.200 ;
        RECT 0.000 3.080 1.120 3.920 ;
      LAYER met2 ;
        RECT 1.120 3.640 3.080 3.920 ;
      LAYER met2 ;
        RECT 3.080 3.640 3.640 3.920 ;
      LAYER met2 ;
        RECT 3.640 3.640 5.600 3.920 ;
      LAYER met2 ;
        RECT 5.600 3.640 7.000 3.920 ;
      LAYER met2 ;
        RECT 7.000 3.640 7.560 3.920 ;
        RECT 1.120 3.360 3.360 3.640 ;
      LAYER met2 ;
        RECT 3.360 3.360 3.640 3.640 ;
      LAYER met2 ;
        RECT 3.640 3.360 5.880 3.640 ;
      LAYER met2 ;
        RECT 5.880 3.360 6.720 3.640 ;
      LAYER met2 ;
        RECT 6.720 3.360 7.560 3.640 ;
      LAYER met2 ;
        RECT 7.560 3.360 9.240 3.920 ;
      LAYER met2 ;
        RECT 9.240 3.360 10.080 3.920 ;
      LAYER met2 ;
        RECT 10.080 3.360 13.720 3.920 ;
      LAYER met2 ;
        RECT 1.120 3.080 3.080 3.360 ;
      LAYER met2 ;
        RECT 3.080 3.080 3.640 3.360 ;
      LAYER met2 ;
        RECT 3.640 3.080 5.600 3.360 ;
      LAYER met2 ;
        RECT 5.600 3.080 6.440 3.360 ;
        RECT 0.000 0.280 1.680 3.080 ;
      LAYER met2 ;
        RECT 1.680 0.280 2.520 3.080 ;
      LAYER met2 ;
        RECT 2.520 0.280 4.200 3.080 ;
      LAYER met2 ;
        RECT 4.200 0.280 5.040 3.080 ;
      LAYER met2 ;
        RECT 5.040 2.800 6.440 3.080 ;
      LAYER met2 ;
        RECT 6.440 2.800 7.560 3.360 ;
      LAYER met2 ;
        RECT 7.560 2.800 8.960 3.360 ;
      LAYER met2 ;
        RECT 8.960 3.080 10.360 3.360 ;
      LAYER met2 ;
        RECT 10.360 3.080 13.720 3.360 ;
      LAYER met2 ;
        RECT 8.960 2.800 9.520 3.080 ;
      LAYER met2 ;
        RECT 5.040 1.120 6.720 2.800 ;
      LAYER met2 ;
        RECT 6.720 1.120 7.560 2.800 ;
      LAYER met2 ;
        RECT 7.560 1.400 8.680 2.800 ;
      LAYER met2 ;
        RECT 8.680 1.400 9.520 2.800 ;
      LAYER met2 ;
        RECT 7.560 1.120 8.960 1.400 ;
      LAYER met2 ;
        RECT 8.960 1.120 9.520 1.400 ;
      LAYER met2 ;
        RECT 9.520 1.120 9.800 3.080 ;
      LAYER met2 ;
        RECT 9.800 1.120 10.640 3.080 ;
      LAYER met2 ;
        RECT 10.640 1.120 13.720 3.080 ;
        RECT 5.040 0.280 6.440 1.120 ;
      LAYER met2 ;
        RECT 6.440 0.840 7.840 1.120 ;
      LAYER met2 ;
        RECT 7.840 0.840 8.960 1.120 ;
      LAYER met2 ;
        RECT 8.960 0.840 10.360 1.120 ;
        RECT 6.440 0.280 8.120 0.840 ;
      LAYER met2 ;
        RECT 8.120 0.280 9.240 0.840 ;
      LAYER met2 ;
        RECT 9.240 0.560 10.360 0.840 ;
      LAYER met2 ;
        RECT 10.360 0.560 13.720 1.120 ;
      LAYER met2 ;
        RECT 9.240 0.280 10.080 0.560 ;
      LAYER met2 ;
        RECT 10.080 0.280 13.720 0.560 ;
        RECT 0.000 0.000 13.720 0.280 ;
      LAYER met3 ;
        RECT 0.000 0.000 13.720 13.720 ;
      LAYER met4 ;
        RECT 0.000 0.000 13.720 13.720 ;
      LAYER met5 ;
        RECT 0.000 0.000 13.720 13.720 ;
  END
END my_logo
END LIBRARY

