module tt_um_jimktrains_vslc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire clknet_0_clk;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire \cur_addr[0] ;
 wire \cur_addr[1] ;
 wire \cur_addr[2] ;
 wire \cur_addr[3] ;
 wire \cur_addr[4] ;
 wire \cur_addr[5] ;
 wire \cur_addr[6] ;
 wire \cur_addr[7] ;
 wire \cycle_end_addr[0] ;
 wire \cycle_end_addr[1] ;
 wire \cycle_end_addr[2] ;
 wire \cycle_end_addr[3] ;
 wire \cycle_end_addr[4] ;
 wire \cycle_end_addr[5] ;
 wire \cycle_end_addr[6] ;
 wire \cycle_end_addr[7] ;
 wire \cycle_start_addr[0] ;
 wire \cycle_start_addr[1] ;
 wire \cycle_start_addr[2] ;
 wire \cycle_start_addr[3] ;
 wire \cycle_start_addr[4] ;
 wire \cycle_start_addr[5] ;
 wire \cycle_start_addr[6] ;
 wire \cycle_start_addr[7] ;
 wire eeprom_copi;
 wire eeprom_cs;
 wire eeprom_oe_copi;
 wire eeprom_sck;
 wire \fetch_count[0] ;
 wire \fetch_count[1] ;
 wire \fetch_count[2] ;
 wire \fetch_prev_state[0] ;
 wire \fetch_prev_state[1] ;
 wire \fetch_prev_state[2] ;
 wire \fetch_prev_state[3] ;
 wire \fetch_state[0] ;
 wire \fetch_state[1] ;
 wire \fetch_state[2] ;
 wire \fetch_state[3] ;
 wire \instr[0] ;
 wire \instr[1] ;
 wire \instr[2] ;
 wire \instr[3] ;
 wire \instr[4] ;
 wire \instr[5] ;
 wire \instr[6] ;
 wire \instr[7] ;
 wire \stack[0] ;
 wire \stack[10] ;
 wire \stack[11] ;
 wire \stack[12] ;
 wire \stack[13] ;
 wire \stack[14] ;
 wire \stack[15] ;
 wire \stack[1] ;
 wire \stack[2] ;
 wire \stack[3] ;
 wire \stack[4] ;
 wire \stack[5] ;
 wire \stack[6] ;
 wire \stack[7] ;
 wire \stack[8] ;
 wire \stack[9] ;
 wire stack_out;
 wire \timer_clock_counter[0] ;
 wire \timer_clock_counter[10] ;
 wire \timer_clock_counter[11] ;
 wire \timer_clock_counter[12] ;
 wire \timer_clock_counter[13] ;
 wire \timer_clock_counter[14] ;
 wire \timer_clock_counter[15] ;
 wire \timer_clock_counter[1] ;
 wire \timer_clock_counter[2] ;
 wire \timer_clock_counter[3] ;
 wire \timer_clock_counter[4] ;
 wire \timer_clock_counter[5] ;
 wire \timer_clock_counter[6] ;
 wire \timer_clock_counter[7] ;
 wire \timer_clock_counter[8] ;
 wire \timer_clock_counter[9] ;
 wire \timer_clock_divisor[0] ;
 wire \timer_clock_divisor[1] ;
 wire \timer_clock_divisor[2] ;
 wire \timer_clock_divisor[3] ;
 wire \timer_counter[0] ;
 wire \timer_counter[10] ;
 wire \timer_counter[11] ;
 wire \timer_counter[12] ;
 wire \timer_counter[13] ;
 wire \timer_counter[14] ;
 wire \timer_counter[15] ;
 wire \timer_counter[1] ;
 wire \timer_counter[2] ;
 wire \timer_counter[3] ;
 wire \timer_counter[4] ;
 wire \timer_counter[5] ;
 wire \timer_counter[6] ;
 wire \timer_counter[7] ;
 wire \timer_counter[8] ;
 wire \timer_counter[9] ;
 wire timer_enabled;
 wire timer_mode;
 wire timer_out;
 wire \timer_period_a[0] ;
 wire \timer_period_a[10] ;
 wire \timer_period_a[11] ;
 wire \timer_period_a[12] ;
 wire \timer_period_a[13] ;
 wire \timer_period_a[14] ;
 wire \timer_period_a[15] ;
 wire \timer_period_a[1] ;
 wire \timer_period_a[2] ;
 wire \timer_period_a[3] ;
 wire \timer_period_a[4] ;
 wire \timer_period_a[5] ;
 wire \timer_period_a[6] ;
 wire \timer_period_a[7] ;
 wire \timer_period_a[8] ;
 wire \timer_period_a[9] ;
 wire \timer_period_b[0] ;
 wire \timer_period_b[10] ;
 wire \timer_period_b[11] ;
 wire \timer_period_b[12] ;
 wire \timer_period_b[13] ;
 wire \timer_period_b[14] ;
 wire \timer_period_b[15] ;
 wire \timer_period_b[1] ;
 wire \timer_period_b[2] ;
 wire \timer_period_b[3] ;
 wire \timer_period_b[4] ;
 wire \timer_period_b[5] ;
 wire \timer_period_b[6] ;
 wire \timer_period_b[7] ;
 wire \timer_period_b[8] ;
 wire \timer_period_b[9] ;
 wire timer_phase;
 wire \ui_in_reg[0] ;
 wire \ui_in_reg[1] ;
 wire \ui_in_reg[2] ;
 wire \ui_in_reg[3] ;
 wire \ui_in_reg[4] ;
 wire \ui_in_reg[5] ;
 wire \ui_in_reg[6] ;
 wire \ui_in_reg[7] ;
 wire \uio_in_reg[3] ;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net68;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;

 sky130_fd_sc_hd__inv_2 _0725_ (.A(net52),
    .Y(_0302_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(\timer_counter[13] ),
    .Y(_0303_));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(\timer_counter[12] ),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(\timer_counter[11] ),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(\timer_counter[10] ),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(\timer_counter[9] ),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_2 _0731_ (.A(\timer_counter[8] ),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(\timer_counter[7] ),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(\timer_counter[4] ),
    .Y(_0310_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(net43),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(net45),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(net47),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(net223),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _0738_ (.A(net242),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(\cur_addr[4] ),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(\cur_addr[3] ),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(net243),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(\fetch_count[2] ),
    .Y(_0319_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(\timer_period_a[0] ),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(\timer_period_a[1] ),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(\timer_period_a[2] ),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(\timer_period_a[14] ),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _0747_ (.A(\timer_period_b[0] ),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(\timer_period_b[1] ),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(\timer_period_b[4] ),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(\timer_period_b[6] ),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(\timer_period_b[10] ),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(\timer_period_b[13] ),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _1309__3 (.A(clknet_4_13_0_clk),
    .Y(net69));
 sky130_fd_sc_hd__nand3_1 _0754_ (.A(\fetch_count[2] ),
    .B(\fetch_count[1] ),
    .C(\fetch_count[0] ),
    .Y(_0330_));
 sky130_fd_sc_hd__or3b_4 _0755_ (.A(\fetch_prev_state[2] ),
    .B(_0330_),
    .C_N(\fetch_prev_state[3] ),
    .X(_0331_));
 sky130_fd_sc_hd__nor3_4 _0756_ (.A(\fetch_prev_state[1] ),
    .B(\fetch_prev_state[0] ),
    .C(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__mux4_1 _0757_ (.A0(\timer_clock_counter[8] ),
    .A1(\timer_clock_counter[9] ),
    .A2(\timer_clock_counter[10] ),
    .A3(\timer_clock_counter[11] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0333_));
 sky130_fd_sc_hd__and2b_1 _0758_ (.A_N(\timer_clock_divisor[2] ),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__mux4_1 _0759_ (.A0(\timer_clock_counter[12] ),
    .A1(\timer_clock_counter[13] ),
    .A2(\timer_clock_counter[14] ),
    .A3(\timer_clock_counter[15] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0335_));
 sky130_fd_sc_hd__a21bo_1 _0760_ (.A1(\timer_clock_divisor[2] ),
    .A2(_0335_),
    .B1_N(\timer_clock_divisor[3] ),
    .X(_0336_));
 sky130_fd_sc_hd__mux4_1 _0761_ (.A0(\timer_clock_counter[0] ),
    .A1(\timer_clock_counter[1] ),
    .A2(\timer_clock_counter[2] ),
    .A3(\timer_clock_counter[3] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0337_));
 sky130_fd_sc_hd__mux4_1 _0762_ (.A0(\timer_clock_counter[4] ),
    .A1(\timer_clock_counter[5] ),
    .A2(\timer_clock_counter[6] ),
    .A3(\timer_clock_counter[7] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _0763_ (.A0(_0337_),
    .A1(_0338_),
    .S(\timer_clock_divisor[2] ),
    .X(_0339_));
 sky130_fd_sc_hd__o22a_1 _0764_ (.A1(_0334_),
    .A2(_0336_),
    .B1(_0339_),
    .B2(\timer_clock_divisor[3] ),
    .X(_0340_));
 sky130_fd_sc_hd__and2b_1 _0765_ (.A_N(\timer_period_b[5] ),
    .B(\timer_counter[5] ),
    .X(_0341_));
 sky130_fd_sc_hd__and2b_1 _0766_ (.A_N(\timer_period_b[12] ),
    .B(\timer_counter[12] ),
    .X(_0342_));
 sky130_fd_sc_hd__nand2b_1 _0767_ (.A_N(\timer_counter[5] ),
    .B(\timer_period_b[5] ),
    .Y(_0343_));
 sky130_fd_sc_hd__xor2_1 _0768_ (.A(\timer_counter[3] ),
    .B(\timer_period_b[3] ),
    .X(_0344_));
 sky130_fd_sc_hd__or2_1 _0769_ (.A(\timer_counter[1] ),
    .B(\timer_period_b[1] ),
    .X(_0345_));
 sky130_fd_sc_hd__nand2_1 _0770_ (.A(\timer_counter[1] ),
    .B(\timer_period_b[1] ),
    .Y(_0346_));
 sky130_fd_sc_hd__or2_1 _0771_ (.A(\timer_counter[11] ),
    .B(\timer_period_b[11] ),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_1 _0772_ (.A(\timer_counter[11] ),
    .B(\timer_period_b[11] ),
    .Y(_0348_));
 sky130_fd_sc_hd__a22o_1 _0773_ (.A1(_0304_),
    .A2(\timer_period_b[12] ),
    .B1(_0329_),
    .B2(\timer_counter[13] ),
    .X(_0349_));
 sky130_fd_sc_hd__and2b_1 _0774_ (.A_N(\timer_counter[4] ),
    .B(\timer_period_b[4] ),
    .X(_0350_));
 sky130_fd_sc_hd__and2b_1 _0775_ (.A_N(\timer_counter[10] ),
    .B(\timer_period_b[10] ),
    .X(_0351_));
 sky130_fd_sc_hd__nand2b_1 _0776_ (.A_N(\timer_counter[2] ),
    .B(\timer_period_b[2] ),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2b_1 _0777_ (.A_N(\timer_period_b[2] ),
    .B(\timer_counter[2] ),
    .Y(_0353_));
 sky130_fd_sc_hd__a2bb2o_1 _0778_ (.A1_N(\timer_counter[6] ),
    .A2_N(_0327_),
    .B1(\timer_period_b[9] ),
    .B2(_0307_),
    .X(_0354_));
 sky130_fd_sc_hd__xnor2_1 _0779_ (.A(\timer_counter[14] ),
    .B(\timer_period_b[14] ),
    .Y(_0355_));
 sky130_fd_sc_hd__o221a_1 _0780_ (.A1(_0308_),
    .A2(\timer_period_b[8] ),
    .B1(_0329_),
    .B2(\timer_counter[13] ),
    .C1(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__xnor2_1 _0781_ (.A(\timer_counter[15] ),
    .B(\timer_period_b[15] ),
    .Y(_0357_));
 sky130_fd_sc_hd__o221a_1 _0782_ (.A1(\timer_counter[0] ),
    .A2(_0324_),
    .B1(\timer_period_b[7] ),
    .B2(_0309_),
    .C1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__a221oi_1 _0783_ (.A1(_0309_),
    .A2(\timer_period_b[7] ),
    .B1(\timer_period_b[8] ),
    .B2(_0308_),
    .C1(_0342_),
    .Y(_0359_));
 sky130_fd_sc_hd__a2111o_1 _0784_ (.A1(\timer_counter[0] ),
    .A2(_0324_),
    .B1(_0341_),
    .C1(_0350_),
    .D1(_0351_),
    .X(_0360_));
 sky130_fd_sc_hd__o2111ai_1 _0785_ (.A1(_0307_),
    .A2(\timer_period_b[9] ),
    .B1(_0343_),
    .C1(_0352_),
    .D1(_0353_),
    .Y(_0361_));
 sky130_fd_sc_hd__a2111o_1 _0786_ (.A1(\timer_counter[6] ),
    .A2(_0327_),
    .B1(_0354_),
    .C1(_0360_),
    .D1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__a221o_1 _0787_ (.A1(_0345_),
    .A2(_0346_),
    .B1(_0347_),
    .B2(_0348_),
    .C1(_0344_),
    .X(_0363_));
 sky130_fd_sc_hd__a221o_1 _0788_ (.A1(\timer_counter[4] ),
    .A2(_0326_),
    .B1(_0328_),
    .B2(\timer_counter[10] ),
    .C1(_0349_),
    .X(_0364_));
 sky130_fd_sc_hd__and4_1 _0789_ (.A(timer_phase),
    .B(_0356_),
    .C(_0358_),
    .D(_0359_),
    .X(_0365_));
 sky130_fd_sc_hd__nor4b_1 _0790_ (.A(_0362_),
    .B(_0363_),
    .C(_0364_),
    .D_N(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__and3_2 _0791_ (.A(timer_mode),
    .B(_0340_),
    .C(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__nor2_2 _0792_ (.A(_0332_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__a32o_1 _0793_ (.A1(net28),
    .A2(\timer_period_b[15] ),
    .A3(_0368_),
    .B1(_0332_),
    .B2(net33),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _0794_ (.A(net49),
    .B(_0369_),
    .X(_0285_));
 sky130_fd_sc_hd__a32o_1 _0795_ (.A1(net27),
    .A2(\timer_period_b[14] ),
    .A3(_0368_),
    .B1(_0332_),
    .B2(\instr[6] ),
    .X(_0370_));
 sky130_fd_sc_hd__and2_1 _0796_ (.A(net49),
    .B(_0370_),
    .X(_0284_));
 sky130_fd_sc_hd__a32o_1 _0797_ (.A1(net27),
    .A2(\timer_period_b[13] ),
    .A3(_0368_),
    .B1(_0332_),
    .B2(net37),
    .X(_0371_));
 sky130_fd_sc_hd__and2_1 _0798_ (.A(net49),
    .B(_0371_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_2 _0799_ (.A(net49),
    .B(net38),
    .X(_0372_));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__and2_1 _0801_ (.A(net51),
    .B(net28),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _0802_ (.A(net55),
    .B(net29),
    .Y(_0375_));
 sky130_fd_sc_hd__a32o_1 _0803_ (.A1(net228),
    .A2(_0368_),
    .A3(_0374_),
    .B1(_0372_),
    .B2(_0332_),
    .X(_0282_));
 sky130_fd_sc_hd__a32o_1 _0804_ (.A1(net27),
    .A2(\timer_period_b[11] ),
    .A3(_0368_),
    .B1(_0332_),
    .B2(net41),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _0805_ (.A(net50),
    .B(_0376_),
    .X(_0281_));
 sky130_fd_sc_hd__a32o_1 _0806_ (.A1(net27),
    .A2(\timer_period_b[10] ),
    .A3(_0368_),
    .B1(_0332_),
    .B2(net44),
    .X(_0377_));
 sky130_fd_sc_hd__and2_1 _0807_ (.A(net50),
    .B(_0377_),
    .X(_0280_));
 sky130_fd_sc_hd__a32o_1 _0808_ (.A1(net27),
    .A2(\timer_period_b[9] ),
    .A3(_0368_),
    .B1(_0332_),
    .B2(net45),
    .X(_0378_));
 sky130_fd_sc_hd__and2_1 _0809_ (.A(net50),
    .B(_0378_),
    .X(_0279_));
 sky130_fd_sc_hd__a32o_1 _0810_ (.A1(net27),
    .A2(\timer_period_b[8] ),
    .A3(_0368_),
    .B1(_0332_),
    .B2(net47),
    .X(_0379_));
 sky130_fd_sc_hd__and2_1 _0811_ (.A(net50),
    .B(_0379_),
    .X(_0278_));
 sky130_fd_sc_hd__nor3b_4 _0812_ (.A(_0331_),
    .B(\fetch_prev_state[1] ),
    .C_N(\fetch_prev_state[0] ),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_2 _0813_ (.A(_0367_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__a32o_1 _0814_ (.A1(net27),
    .A2(\timer_period_b[7] ),
    .A3(_0381_),
    .B1(_0380_),
    .B2(net33),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _0815_ (.A(net49),
    .B(_0382_),
    .X(_0277_));
 sky130_fd_sc_hd__a32o_1 _0816_ (.A1(net28),
    .A2(\timer_period_b[6] ),
    .A3(_0381_),
    .B1(_0380_),
    .B2(\instr[6] ),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _0817_ (.A(net49),
    .B(_0383_),
    .X(_0276_));
 sky130_fd_sc_hd__a32o_1 _0818_ (.A1(net27),
    .A2(\timer_period_b[5] ),
    .A3(_0381_),
    .B1(_0380_),
    .B2(net37),
    .X(_0384_));
 sky130_fd_sc_hd__and2_1 _0819_ (.A(net49),
    .B(_0384_),
    .X(_0275_));
 sky130_fd_sc_hd__a32o_1 _0820_ (.A1(net241),
    .A2(_0374_),
    .A3(_0381_),
    .B1(_0380_),
    .B2(_0372_),
    .X(_0274_));
 sky130_fd_sc_hd__a32o_1 _0821_ (.A1(net27),
    .A2(\timer_period_b[3] ),
    .A3(_0381_),
    .B1(_0380_),
    .B2(net41),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _0822_ (.A(net49),
    .B(_0385_),
    .X(_0273_));
 sky130_fd_sc_hd__a32o_1 _0823_ (.A1(net27),
    .A2(\timer_period_b[2] ),
    .A3(_0381_),
    .B1(_0380_),
    .B2(net44),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _0824_ (.A(net49),
    .B(_0386_),
    .X(_0272_));
 sky130_fd_sc_hd__a32o_1 _0825_ (.A1(net28),
    .A2(_0325_),
    .A3(_0381_),
    .B1(_0380_),
    .B2(_0312_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _0826_ (.A(net49),
    .B(_0387_),
    .Y(_0271_));
 sky130_fd_sc_hd__a32o_1 _0827_ (.A1(net28),
    .A2(\timer_period_b[0] ),
    .A3(_0381_),
    .B1(_0380_),
    .B2(net47),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _0828_ (.A(net50),
    .B(_0388_),
    .X(_0270_));
 sky130_fd_sc_hd__nor2_1 _0829_ (.A(\timer_counter[14] ),
    .B(_0323_),
    .Y(_0389_));
 sky130_fd_sc_hd__xnor2_1 _0830_ (.A(\timer_counter[8] ),
    .B(\timer_period_a[8] ),
    .Y(_0390_));
 sky130_fd_sc_hd__xor2_1 _0831_ (.A(\timer_counter[6] ),
    .B(\timer_period_a[6] ),
    .X(_0391_));
 sky130_fd_sc_hd__nand2b_1 _0832_ (.A_N(\timer_counter[7] ),
    .B(\timer_period_a[7] ),
    .Y(_0392_));
 sky130_fd_sc_hd__and2b_1 _0833_ (.A_N(\timer_counter[2] ),
    .B(\timer_period_a[2] ),
    .X(_0393_));
 sky130_fd_sc_hd__xor2_1 _0834_ (.A(\timer_counter[15] ),
    .B(\timer_period_a[15] ),
    .X(_0394_));
 sky130_fd_sc_hd__a221o_1 _0835_ (.A1(_0304_),
    .A2(\timer_period_a[12] ),
    .B1(\timer_period_a[13] ),
    .B2(_0303_),
    .C1(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__a2111o_1 _0836_ (.A1(_0310_),
    .A2(\timer_period_a[4] ),
    .B1(_0389_),
    .C1(_0395_),
    .D1(timer_phase),
    .X(_0396_));
 sky130_fd_sc_hd__a221o_1 _0837_ (.A1(_0306_),
    .A2(\timer_period_a[10] ),
    .B1(\timer_period_a[11] ),
    .B2(_0305_),
    .C1(_0391_),
    .X(_0397_));
 sky130_fd_sc_hd__a2bb2o_1 _0838_ (.A1_N(\timer_counter[0] ),
    .A2_N(_0320_),
    .B1(_0322_),
    .B2(\timer_counter[2] ),
    .X(_0398_));
 sky130_fd_sc_hd__a2bb2o_1 _0839_ (.A1_N(_0309_),
    .A2_N(\timer_period_a[7] ),
    .B1(\timer_counter[1] ),
    .B2(_0321_),
    .X(_0399_));
 sky130_fd_sc_hd__a221o_1 _0840_ (.A1(\timer_counter[0] ),
    .A2(_0320_),
    .B1(_0323_),
    .B2(\timer_counter[14] ),
    .C1(_0393_),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _0841_ (.A(_0397_),
    .B(_0398_),
    .C(_0399_),
    .D(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__xnor2_1 _0842_ (.A(\timer_counter[5] ),
    .B(\timer_period_a[5] ),
    .Y(_0402_));
 sky130_fd_sc_hd__o221a_1 _0843_ (.A1(\timer_counter[1] ),
    .A2(_0321_),
    .B1(\timer_period_a[13] ),
    .B2(_0303_),
    .C1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__xor2_1 _0844_ (.A(\timer_counter[3] ),
    .B(\timer_period_a[3] ),
    .X(_0404_));
 sky130_fd_sc_hd__xor2_1 _0845_ (.A(\timer_counter[9] ),
    .B(\timer_period_a[9] ),
    .X(_0405_));
 sky130_fd_sc_hd__nor2_1 _0846_ (.A(_0404_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__o221a_1 _0847_ (.A1(_0310_),
    .A2(\timer_period_a[4] ),
    .B1(\timer_period_a[12] ),
    .B2(_0304_),
    .C1(_0390_),
    .X(_0407_));
 sky130_fd_sc_hd__o221a_1 _0848_ (.A1(_0306_),
    .A2(\timer_period_a[10] ),
    .B1(\timer_period_a[11] ),
    .B2(_0305_),
    .C1(_0392_),
    .X(_0408_));
 sky130_fd_sc_hd__nand4_1 _0849_ (.A(_0403_),
    .B(_0406_),
    .C(_0407_),
    .D(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__nor3_1 _0850_ (.A(_0396_),
    .B(_0401_),
    .C(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__o21a_1 _0851_ (.A1(_0366_),
    .A2(_0410_),
    .B1(_0340_),
    .X(_0411_));
 sky130_fd_sc_hd__a21oi_1 _0852_ (.A1(timer_phase),
    .A2(_0411_),
    .B1(_0375_),
    .Y(_0412_));
 sky130_fd_sc_hd__o21a_1 _0853_ (.A1(net231),
    .A2(_0411_),
    .B1(_0412_),
    .X(_0269_));
 sky130_fd_sc_hd__or3b_4 _0854_ (.A(_0330_),
    .B(\fetch_prev_state[3] ),
    .C_N(\fetch_prev_state[2] ),
    .X(_0413_));
 sky130_fd_sc_hd__or3b_4 _0855_ (.A(_0413_),
    .B(\fetch_prev_state[1] ),
    .C_N(\fetch_prev_state[0] ),
    .X(_0414_));
 sky130_fd_sc_hd__or4b_1 _0856_ (.A(net34),
    .B(net31),
    .C(\stack[0] ),
    .D_N(net36),
    .X(_0415_));
 sky130_fd_sc_hd__nor2_1 _0857_ (.A(net36),
    .B(net38),
    .Y(_0416_));
 sky130_fd_sc_hd__nor3_2 _0858_ (.A(net34),
    .B(net31),
    .C(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__or3_1 _0859_ (.A(net34),
    .B(net32),
    .C(_0416_),
    .X(_0418_));
 sky130_fd_sc_hd__or4b_1 _0860_ (.A(net39),
    .B(_0414_),
    .C(net20),
    .D_N(_0415_),
    .X(_0419_));
 sky130_fd_sc_hd__o31a_1 _0861_ (.A1(net40),
    .A2(_0414_),
    .A3(_0415_),
    .B1(_0367_),
    .X(_0420_));
 sky130_fd_sc_hd__or3b_1 _0862_ (.A(_0420_),
    .B(_0375_),
    .C_N(_0419_),
    .X(_0421_));
 sky130_fd_sc_hd__and2b_1 _0863_ (.A_N(net38),
    .B(net37),
    .X(_0422_));
 sky130_fd_sc_hd__nand2b_2 _0864_ (.A_N(net38),
    .B(net37),
    .Y(_0423_));
 sky130_fd_sc_hd__or2_1 _0865_ (.A(\stack[0] ),
    .B(net26),
    .X(_0424_));
 sky130_fd_sc_hd__nand2_1 _0866_ (.A(net36),
    .B(net38),
    .Y(_0425_));
 sky130_fd_sc_hd__nand4_1 _0867_ (.A(net58),
    .B(_0417_),
    .C(_0424_),
    .D(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__o21ai_1 _0868_ (.A1(_0419_),
    .A2(_0426_),
    .B1(_0421_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2b_2 _0869_ (.A_N(\fetch_prev_state[0] ),
    .B(\fetch_prev_state[1] ),
    .Y(_0427_));
 sky130_fd_sc_hd__nor2_4 _0870_ (.A(_0413_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__nor2_2 _0871_ (.A(_0367_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__a32o_1 _0872_ (.A1(net28),
    .A2(\timer_period_a[15] ),
    .A3(_0429_),
    .B1(_0428_),
    .B2(net33),
    .X(_0430_));
 sky130_fd_sc_hd__and2_1 _0873_ (.A(net51),
    .B(_0430_),
    .X(_0267_));
 sky130_fd_sc_hd__a32o_1 _0874_ (.A1(net30),
    .A2(\timer_period_a[14] ),
    .A3(_0429_),
    .B1(_0428_),
    .B2(net35),
    .X(_0431_));
 sky130_fd_sc_hd__and2_1 _0875_ (.A(net51),
    .B(_0431_),
    .X(_0266_));
 sky130_fd_sc_hd__a32o_1 _0876_ (.A1(net30),
    .A2(\timer_period_a[13] ),
    .A3(_0429_),
    .B1(_0428_),
    .B2(net36),
    .X(_0432_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(net51),
    .B(_0432_),
    .X(_0265_));
 sky130_fd_sc_hd__a32o_1 _0878_ (.A1(net226),
    .A2(_0374_),
    .A3(_0429_),
    .B1(_0428_),
    .B2(_0372_),
    .X(_0264_));
 sky130_fd_sc_hd__a32o_1 _0879_ (.A1(net30),
    .A2(\timer_period_a[11] ),
    .A3(_0429_),
    .B1(_0428_),
    .B2(net39),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _0880_ (.A(net51),
    .B(_0433_),
    .X(_0263_));
 sky130_fd_sc_hd__a32o_1 _0881_ (.A1(net30),
    .A2(\timer_period_a[10] ),
    .A3(_0429_),
    .B1(_0428_),
    .B2(net43),
    .X(_0434_));
 sky130_fd_sc_hd__and2_1 _0882_ (.A(net51),
    .B(_0434_),
    .X(_0262_));
 sky130_fd_sc_hd__a32o_1 _0883_ (.A1(net30),
    .A2(\timer_period_a[9] ),
    .A3(_0429_),
    .B1(_0428_),
    .B2(\instr[1] ),
    .X(_0435_));
 sky130_fd_sc_hd__and2_1 _0884_ (.A(net51),
    .B(_0435_),
    .X(_0261_));
 sky130_fd_sc_hd__a32o_1 _0885_ (.A1(net28),
    .A2(\timer_period_a[8] ),
    .A3(_0429_),
    .B1(_0428_),
    .B2(net47),
    .X(_0436_));
 sky130_fd_sc_hd__and2_1 _0886_ (.A(net51),
    .B(_0436_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_2 _0887_ (.A(\fetch_prev_state[1] ),
    .B(\fetch_prev_state[0] ),
    .Y(_0437_));
 sky130_fd_sc_hd__nor2_4 _0888_ (.A(_0413_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor2_2 _0889_ (.A(_0367_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a32o_1 _0890_ (.A1(net29),
    .A2(\timer_period_a[7] ),
    .A3(_0439_),
    .B1(_0438_),
    .B2(net32),
    .X(_0440_));
 sky130_fd_sc_hd__and2_1 _0891_ (.A(net55),
    .B(_0440_),
    .X(_0259_));
 sky130_fd_sc_hd__a32o_1 _0892_ (.A1(net29),
    .A2(\timer_period_a[6] ),
    .A3(_0439_),
    .B1(_0438_),
    .B2(net34),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _0893_ (.A(net55),
    .B(_0441_),
    .X(_0258_));
 sky130_fd_sc_hd__a32o_1 _0894_ (.A1(net30),
    .A2(\timer_period_a[5] ),
    .A3(_0439_),
    .B1(_0438_),
    .B2(net36),
    .X(_0442_));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(net56),
    .B(_0442_),
    .X(_0257_));
 sky130_fd_sc_hd__a32o_1 _0896_ (.A1(net225),
    .A2(_0374_),
    .A3(_0439_),
    .B1(_0438_),
    .B2(_0372_),
    .X(_0256_));
 sky130_fd_sc_hd__a32o_1 _0897_ (.A1(net29),
    .A2(\timer_period_a[3] ),
    .A3(_0439_),
    .B1(_0438_),
    .B2(net39),
    .X(_0443_));
 sky130_fd_sc_hd__and2_1 _0898_ (.A(net55),
    .B(_0443_),
    .X(_0255_));
 sky130_fd_sc_hd__a32o_1 _0899_ (.A1(net29),
    .A2(\timer_period_a[2] ),
    .A3(_0439_),
    .B1(_0438_),
    .B2(net43),
    .X(_0444_));
 sky130_fd_sc_hd__and2_1 _0900_ (.A(net55),
    .B(_0444_),
    .X(_0254_));
 sky130_fd_sc_hd__a32o_1 _0901_ (.A1(net29),
    .A2(\timer_period_a[1] ),
    .A3(_0439_),
    .B1(_0438_),
    .B2(\instr[1] ),
    .X(_0445_));
 sky130_fd_sc_hd__and2_1 _0902_ (.A(net55),
    .B(_0445_),
    .X(_0253_));
 sky130_fd_sc_hd__a32o_1 _0903_ (.A1(net30),
    .A2(_0320_),
    .A3(_0439_),
    .B1(_0438_),
    .B2(_0313_),
    .X(_0446_));
 sky130_fd_sc_hd__nand2_1 _0904_ (.A(net51),
    .B(_0446_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2b_1 _0905_ (.A_N(net31),
    .B(net35),
    .Y(_0447_));
 sky130_fd_sc_hd__and4bb_2 _0906_ (.A_N(net31),
    .B_N(_0414_),
    .C(_0416_),
    .D(net34),
    .X(_0448_));
 sky130_fd_sc_hd__nor2_1 _0907_ (.A(_0367_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__a32o_1 _0908_ (.A1(net29),
    .A2(\timer_clock_divisor[3] ),
    .A3(_0449_),
    .B1(_0448_),
    .B2(net39),
    .X(_0450_));
 sky130_fd_sc_hd__and2_1 _0909_ (.A(net55),
    .B(_0450_),
    .X(_0251_));
 sky130_fd_sc_hd__a32o_1 _0910_ (.A1(net29),
    .A2(\timer_clock_divisor[2] ),
    .A3(_0449_),
    .B1(_0448_),
    .B2(net43),
    .X(_0451_));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(net55),
    .B(_0451_),
    .X(_0250_));
 sky130_fd_sc_hd__a32o_1 _0912_ (.A1(net29),
    .A2(\timer_clock_divisor[1] ),
    .A3(_0449_),
    .B1(_0448_),
    .B2(\instr[1] ),
    .X(_0452_));
 sky130_fd_sc_hd__and2_1 _0913_ (.A(net55),
    .B(_0452_),
    .X(_0249_));
 sky130_fd_sc_hd__a32o_1 _0914_ (.A1(net29),
    .A2(\timer_clock_divisor[0] ),
    .A3(_0449_),
    .B1(_0448_),
    .B2(net46),
    .X(_0453_));
 sky130_fd_sc_hd__and2_1 _0915_ (.A(net55),
    .B(_0453_),
    .X(_0248_));
 sky130_fd_sc_hd__o221a_2 _0916_ (.A1(_0334_),
    .A2(_0336_),
    .B1(_0339_),
    .B2(\timer_clock_divisor[3] ),
    .C1(\timer_counter[0] ),
    .X(_0454_));
 sky130_fd_sc_hd__and4_1 _0917_ (.A(\timer_counter[4] ),
    .B(\timer_counter[3] ),
    .C(\timer_counter[2] ),
    .D(\timer_counter[1] ),
    .X(_0455_));
 sky130_fd_sc_hd__and4_1 _0918_ (.A(\timer_counter[8] ),
    .B(\timer_counter[7] ),
    .C(\timer_counter[6] ),
    .D(\timer_counter[5] ),
    .X(_0456_));
 sky130_fd_sc_hd__and3_1 _0919_ (.A(_0454_),
    .B(_0455_),
    .C(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__inv_2 _0920_ (.A(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__and4_1 _0921_ (.A(\timer_counter[9] ),
    .B(_0454_),
    .C(_0455_),
    .D(_0456_),
    .X(_0459_));
 sky130_fd_sc_hd__inv_2 _0922_ (.A(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand2_1 _0923_ (.A(\timer_counter[10] ),
    .B(_0459_),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_1 _0924_ (.A(_0305_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__and4_1 _0925_ (.A(\timer_counter[12] ),
    .B(\timer_counter[11] ),
    .C(\timer_counter[10] ),
    .D(_0459_),
    .X(_0463_));
 sky130_fd_sc_hd__inv_2 _0926_ (.A(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand2_1 _0927_ (.A(\timer_counter[13] ),
    .B(_0463_),
    .Y(_0465_));
 sky130_fd_sc_hd__and3_1 _0928_ (.A(\timer_counter[14] ),
    .B(\timer_counter[13] ),
    .C(_0463_),
    .X(_0466_));
 sky130_fd_sc_hd__or2_1 _0929_ (.A(\timer_counter[15] ),
    .B(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__nor2_1 _0930_ (.A(_0375_),
    .B(_0411_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _0931_ (.A(\timer_counter[15] ),
    .B(_0466_),
    .Y(_0469_));
 sky130_fd_sc_hd__and3_1 _0932_ (.A(_0467_),
    .B(net11),
    .C(_0469_),
    .X(_0247_));
 sky130_fd_sc_hd__a21o_1 _0933_ (.A1(\timer_counter[13] ),
    .A2(_0463_),
    .B1(\timer_counter[14] ),
    .X(_0470_));
 sky130_fd_sc_hd__and3b_1 _0934_ (.A_N(_0466_),
    .B(net11),
    .C(_0470_),
    .X(_0246_));
 sky130_fd_sc_hd__o211a_1 _0935_ (.A1(\timer_counter[13] ),
    .A2(_0463_),
    .B1(_0465_),
    .C1(net11),
    .X(_0245_));
 sky130_fd_sc_hd__o211a_1 _0936_ (.A1(net250),
    .A2(_0462_),
    .B1(_0464_),
    .C1(net11),
    .X(_0244_));
 sky130_fd_sc_hd__nand2_1 _0937_ (.A(_0305_),
    .B(_0461_),
    .Y(_0471_));
 sky130_fd_sc_hd__and3b_1 _0938_ (.A_N(_0462_),
    .B(net11),
    .C(_0471_),
    .X(_0243_));
 sky130_fd_sc_hd__o211a_1 _0939_ (.A1(\timer_counter[10] ),
    .A2(_0459_),
    .B1(_0461_),
    .C1(net11),
    .X(_0242_));
 sky130_fd_sc_hd__o211a_1 _0940_ (.A1(\timer_counter[9] ),
    .A2(_0457_),
    .B1(_0460_),
    .C1(net11),
    .X(_0241_));
 sky130_fd_sc_hd__and2_1 _0941_ (.A(\timer_counter[1] ),
    .B(_0454_),
    .X(_0472_));
 sky130_fd_sc_hd__and3_1 _0942_ (.A(\timer_counter[2] ),
    .B(\timer_counter[1] ),
    .C(_0454_),
    .X(_0473_));
 sky130_fd_sc_hd__and2_1 _0943_ (.A(_0454_),
    .B(_0455_),
    .X(_0474_));
 sky130_fd_sc_hd__and3_1 _0944_ (.A(\timer_counter[5] ),
    .B(_0454_),
    .C(_0455_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _0945_ (.A(\timer_counter[6] ),
    .B(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__and3_1 _0946_ (.A(\timer_counter[7] ),
    .B(\timer_counter[6] ),
    .C(_0475_),
    .X(_0477_));
 sky130_fd_sc_hd__o211a_1 _0947_ (.A1(\timer_counter[8] ),
    .A2(_0477_),
    .B1(net12),
    .C1(_0458_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _0948_ (.A(\timer_counter[7] ),
    .B(_0476_),
    .X(_0478_));
 sky130_fd_sc_hd__and3b_1 _0949_ (.A_N(_0477_),
    .B(_0478_),
    .C(net12),
    .X(_0239_));
 sky130_fd_sc_hd__o21ai_1 _0950_ (.A1(\timer_counter[6] ),
    .A2(_0475_),
    .B1(net11),
    .Y(_0479_));
 sky130_fd_sc_hd__nor2_1 _0951_ (.A(_0476_),
    .B(_0479_),
    .Y(_0238_));
 sky130_fd_sc_hd__or2_1 _0952_ (.A(\timer_counter[5] ),
    .B(_0474_),
    .X(_0480_));
 sky130_fd_sc_hd__and3b_1 _0953_ (.A_N(_0475_),
    .B(_0480_),
    .C(net12),
    .X(_0237_));
 sky130_fd_sc_hd__a21o_1 _0954_ (.A1(\timer_counter[3] ),
    .A2(_0473_),
    .B1(\timer_counter[4] ),
    .X(_0481_));
 sky130_fd_sc_hd__and3b_1 _0955_ (.A_N(_0474_),
    .B(_0481_),
    .C(net11),
    .X(_0236_));
 sky130_fd_sc_hd__o21ai_1 _0956_ (.A1(net220),
    .A2(_0473_),
    .B1(net12),
    .Y(_0482_));
 sky130_fd_sc_hd__a21oi_1 _0957_ (.A1(net220),
    .A2(_0473_),
    .B1(_0482_),
    .Y(_0235_));
 sky130_fd_sc_hd__or2_1 _0958_ (.A(\timer_counter[2] ),
    .B(_0472_),
    .X(_0483_));
 sky130_fd_sc_hd__and3b_1 _0959_ (.A_N(_0473_),
    .B(_0483_),
    .C(net11),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _0960_ (.A(\timer_counter[1] ),
    .B(_0454_),
    .X(_0484_));
 sky130_fd_sc_hd__and3b_1 _0961_ (.A_N(_0472_),
    .B(_0484_),
    .C(net12),
    .X(_0233_));
 sky130_fd_sc_hd__or2_1 _0962_ (.A(\timer_counter[0] ),
    .B(_0340_),
    .X(_0485_));
 sky130_fd_sc_hd__and3b_1 _0963_ (.A_N(_0454_),
    .B(net12),
    .C(_0485_),
    .X(_0232_));
 sky130_fd_sc_hd__nand3_1 _0964_ (.A(\timer_clock_counter[0] ),
    .B(\timer_clock_counter[1] ),
    .C(\timer_clock_counter[2] ),
    .Y(_0486_));
 sky130_fd_sc_hd__and4_1 _0965_ (.A(\timer_clock_counter[0] ),
    .B(\timer_clock_counter[1] ),
    .C(\timer_clock_counter[2] ),
    .D(\timer_clock_counter[3] ),
    .X(_0487_));
 sky130_fd_sc_hd__and3_1 _0966_ (.A(\timer_clock_counter[4] ),
    .B(\timer_clock_counter[5] ),
    .C(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__and4_1 _0967_ (.A(\timer_clock_counter[4] ),
    .B(\timer_clock_counter[5] ),
    .C(\timer_clock_counter[6] ),
    .D(_0487_),
    .X(_0489_));
 sky130_fd_sc_hd__and2_1 _0968_ (.A(\timer_clock_counter[7] ),
    .B(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__and3_1 _0969_ (.A(\timer_clock_counter[7] ),
    .B(\timer_clock_counter[8] ),
    .C(_0489_),
    .X(_0491_));
 sky130_fd_sc_hd__and2_1 _0970_ (.A(\timer_clock_counter[9] ),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__and3_1 _0971_ (.A(\timer_clock_counter[10] ),
    .B(\timer_clock_counter[11] ),
    .C(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _0972_ (.A(\timer_clock_counter[12] ),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and3_1 _0973_ (.A(\timer_clock_counter[13] ),
    .B(\timer_clock_counter[14] ),
    .C(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nor2_1 _0974_ (.A(_0340_),
    .B(_0375_),
    .Y(_0496_));
 sky130_fd_sc_hd__o21a_1 _0975_ (.A1(net211),
    .A2(_0495_),
    .B1(net15),
    .X(_0231_));
 sky130_fd_sc_hd__a31o_1 _0976_ (.A1(\timer_clock_counter[12] ),
    .A2(\timer_clock_counter[13] ),
    .A3(_0493_),
    .B1(\timer_clock_counter[14] ),
    .X(_0497_));
 sky130_fd_sc_hd__and3b_1 _0977_ (.A_N(_0495_),
    .B(net15),
    .C(_0497_),
    .X(_0230_));
 sky130_fd_sc_hd__o21ai_1 _0978_ (.A1(net215),
    .A2(_0494_),
    .B1(net15),
    .Y(_0498_));
 sky130_fd_sc_hd__a21oi_1 _0979_ (.A1(net215),
    .A2(_0494_),
    .B1(_0498_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ai_1 _0980_ (.A1(net236),
    .A2(_0493_),
    .B1(net15),
    .Y(_0499_));
 sky130_fd_sc_hd__nor2_1 _0981_ (.A(_0494_),
    .B(_0499_),
    .Y(_0228_));
 sky130_fd_sc_hd__a31o_1 _0982_ (.A1(\timer_clock_counter[9] ),
    .A2(\timer_clock_counter[10] ),
    .A3(_0491_),
    .B1(\timer_clock_counter[11] ),
    .X(_0500_));
 sky130_fd_sc_hd__and3b_1 _0983_ (.A_N(_0493_),
    .B(net15),
    .C(_0500_),
    .X(_0227_));
 sky130_fd_sc_hd__o21ai_1 _0984_ (.A1(net216),
    .A2(_0492_),
    .B1(net15),
    .Y(_0501_));
 sky130_fd_sc_hd__a21oi_1 _0985_ (.A1(net216),
    .A2(_0492_),
    .B1(_0501_),
    .Y(_0226_));
 sky130_fd_sc_hd__o21ai_1 _0986_ (.A1(net233),
    .A2(_0491_),
    .B1(net15),
    .Y(_0502_));
 sky130_fd_sc_hd__nor2_1 _0987_ (.A(_0492_),
    .B(_0502_),
    .Y(_0225_));
 sky130_fd_sc_hd__o21ai_1 _0988_ (.A1(net218),
    .A2(_0490_),
    .B1(net15),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_1 _0989_ (.A(_0491_),
    .B(_0503_),
    .Y(_0224_));
 sky130_fd_sc_hd__o21ai_1 _0990_ (.A1(net227),
    .A2(_0489_),
    .B1(net15),
    .Y(_0504_));
 sky130_fd_sc_hd__nor2_1 _0991_ (.A(_0490_),
    .B(_0504_),
    .Y(_0223_));
 sky130_fd_sc_hd__o21ai_1 _0992_ (.A1(net219),
    .A2(_0488_),
    .B1(net15),
    .Y(_0505_));
 sky130_fd_sc_hd__nor2_1 _0993_ (.A(_0489_),
    .B(_0505_),
    .Y(_0222_));
 sky130_fd_sc_hd__a21o_1 _0994_ (.A1(\timer_clock_counter[4] ),
    .A2(_0487_),
    .B1(\timer_clock_counter[5] ),
    .X(_0506_));
 sky130_fd_sc_hd__and3b_1 _0995_ (.A_N(_0488_),
    .B(net16),
    .C(_0506_),
    .X(_0221_));
 sky130_fd_sc_hd__o21ai_1 _0996_ (.A1(net221),
    .A2(_0487_),
    .B1(net16),
    .Y(_0507_));
 sky130_fd_sc_hd__a21oi_1 _0997_ (.A1(net221),
    .A2(_0487_),
    .B1(_0507_),
    .Y(_0220_));
 sky130_fd_sc_hd__a31o_1 _0998_ (.A1(\timer_clock_counter[0] ),
    .A2(\timer_clock_counter[1] ),
    .A3(\timer_clock_counter[2] ),
    .B1(\timer_clock_counter[3] ),
    .X(_0508_));
 sky130_fd_sc_hd__and3b_1 _0999_ (.A_N(_0487_),
    .B(net16),
    .C(_0508_),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_1 _1000_ (.A1(\timer_clock_counter[0] ),
    .A2(\timer_clock_counter[1] ),
    .B1(\timer_clock_counter[2] ),
    .X(_0509_));
 sky130_fd_sc_hd__and3_1 _1001_ (.A(_0486_),
    .B(net16),
    .C(_0509_),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1002_ (.A1(\timer_clock_counter[0] ),
    .A2(\timer_clock_counter[1] ),
    .B1(net16),
    .Y(_0510_));
 sky130_fd_sc_hd__a21oi_1 _1003_ (.A1(net239),
    .A2(\timer_clock_counter[1] ),
    .B1(_0510_),
    .Y(_0217_));
 sky130_fd_sc_hd__and2b_1 _1004_ (.A_N(\timer_clock_counter[0] ),
    .B(net16),
    .X(_0216_));
 sky130_fd_sc_hd__nor2_1 _1005_ (.A(net34),
    .B(_0414_),
    .Y(_0511_));
 sky130_fd_sc_hd__or2_1 _1006_ (.A(net34),
    .B(_0414_),
    .X(_0512_));
 sky130_fd_sc_hd__or3b_1 _1007_ (.A(_0512_),
    .B(\stack[14] ),
    .C_N(_0416_),
    .X(_0513_));
 sky130_fd_sc_hd__a21o_1 _1008_ (.A1(_0416_),
    .A2(_0511_),
    .B1(\stack[15] ),
    .X(_0514_));
 sky130_fd_sc_hd__and3_1 _1009_ (.A(net58),
    .B(_0513_),
    .C(_0514_),
    .X(_0215_));
 sky130_fd_sc_hd__and2b_1 _1010_ (.A_N(\fetch_state[2] ),
    .B(net48),
    .X(_0515_));
 sky130_fd_sc_hd__nor2_1 _1011_ (.A(\fetch_state[1] ),
    .B(\fetch_state[0] ),
    .Y(_0516_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(\fetch_state[1] ),
    .B(\fetch_state[0] ),
    .X(_0517_));
 sky130_fd_sc_hd__and2b_1 _1013_ (.A_N(net48),
    .B(\fetch_state[2] ),
    .X(_0518_));
 sky130_fd_sc_hd__a21oi_2 _1014_ (.A1(_0517_),
    .A2(_0518_),
    .B1(_0515_),
    .Y(_0519_));
 sky130_fd_sc_hd__a21o_2 _1015_ (.A1(_0517_),
    .A2(_0518_),
    .B1(_0515_),
    .X(_0520_));
 sky130_fd_sc_hd__or2_1 _1016_ (.A(net35),
    .B(_0519_),
    .X(_0521_));
 sky130_fd_sc_hd__o211a_1 _1017_ (.A1(net31),
    .A2(net18),
    .B1(_0521_),
    .C1(net53),
    .X(_0214_));
 sky130_fd_sc_hd__or2_1 _1018_ (.A(net36),
    .B(_0519_),
    .X(_0522_));
 sky130_fd_sc_hd__o211a_1 _1019_ (.A1(net35),
    .A2(net18),
    .B1(_0522_),
    .C1(net58),
    .X(_0213_));
 sky130_fd_sc_hd__or2_1 _1020_ (.A(net38),
    .B(_0519_),
    .X(_0523_));
 sky130_fd_sc_hd__o211a_1 _1021_ (.A1(net36),
    .A2(net18),
    .B1(_0523_),
    .C1(net53),
    .X(_0212_));
 sky130_fd_sc_hd__nand2_1 _1022_ (.A(net56),
    .B(net18),
    .Y(_0524_));
 sky130_fd_sc_hd__a2bb2oi_1 _1023_ (.A1_N(net39),
    .A2_N(_0519_),
    .B1(_0524_),
    .B2(_0373_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _1024_ (.A(_0311_),
    .B(_0520_),
    .Y(_0525_));
 sky130_fd_sc_hd__o211a_1 _1025_ (.A1(net39),
    .A2(_0520_),
    .B1(_0525_),
    .C1(net58),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _1026_ (.A(_0312_),
    .B(net18),
    .Y(_0526_));
 sky130_fd_sc_hd__o211a_1 _1027_ (.A1(net44),
    .A2(net18),
    .B1(_0526_),
    .C1(net53),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _1028_ (.A(_0313_),
    .B(net18),
    .Y(_0527_));
 sky130_fd_sc_hd__o211a_1 _1029_ (.A1(net45),
    .A2(net18),
    .B1(_0527_),
    .C1(net56),
    .X(_0208_));
 sky130_fd_sc_hd__or2_1 _1030_ (.A(\uio_in_reg[3] ),
    .B(_0519_),
    .X(_0528_));
 sky130_fd_sc_hd__o211a_1 _1031_ (.A1(net46),
    .A2(net18),
    .B1(_0528_),
    .C1(net58),
    .X(_0207_));
 sky130_fd_sc_hd__nor2_1 _1032_ (.A(_0331_),
    .B(_0427_),
    .Y(_0529_));
 sky130_fd_sc_hd__or2_2 _1033_ (.A(_0331_),
    .B(_0427_),
    .X(_0530_));
 sky130_fd_sc_hd__or2_1 _1034_ (.A(\cycle_end_addr[7] ),
    .B(_0529_),
    .X(_0531_));
 sky130_fd_sc_hd__o211a_1 _1035_ (.A1(net32),
    .A2(_0530_),
    .B1(_0531_),
    .C1(net57),
    .X(_0206_));
 sky130_fd_sc_hd__or2_1 _1036_ (.A(net261),
    .B(_0529_),
    .X(_0532_));
 sky130_fd_sc_hd__o211a_1 _1037_ (.A1(net34),
    .A2(_0530_),
    .B1(_0532_),
    .C1(net56),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _1038_ (.A(\cycle_end_addr[5] ),
    .B(_0529_),
    .X(_0533_));
 sky130_fd_sc_hd__o211a_1 _1039_ (.A1(net36),
    .A2(_0530_),
    .B1(_0533_),
    .C1(net56),
    .X(_0204_));
 sky130_fd_sc_hd__or2_1 _1040_ (.A(\cycle_end_addr[4] ),
    .B(_0529_),
    .X(_0534_));
 sky130_fd_sc_hd__o211a_1 _1041_ (.A1(net38),
    .A2(_0530_),
    .B1(_0534_),
    .C1(net57),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _1042_ (.A(\cycle_end_addr[3] ),
    .B(_0529_),
    .X(_0535_));
 sky130_fd_sc_hd__o211a_1 _1043_ (.A1(net39),
    .A2(_0530_),
    .B1(_0535_),
    .C1(net56),
    .X(_0202_));
 sky130_fd_sc_hd__or2_1 _1044_ (.A(\cycle_end_addr[2] ),
    .B(_0529_),
    .X(_0536_));
 sky130_fd_sc_hd__o211a_1 _1045_ (.A1(net43),
    .A2(_0530_),
    .B1(_0536_),
    .C1(net57),
    .X(_0201_));
 sky130_fd_sc_hd__or2_1 _1046_ (.A(net253),
    .B(_0529_),
    .X(_0537_));
 sky130_fd_sc_hd__o211a_1 _1047_ (.A1(\instr[1] ),
    .A2(_0530_),
    .B1(_0537_),
    .C1(net57),
    .X(_0200_));
 sky130_fd_sc_hd__or2_1 _1048_ (.A(net238),
    .B(_0529_),
    .X(_0538_));
 sky130_fd_sc_hd__o211a_1 _1049_ (.A1(net46),
    .A2(_0530_),
    .B1(_0538_),
    .C1(net56),
    .X(_0199_));
 sky130_fd_sc_hd__nor2_1 _1050_ (.A(_0331_),
    .B(_0437_),
    .Y(_0539_));
 sky130_fd_sc_hd__or2_2 _1051_ (.A(_0331_),
    .B(_0437_),
    .X(_0540_));
 sky130_fd_sc_hd__or2_1 _1052_ (.A(net257),
    .B(_0539_),
    .X(_0541_));
 sky130_fd_sc_hd__o211a_1 _1053_ (.A1(net33),
    .A2(_0540_),
    .B1(_0541_),
    .C1(net52),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _1054_ (.A(net260),
    .B(_0539_),
    .X(_0542_));
 sky130_fd_sc_hd__o211a_1 _1055_ (.A1(\instr[6] ),
    .A2(_0540_),
    .B1(_0542_),
    .C1(net52),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _1056_ (.A(net262),
    .B(_0539_),
    .X(_0543_));
 sky130_fd_sc_hd__o211a_1 _1057_ (.A1(net37),
    .A2(_0540_),
    .B1(_0543_),
    .C1(net52),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _1058_ (.A(net256),
    .B(_0539_),
    .X(_0544_));
 sky130_fd_sc_hd__o211a_1 _1059_ (.A1(net38),
    .A2(_0540_),
    .B1(_0544_),
    .C1(net52),
    .X(_0195_));
 sky130_fd_sc_hd__or2_1 _1060_ (.A(\cycle_start_addr[3] ),
    .B(_0539_),
    .X(_0545_));
 sky130_fd_sc_hd__o211a_1 _1061_ (.A1(net41),
    .A2(_0540_),
    .B1(_0545_),
    .C1(net52),
    .X(_0194_));
 sky130_fd_sc_hd__or2_1 _1062_ (.A(net255),
    .B(_0539_),
    .X(_0546_));
 sky130_fd_sc_hd__o211a_1 _1063_ (.A1(net44),
    .A2(_0540_),
    .B1(_0546_),
    .C1(net52),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _1064_ (.A(net263),
    .B(_0539_),
    .X(_0547_));
 sky130_fd_sc_hd__o211a_1 _1065_ (.A1(net45),
    .A2(_0540_),
    .B1(_0547_),
    .C1(net52),
    .X(_0192_));
 sky130_fd_sc_hd__or2_1 _1066_ (.A(net254),
    .B(_0539_),
    .X(_0548_));
 sky130_fd_sc_hd__o211a_1 _1067_ (.A1(net47),
    .A2(_0540_),
    .B1(_0548_),
    .C1(net52),
    .X(_0191_));
 sky130_fd_sc_hd__or2_1 _1068_ (.A(_0302_),
    .B(net224),
    .X(_0190_));
 sky130_fd_sc_hd__nor2_2 _1069_ (.A(_0312_),
    .B(_0313_),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_1 _1070_ (.A(net45),
    .B(net46),
    .Y(_0550_));
 sky130_fd_sc_hd__or4bb_1 _1071_ (.A(net34),
    .B(net31),
    .C_N(net37),
    .D_N(net38),
    .X(_0551_));
 sky130_fd_sc_hd__nor2_2 _1072_ (.A(_0312_),
    .B(net46),
    .Y(_0552_));
 sky130_fd_sc_hd__and2b_2 _1073_ (.A_N(net45),
    .B(net46),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_1 _1074_ (.A1(uo_out[7]),
    .A2(_0549_),
    .B1(_0553_),
    .B2(uo_out[5]),
    .X(_0554_));
 sky130_fd_sc_hd__nor2_2 _1075_ (.A(net45),
    .B(net46),
    .Y(_0555_));
 sky130_fd_sc_hd__a221o_1 _1076_ (.A1(uo_out[6]),
    .A2(_0552_),
    .B1(_0555_),
    .B2(uo_out[4]),
    .C1(_0311_),
    .X(_0556_));
 sky130_fd_sc_hd__a22o_1 _1077_ (.A1(uo_out[1]),
    .A2(_0553_),
    .B1(_0555_),
    .B2(uo_out[0]),
    .X(_0557_));
 sky130_fd_sc_hd__a221o_1 _1078_ (.A1(uo_out[3]),
    .A2(_0549_),
    .B1(_0552_),
    .B2(uo_out[2]),
    .C1(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__o22ai_1 _1079_ (.A1(_0554_),
    .A2(_0556_),
    .B1(_0558_),
    .B2(net42),
    .Y(_0559_));
 sky130_fd_sc_hd__a2bb2o_2 _1080_ (.A1_N(_0415_),
    .A2_N(_0559_),
    .B1(_0551_),
    .B2(\stack[0] ),
    .X(_0560_));
 sky130_fd_sc_hd__and2b_1 _1081_ (.A_N(net34),
    .B(net31),
    .X(_0561_));
 sky130_fd_sc_hd__nand2b_1 _1082_ (.A_N(net35),
    .B(net31),
    .Y(_0562_));
 sky130_fd_sc_hd__a31o_1 _1083_ (.A1(net42),
    .A2(net45),
    .A3(net46),
    .B1(uo_out[7]),
    .X(_0563_));
 sky130_fd_sc_hd__o311a_1 _1084_ (.A1(_0311_),
    .A2(_0550_),
    .A3(_0560_),
    .B1(net22),
    .C1(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__o21a_1 _1085_ (.A1(net36),
    .A2(net38),
    .B1(net39),
    .X(_0565_));
 sky130_fd_sc_hd__o21a_1 _1086_ (.A1(net31),
    .A2(_0565_),
    .B1(_0511_),
    .X(_0566_));
 sky130_fd_sc_hd__o21ai_2 _1087_ (.A1(net31),
    .A2(_0565_),
    .B1(_0511_),
    .Y(_0567_));
 sky130_fd_sc_hd__a211o_1 _1088_ (.A1(net40),
    .A2(net24),
    .B1(_0564_),
    .C1(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__o211a_1 _1089_ (.A1(uo_out[7]),
    .A2(_0566_),
    .B1(_0568_),
    .C1(net53),
    .X(_0189_));
 sky130_fd_sc_hd__nand2_1 _1090_ (.A(net42),
    .B(_0552_),
    .Y(_0569_));
 sky130_fd_sc_hd__a21o_1 _1091_ (.A1(net42),
    .A2(_0552_),
    .B1(uo_out[6]),
    .X(_0570_));
 sky130_fd_sc_hd__o211a_1 _1092_ (.A1(_0560_),
    .A2(_0569_),
    .B1(_0570_),
    .C1(net22),
    .X(_0571_));
 sky130_fd_sc_hd__a21o_1 _1093_ (.A1(net42),
    .A2(net24),
    .B1(_0567_),
    .X(_0572_));
 sky130_fd_sc_hd__o221a_1 _1094_ (.A1(uo_out[6]),
    .A2(_0566_),
    .B1(_0571_),
    .B2(_0572_),
    .C1(net53),
    .X(_0188_));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(net42),
    .B(_0553_),
    .Y(_0573_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(_0560_),
    .A1(uo_out[5]),
    .S(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__or2_1 _1097_ (.A(uo_out[5]),
    .B(_0566_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _1098_ (.A0(net45),
    .A1(_0574_),
    .S(net22),
    .X(_0576_));
 sky130_fd_sc_hd__o211a_1 _1099_ (.A1(_0567_),
    .A2(_0576_),
    .B1(_0575_),
    .C1(net58),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_1 _1100_ (.A(net42),
    .B(_0555_),
    .Y(_0577_));
 sky130_fd_sc_hd__a21o_1 _1101_ (.A1(net42),
    .A2(_0555_),
    .B1(uo_out[4]),
    .X(_0578_));
 sky130_fd_sc_hd__o211a_1 _1102_ (.A1(_0560_),
    .A2(_0577_),
    .B1(_0578_),
    .C1(net22),
    .X(_0579_));
 sky130_fd_sc_hd__a211o_1 _1103_ (.A1(net46),
    .A2(net24),
    .B1(_0567_),
    .C1(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__o211a_1 _1104_ (.A1(uo_out[4]),
    .A2(_0566_),
    .B1(_0580_),
    .C1(net53),
    .X(_0186_));
 sky130_fd_sc_hd__and4_1 _1105_ (.A(net57),
    .B(\cur_addr[1] ),
    .C(\cur_addr[0] ),
    .D(_0520_),
    .X(_0581_));
 sky130_fd_sc_hd__and3_1 _1106_ (.A(\cur_addr[3] ),
    .B(\cur_addr[2] ),
    .C(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__and2_1 _1107_ (.A(\cur_addr[4] ),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__and3_1 _1108_ (.A(\cur_addr[6] ),
    .B(\cur_addr[5] ),
    .C(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__xnor2_1 _1109_ (.A(_0314_),
    .B(_0584_),
    .Y(_0185_));
 sky130_fd_sc_hd__a21oi_1 _1110_ (.A1(\cur_addr[5] ),
    .A2(_0583_),
    .B1(net234),
    .Y(_0585_));
 sky130_fd_sc_hd__nor2_1 _1111_ (.A(_0584_),
    .B(net235),
    .Y(_0184_));
 sky130_fd_sc_hd__xnor2_1 _1112_ (.A(_0315_),
    .B(_0583_),
    .Y(_0183_));
 sky130_fd_sc_hd__nor2_1 _1113_ (.A(net232),
    .B(_0582_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_1 _1114_ (.A(_0583_),
    .B(_0586_),
    .Y(_0182_));
 sky130_fd_sc_hd__a21oi_1 _1115_ (.A1(\cur_addr[2] ),
    .A2(_0581_),
    .B1(net229),
    .Y(_0587_));
 sky130_fd_sc_hd__nor2_1 _1116_ (.A(_0582_),
    .B(net230),
    .Y(_0181_));
 sky130_fd_sc_hd__xnor2_1 _1117_ (.A(_0318_),
    .B(_0581_),
    .Y(_0180_));
 sky130_fd_sc_hd__a31o_1 _1118_ (.A1(net57),
    .A2(\cur_addr[0] ),
    .A3(_0520_),
    .B1(\cur_addr[1] ),
    .X(_0588_));
 sky130_fd_sc_hd__and2b_1 _1119_ (.A_N(_0581_),
    .B(_0588_),
    .X(_0179_));
 sky130_fd_sc_hd__xnor2_1 _1120_ (.A(net246),
    .B(_0524_),
    .Y(_0178_));
 sky130_fd_sc_hd__and2b_1 _1121_ (.A_N(\fetch_state[0] ),
    .B(\fetch_state[1] ),
    .X(_0589_));
 sky130_fd_sc_hd__or3_2 _1122_ (.A(net48),
    .B(\fetch_state[2] ),
    .C(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__inv_2 _1123_ (.A(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__o31ai_4 _1124_ (.A1(\fetch_count[2] ),
    .A2(\fetch_count[1] ),
    .A3(\fetch_count[0] ),
    .B1(_0590_),
    .Y(_0592_));
 sky130_fd_sc_hd__inv_2 _1125_ (.A(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _1126_ (.A(net52),
    .B(_0592_),
    .Y(_0594_));
 sky130_fd_sc_hd__mux2_1 _1127_ (.A0(net48),
    .A1(net217),
    .S(_0594_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _1128_ (.A0(\fetch_state[2] ),
    .A1(net213),
    .S(_0594_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _1129_ (.A0(net248),
    .A1(\fetch_prev_state[1] ),
    .S(_0594_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _1130_ (.A0(\fetch_state[0] ),
    .A1(net258),
    .S(_0594_),
    .X(_0174_));
 sky130_fd_sc_hd__and3_1 _1131_ (.A(net48),
    .B(\fetch_state[2] ),
    .C(_0516_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _1132_ (.A(\fetch_state[1] ),
    .B(\fetch_state[0] ),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_1 _1133_ (.A(\fetch_state[2] ),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__and2b_1 _1134_ (.A_N(\fetch_state[1] ),
    .B(\fetch_state[0] ),
    .X(_0598_));
 sky130_fd_sc_hd__and4bb_1 _1135_ (.A_N(net48),
    .B_N(\fetch_state[2] ),
    .C(\fetch_state[1] ),
    .D(\fetch_state[0] ),
    .X(_0599_));
 sky130_fd_sc_hd__a31o_1 _1136_ (.A1(net48),
    .A2(\fetch_state[2] ),
    .A3(_0598_),
    .B1(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__or2_1 _1137_ (.A(_0595_),
    .B(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__nor2_1 _1138_ (.A(net18),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__or2_1 _1139_ (.A(\fetch_count[0] ),
    .B(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__or2_1 _1140_ (.A(\fetch_count[1] ),
    .B(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__o21ai_1 _1141_ (.A1(\fetch_count[2] ),
    .A2(_0604_),
    .B1(net53),
    .Y(_0605_));
 sky130_fd_sc_hd__a21o_1 _1142_ (.A1(\fetch_count[2] ),
    .A2(_0604_),
    .B1(_0605_),
    .X(_0173_));
 sky130_fd_sc_hd__a21oi_1 _1143_ (.A1(\fetch_count[1] ),
    .A2(_0603_),
    .B1(_0302_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _1144_ (.A(_0604_),
    .B(_0606_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _1145_ (.A(net53),
    .B(_0603_),
    .Y(_0607_));
 sky130_fd_sc_hd__a21o_1 _1146_ (.A1(\fetch_count[0] ),
    .A2(_0602_),
    .B1(_0607_),
    .X(_0171_));
 sky130_fd_sc_hd__or4_1 _1147_ (.A(\cycle_start_addr[3] ),
    .B(\cycle_start_addr[2] ),
    .C(\cycle_start_addr[1] ),
    .D(\cycle_start_addr[0] ),
    .X(_0608_));
 sky130_fd_sc_hd__or4_1 _1148_ (.A(\cycle_start_addr[7] ),
    .B(\cycle_start_addr[6] ),
    .C(\cycle_start_addr[5] ),
    .D(\cycle_start_addr[4] ),
    .X(_0609_));
 sky130_fd_sc_hd__nor2_1 _1149_ (.A(_0608_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__a22o_1 _1150_ (.A1(net48),
    .A2(_0597_),
    .B1(_0610_),
    .B2(_0595_),
    .X(_0611_));
 sky130_fd_sc_hd__a2111o_1 _1151_ (.A1(_0515_),
    .A2(_0516_),
    .B1(_0593_),
    .C1(_0600_),
    .D1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__and2_1 _1152_ (.A(_0518_),
    .B(_0598_),
    .X(_0613_));
 sky130_fd_sc_hd__nand2b_1 _1153_ (.A_N(\cycle_end_addr[6] ),
    .B(\cur_addr[6] ),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2b_1 _1154_ (.A_N(\cycle_end_addr[1] ),
    .B(\cur_addr[1] ),
    .Y(_0615_));
 sky130_fd_sc_hd__and2b_1 _1155_ (.A_N(\cur_addr[1] ),
    .B(\cycle_end_addr[1] ),
    .X(_0616_));
 sky130_fd_sc_hd__nand2b_1 _1156_ (.A_N(\cycle_end_addr[0] ),
    .B(\cur_addr[0] ),
    .Y(_0617_));
 sky130_fd_sc_hd__a221o_1 _1157_ (.A1(\cycle_end_addr[2] ),
    .A2(_0318_),
    .B1(_0615_),
    .B2(_0617_),
    .C1(_0616_),
    .X(_0618_));
 sky130_fd_sc_hd__o22a_1 _1158_ (.A1(\cycle_end_addr[3] ),
    .A2(_0317_),
    .B1(_0318_),
    .B2(\cycle_end_addr[2] ),
    .X(_0619_));
 sky130_fd_sc_hd__a22o_1 _1159_ (.A1(\cycle_end_addr[4] ),
    .A2(_0316_),
    .B1(_0317_),
    .B2(\cycle_end_addr[3] ),
    .X(_0620_));
 sky130_fd_sc_hd__a21o_1 _1160_ (.A1(_0618_),
    .A2(_0619_),
    .B1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__o22a_1 _1161_ (.A1(\cycle_end_addr[5] ),
    .A2(_0315_),
    .B1(_0316_),
    .B2(\cycle_end_addr[4] ),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _1162_ (.A1(\cycle_end_addr[5] ),
    .A2(_0315_),
    .B1(_0621_),
    .B2(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__and2b_1 _1163_ (.A_N(\cur_addr[6] ),
    .B(\cycle_end_addr[6] ),
    .X(_0624_));
 sky130_fd_sc_hd__a221o_1 _1164_ (.A1(\cycle_end_addr[7] ),
    .A2(_0314_),
    .B1(_0614_),
    .B2(_0623_),
    .C1(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__or4_1 _1165_ (.A(\cur_addr[3] ),
    .B(\cur_addr[2] ),
    .C(\cur_addr[1] ),
    .D(\cur_addr[0] ),
    .X(_0626_));
 sky130_fd_sc_hd__or4_1 _1166_ (.A(\cur_addr[7] ),
    .B(\cur_addr[6] ),
    .C(\cur_addr[5] ),
    .D(\cur_addr[4] ),
    .X(_0627_));
 sky130_fd_sc_hd__o22a_1 _1167_ (.A1(\cycle_end_addr[7] ),
    .A2(_0314_),
    .B1(_0626_),
    .B2(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__and3_1 _1168_ (.A(_0613_),
    .B(_0625_),
    .C(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__nor4_2 _1169_ (.A(net41),
    .B(net42),
    .C(_0425_),
    .D(_0447_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_1 _1170_ (.A(_0553_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__a31o_1 _1171_ (.A1(_0553_),
    .A2(_0629_),
    .A3(_0630_),
    .B1(_0612_),
    .X(_0632_));
 sky130_fd_sc_hd__o211a_1 _1172_ (.A1(net48),
    .A2(_0592_),
    .B1(_0632_),
    .C1(net54),
    .X(_0170_));
 sky130_fd_sc_hd__and3_1 _1173_ (.A(_0515_),
    .B(_0517_),
    .C(_0596_),
    .X(_0633_));
 sky130_fd_sc_hd__a211o_1 _1174_ (.A1(\fetch_state[1] ),
    .A2(_0518_),
    .B1(_0593_),
    .C1(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__and2b_1 _1175_ (.A_N(_0610_),
    .B(_0595_),
    .X(_0635_));
 sky130_fd_sc_hd__a2111o_1 _1176_ (.A1(_0629_),
    .A2(_0631_),
    .B1(_0634_),
    .C1(_0635_),
    .D1(_0600_),
    .X(_0636_));
 sky130_fd_sc_hd__o211a_1 _1177_ (.A1(\fetch_state[2] ),
    .A2(_0592_),
    .B1(_0636_),
    .C1(net53),
    .X(_0169_));
 sky130_fd_sc_hd__nor3b_1 _1178_ (.A(net48),
    .B(\fetch_state[2] ),
    .C_N(_0598_),
    .Y(_0637_));
 sky130_fd_sc_hd__a2111o_1 _1179_ (.A1(_0518_),
    .A2(_0589_),
    .B1(_0593_),
    .C1(_0611_),
    .D1(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__a31o_1 _1180_ (.A1(_0555_),
    .A2(_0629_),
    .A3(_0630_),
    .B1(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__o211a_1 _1181_ (.A1(net248),
    .A2(_0592_),
    .B1(_0639_),
    .C1(net54),
    .X(_0168_));
 sky130_fd_sc_hd__and3_1 _1182_ (.A(_0625_),
    .B(_0628_),
    .C(_0630_),
    .X(_0640_));
 sky130_fd_sc_hd__a21boi_1 _1183_ (.A1(_0312_),
    .A2(_0640_),
    .B1_N(_0613_),
    .Y(_0641_));
 sky130_fd_sc_hd__a211o_1 _1184_ (.A1(\fetch_state[3] ),
    .A2(_0516_),
    .B1(_0591_),
    .C1(_0634_),
    .X(_0642_));
 sky130_fd_sc_hd__o221a_1 _1185_ (.A1(\fetch_state[0] ),
    .A2(_0592_),
    .B1(_0641_),
    .B2(_0642_),
    .C1(net54),
    .X(_0167_));
 sky130_fd_sc_hd__a211o_1 _1186_ (.A1(net222),
    .A2(_0602_),
    .B1(_0637_),
    .C1(_0302_),
    .X(_0166_));
 sky130_fd_sc_hd__or4_1 _1187_ (.A(\timer_period_b[1] ),
    .B(\timer_period_b[2] ),
    .C(\timer_period_b[3] ),
    .D(\timer_period_b[4] ),
    .X(_0643_));
 sky130_fd_sc_hd__or3_1 _1188_ (.A(\timer_period_b[13] ),
    .B(\timer_period_b[14] ),
    .C(\timer_period_b[15] ),
    .X(_0644_));
 sky130_fd_sc_hd__or4_1 _1189_ (.A(\timer_period_b[9] ),
    .B(\timer_period_b[10] ),
    .C(\timer_period_b[11] ),
    .D(\timer_period_b[12] ),
    .X(_0645_));
 sky130_fd_sc_hd__or4_1 _1190_ (.A(\timer_period_b[5] ),
    .B(\timer_period_b[6] ),
    .C(\timer_period_b[7] ),
    .D(\timer_period_b[8] ),
    .X(_0646_));
 sky130_fd_sc_hd__nor3_1 _1191_ (.A(_0644_),
    .B(_0645_),
    .C(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _1192_ (.A(net17),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__o41a_1 _1193_ (.A1(timer_mode),
    .A2(\timer_period_b[0] ),
    .A3(_0643_),
    .A4(_0648_),
    .B1(_0411_),
    .X(_0649_));
 sky130_fd_sc_hd__a21oi_1 _1194_ (.A1(timer_mode),
    .A2(net17),
    .B1(timer_out),
    .Y(_0650_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(timer_out),
    .A1(_0650_),
    .S(_0649_),
    .X(_0651_));
 sky130_fd_sc_hd__and3_1 _1196_ (.A(net54),
    .B(net28),
    .C(_0651_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _1197_ (.A0(\cycle_start_addr[2] ),
    .A1(\cycle_start_addr[3] ),
    .S(\fetch_count[0] ),
    .X(_0652_));
 sky130_fd_sc_hd__mux4_1 _1198_ (.A0(\cycle_start_addr[4] ),
    .A1(\cycle_start_addr[5] ),
    .A2(\cycle_start_addr[6] ),
    .A3(\cycle_start_addr[7] ),
    .S0(\fetch_count[0] ),
    .S1(\fetch_count[1] ),
    .X(_0653_));
 sky130_fd_sc_hd__nand3_1 _1199_ (.A(\fetch_count[2] ),
    .B(_0595_),
    .C(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(\cycle_start_addr[0] ),
    .A1(\cycle_start_addr[1] ),
    .S(\fetch_count[0] ),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _1201_ (.A(_0595_),
    .B(_0652_),
    .Y(_0656_));
 sky130_fd_sc_hd__nor2_1 _1202_ (.A(\fetch_count[1] ),
    .B(_0655_),
    .Y(_0657_));
 sky130_fd_sc_hd__a221o_1 _1203_ (.A1(\fetch_count[1] ),
    .A2(_0656_),
    .B1(_0657_),
    .B2(_0595_),
    .C1(\fetch_count[2] ),
    .X(_0658_));
 sky130_fd_sc_hd__a31o_1 _1204_ (.A1(_0601_),
    .A2(_0654_),
    .A3(_0658_),
    .B1(_0302_),
    .X(_0659_));
 sky130_fd_sc_hd__o21ba_1 _1205_ (.A1(net212),
    .A2(_0601_),
    .B1_N(_0659_),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _1206_ (.A1(\ui_in_reg[3] ),
    .A2(_0549_),
    .B1(_0555_),
    .B2(\ui_in_reg[0] ),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_1 _1207_ (.A(net40),
    .B(_0559_),
    .Y(_0661_));
 sky130_fd_sc_hd__a211o_1 _1208_ (.A1(\ui_in_reg[4] ),
    .A2(_0555_),
    .B1(net40),
    .C1(_0311_),
    .X(_0662_));
 sky130_fd_sc_hd__a22o_1 _1209_ (.A1(\ui_in_reg[6] ),
    .A2(_0552_),
    .B1(_0553_),
    .B2(\ui_in_reg[5] ),
    .X(_0663_));
 sky130_fd_sc_hd__a211o_1 _1210_ (.A1(\ui_in_reg[7] ),
    .A2(_0549_),
    .B1(_0662_),
    .C1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__a211o_1 _1211_ (.A1(\ui_in_reg[2] ),
    .A2(_0552_),
    .B1(net40),
    .C1(net42),
    .X(_0665_));
 sky130_fd_sc_hd__a211o_1 _1212_ (.A1(\ui_in_reg[1] ),
    .A2(_0553_),
    .B1(_0660_),
    .C1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__a31o_1 _1213_ (.A1(_0661_),
    .A2(_0664_),
    .A3(_0666_),
    .B1(_0417_),
    .X(_0667_));
 sky130_fd_sc_hd__o211a_1 _1214_ (.A1(\stack[1] ),
    .A2(net20),
    .B1(net22),
    .C1(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__mux4_1 _1215_ (.A0(net39),
    .A1(net43),
    .A2(net45),
    .A3(net46),
    .S0(\stack[0] ),
    .S1(\stack[1] ),
    .X(_0669_));
 sky130_fd_sc_hd__a21o_1 _1216_ (.A1(net24),
    .A2(_0669_),
    .B1(_0512_),
    .X(_0670_));
 sky130_fd_sc_hd__o221a_1 _1217_ (.A1(\stack[0] ),
    .A2(_0511_),
    .B1(_0668_),
    .B2(_0670_),
    .C1(net58),
    .X(_0163_));
 sky130_fd_sc_hd__a21oi_2 _1218_ (.A1(net32),
    .A2(\instr[4] ),
    .B1(_0512_),
    .Y(_0671_));
 sky130_fd_sc_hd__a21o_1 _1219_ (.A1(net32),
    .A2(\instr[4] ),
    .B1(_0512_),
    .X(_0672_));
 sky130_fd_sc_hd__or2_1 _1220_ (.A(\stack[13] ),
    .B(net26),
    .X(_0673_));
 sky130_fd_sc_hd__o211a_1 _1221_ (.A1(\stack[15] ),
    .A2(net25),
    .B1(net23),
    .C1(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _1222_ (.A0(\stack[15] ),
    .A1(\stack[13] ),
    .S(net20),
    .X(_0675_));
 sky130_fd_sc_hd__a211o_1 _1223_ (.A1(net21),
    .A2(_0675_),
    .B1(_0674_),
    .C1(net13),
    .X(_0676_));
 sky130_fd_sc_hd__o211a_1 _1224_ (.A1(net237),
    .A2(net14),
    .B1(_0676_),
    .C1(net59),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _1225_ (.A(\stack[12] ),
    .B(net26),
    .X(_0677_));
 sky130_fd_sc_hd__o211a_1 _1226_ (.A1(\stack[14] ),
    .A2(net25),
    .B1(net23),
    .C1(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _1227_ (.A0(\stack[14] ),
    .A1(\stack[12] ),
    .S(net19),
    .X(_0679_));
 sky130_fd_sc_hd__a211o_1 _1228_ (.A1(net21),
    .A2(_0679_),
    .B1(_0678_),
    .C1(net13),
    .X(_0680_));
 sky130_fd_sc_hd__o211a_1 _1229_ (.A1(net249),
    .A2(net14),
    .B1(_0680_),
    .C1(net59),
    .X(_0161_));
 sky130_fd_sc_hd__or2_1 _1230_ (.A(\stack[11] ),
    .B(net26),
    .X(_0681_));
 sky130_fd_sc_hd__o211a_1 _1231_ (.A1(\stack[13] ),
    .A2(_0423_),
    .B1(net23),
    .C1(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _1232_ (.A0(\stack[13] ),
    .A1(\stack[11] ),
    .S(net19),
    .X(_0683_));
 sky130_fd_sc_hd__a211o_1 _1233_ (.A1(net21),
    .A2(_0683_),
    .B1(_0682_),
    .C1(net13),
    .X(_0684_));
 sky130_fd_sc_hd__o211a_1 _1234_ (.A1(net259),
    .A2(net14),
    .B1(_0684_),
    .C1(net59),
    .X(_0160_));
 sky130_fd_sc_hd__or2_1 _1235_ (.A(\stack[10] ),
    .B(_0422_),
    .X(_0685_));
 sky130_fd_sc_hd__o211a_1 _1236_ (.A1(\stack[12] ),
    .A2(_0423_),
    .B1(net23),
    .C1(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _1237_ (.A0(\stack[12] ),
    .A1(\stack[10] ),
    .S(net19),
    .X(_0687_));
 sky130_fd_sc_hd__a211o_1 _1238_ (.A1(net21),
    .A2(_0687_),
    .B1(_0686_),
    .C1(_0672_),
    .X(_0688_));
 sky130_fd_sc_hd__o211a_1 _1239_ (.A1(net252),
    .A2(_0671_),
    .B1(_0688_),
    .C1(net59),
    .X(_0159_));
 sky130_fd_sc_hd__or2_1 _1240_ (.A(\stack[9] ),
    .B(_0422_),
    .X(_0689_));
 sky130_fd_sc_hd__o211a_1 _1241_ (.A1(\stack[11] ),
    .A2(_0423_),
    .B1(net23),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _1242_ (.A0(\stack[11] ),
    .A1(\stack[9] ),
    .S(net19),
    .X(_0691_));
 sky130_fd_sc_hd__a211o_1 _1243_ (.A1(net21),
    .A2(_0691_),
    .B1(_0690_),
    .C1(net13),
    .X(_0692_));
 sky130_fd_sc_hd__o211a_1 _1244_ (.A1(net251),
    .A2(_0671_),
    .B1(_0692_),
    .C1(net59),
    .X(_0158_));
 sky130_fd_sc_hd__or2_1 _1245_ (.A(\stack[8] ),
    .B(_0422_),
    .X(_0693_));
 sky130_fd_sc_hd__o211a_1 _1246_ (.A1(\stack[10] ),
    .A2(_0423_),
    .B1(net23),
    .C1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _1247_ (.A0(\stack[10] ),
    .A1(\stack[8] ),
    .S(net19),
    .X(_0695_));
 sky130_fd_sc_hd__a211o_1 _1248_ (.A1(net21),
    .A2(_0695_),
    .B1(_0694_),
    .C1(net13),
    .X(_0696_));
 sky130_fd_sc_hd__o211a_1 _1249_ (.A1(net247),
    .A2(net14),
    .B1(_0696_),
    .C1(net59),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _1250_ (.A(\stack[7] ),
    .B(net26),
    .X(_0697_));
 sky130_fd_sc_hd__o211a_1 _1251_ (.A1(\stack[9] ),
    .A2(net25),
    .B1(net24),
    .C1(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _1252_ (.A0(\stack[9] ),
    .A1(\stack[7] ),
    .S(net19),
    .X(_0699_));
 sky130_fd_sc_hd__a211o_1 _1253_ (.A1(net21),
    .A2(_0699_),
    .B1(_0698_),
    .C1(net13),
    .X(_0700_));
 sky130_fd_sc_hd__o211a_1 _1254_ (.A1(net245),
    .A2(net14),
    .B1(_0700_),
    .C1(net59),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _1255_ (.A(\stack[6] ),
    .B(net26),
    .X(_0701_));
 sky130_fd_sc_hd__o211a_1 _1256_ (.A1(\stack[8] ),
    .A2(net25),
    .B1(net23),
    .C1(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _1257_ (.A0(\stack[8] ),
    .A1(\stack[6] ),
    .S(net19),
    .X(_0703_));
 sky130_fd_sc_hd__a211o_1 _1258_ (.A1(net22),
    .A2(_0703_),
    .B1(_0702_),
    .C1(_0672_),
    .X(_0704_));
 sky130_fd_sc_hd__o211a_1 _1259_ (.A1(\stack[7] ),
    .A2(_0671_),
    .B1(_0704_),
    .C1(net59),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _1260_ (.A(\stack[5] ),
    .B(net26),
    .X(_0705_));
 sky130_fd_sc_hd__o211a_1 _1261_ (.A1(\stack[7] ),
    .A2(net25),
    .B1(net24),
    .C1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _1262_ (.A0(\stack[7] ),
    .A1(\stack[5] ),
    .S(net19),
    .X(_0707_));
 sky130_fd_sc_hd__a211o_1 _1263_ (.A1(net22),
    .A2(_0707_),
    .B1(_0706_),
    .C1(_0672_),
    .X(_0708_));
 sky130_fd_sc_hd__o211a_1 _1264_ (.A1(\stack[6] ),
    .A2(_0671_),
    .B1(_0708_),
    .C1(net60),
    .X(_0154_));
 sky130_fd_sc_hd__or2_1 _1265_ (.A(\stack[4] ),
    .B(net26),
    .X(_0709_));
 sky130_fd_sc_hd__o211a_1 _1266_ (.A1(\stack[6] ),
    .A2(net25),
    .B1(net24),
    .C1(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _1267_ (.A0(\stack[6] ),
    .A1(\stack[4] ),
    .S(net19),
    .X(_0711_));
 sky130_fd_sc_hd__a211o_1 _1268_ (.A1(net22),
    .A2(_0711_),
    .B1(_0710_),
    .C1(_0672_),
    .X(_0712_));
 sky130_fd_sc_hd__o211a_1 _1269_ (.A1(\stack[5] ),
    .A2(net14),
    .B1(_0712_),
    .C1(net60),
    .X(_0153_));
 sky130_fd_sc_hd__or2_1 _1270_ (.A(\stack[3] ),
    .B(net26),
    .X(_0713_));
 sky130_fd_sc_hd__o211a_1 _1271_ (.A1(\stack[5] ),
    .A2(net25),
    .B1(net23),
    .C1(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _1272_ (.A0(\stack[5] ),
    .A1(\stack[3] ),
    .S(net20),
    .X(_0715_));
 sky130_fd_sc_hd__a211o_1 _1273_ (.A1(net21),
    .A2(_0715_),
    .B1(_0714_),
    .C1(net13),
    .X(_0716_));
 sky130_fd_sc_hd__o211a_1 _1274_ (.A1(net264),
    .A2(net14),
    .B1(_0716_),
    .C1(net60),
    .X(_0152_));
 sky130_fd_sc_hd__or2_1 _1275_ (.A(\stack[2] ),
    .B(_0422_),
    .X(_0717_));
 sky130_fd_sc_hd__o211a_1 _1276_ (.A1(\stack[4] ),
    .A2(net25),
    .B1(net23),
    .C1(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _1277_ (.A0(\stack[4] ),
    .A1(\stack[2] ),
    .S(net19),
    .X(_0719_));
 sky130_fd_sc_hd__a211o_1 _1278_ (.A1(net21),
    .A2(_0719_),
    .B1(_0718_),
    .C1(net13),
    .X(_0720_));
 sky130_fd_sc_hd__o211a_1 _1279_ (.A1(\stack[3] ),
    .A2(net14),
    .B1(_0720_),
    .C1(net59),
    .X(_0151_));
 sky130_fd_sc_hd__or2_1 _1280_ (.A(\stack[1] ),
    .B(net26),
    .X(_0721_));
 sky130_fd_sc_hd__o211a_1 _1281_ (.A1(\stack[3] ),
    .A2(net25),
    .B1(net23),
    .C1(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(\stack[3] ),
    .A1(\stack[1] ),
    .S(net20),
    .X(_0723_));
 sky130_fd_sc_hd__a211o_1 _1283_ (.A1(net21),
    .A2(_0723_),
    .B1(_0722_),
    .C1(net13),
    .X(_0724_));
 sky130_fd_sc_hd__o211a_1 _1284_ (.A1(\stack[2] ),
    .A2(net14),
    .B1(_0724_),
    .C1(net59),
    .X(_0150_));
 sky130_fd_sc_hd__o211a_1 _1285_ (.A1(\stack[2] ),
    .A2(net25),
    .B1(_0424_),
    .C1(net24),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _1286_ (.A0(\stack[0] ),
    .A1(\stack[2] ),
    .S(_0417_),
    .X(_0287_));
 sky130_fd_sc_hd__a211o_1 _1287_ (.A1(net22),
    .A2(_0287_),
    .B1(_0286_),
    .C1(net13),
    .X(_0288_));
 sky130_fd_sc_hd__o211a_1 _1288_ (.A1(\stack[1] ),
    .A2(net14),
    .B1(_0288_),
    .C1(net58),
    .X(_0149_));
 sky130_fd_sc_hd__or4_1 _1289_ (.A(net36),
    .B(_0373_),
    .C(_0414_),
    .D(_0447_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(net47),
    .A1(net244),
    .S(_0289_),
    .X(_0148_));
 sky130_fd_sc_hd__and4bb_2 _1291_ (.A_N(net43),
    .B_N(_0414_),
    .C(_0417_),
    .D(net39),
    .X(_0290_));
 sky130_fd_sc_hd__or3b_1 _1292_ (.A(_0550_),
    .B(_0560_),
    .C_N(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__a21o_1 _1293_ (.A1(_0549_),
    .A2(_0290_),
    .B1(uo_out[3]),
    .X(_0292_));
 sky130_fd_sc_hd__and3_1 _1294_ (.A(net58),
    .B(_0291_),
    .C(_0292_),
    .X(_0147_));
 sky130_fd_sc_hd__nand2_1 _1295_ (.A(_0552_),
    .B(_0290_),
    .Y(_0293_));
 sky130_fd_sc_hd__a21o_1 _1296_ (.A1(_0552_),
    .A2(_0290_),
    .B1(uo_out[2]),
    .X(_0294_));
 sky130_fd_sc_hd__o211a_1 _1297_ (.A1(_0560_),
    .A2(_0293_),
    .B1(_0294_),
    .C1(net58),
    .X(_0146_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0553_),
    .B(_0290_),
    .Y(_0295_));
 sky130_fd_sc_hd__a21o_1 _1299_ (.A1(_0553_),
    .A2(_0290_),
    .B1(uo_out[1]),
    .X(_0296_));
 sky130_fd_sc_hd__o211a_1 _1300_ (.A1(_0560_),
    .A2(_0295_),
    .B1(_0296_),
    .C1(net60),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_1 _1301_ (.A(_0555_),
    .B(_0290_),
    .Y(_0297_));
 sky130_fd_sc_hd__a21o_1 _1302_ (.A1(_0555_),
    .A2(_0290_),
    .B1(uo_out[0]),
    .X(_0298_));
 sky130_fd_sc_hd__o211a_1 _1303_ (.A1(_0560_),
    .A2(_0297_),
    .B1(_0298_),
    .C1(net60),
    .X(_0144_));
 sky130_fd_sc_hd__mux4_1 _1304_ (.A0(\stack[7] ),
    .A1(\stack[6] ),
    .A2(\stack[5] ),
    .A3(\stack[4] ),
    .S0(\fetch_count[0] ),
    .S1(\fetch_count[1] ),
    .X(_0299_));
 sky130_fd_sc_hd__mux4_1 _1305_ (.A0(\stack[3] ),
    .A1(\stack[2] ),
    .A2(\stack[1] ),
    .A3(\stack[0] ),
    .S0(\fetch_count[0] ),
    .S1(\fetch_count[1] ),
    .X(_0300_));
 sky130_fd_sc_hd__or2_1 _1306_ (.A(_0319_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_1 _1307_ (.A1(\fetch_count[2] ),
    .A2(_0299_),
    .B1(_0301_),
    .C1(net54),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_2 _1308_ (.A(eeprom_cs),
    .B(net68),
    .Y(eeprom_sck));
 sky130_fd_sc_hd__inv_2 _1310__4 (.A(clknet_4_13_0_clk),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _1311__5 (.A(clknet_4_7_0_clk),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _1312__6 (.A(clknet_4_7_0_clk),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _1313__7 (.A(clknet_4_6_0_clk),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _1314__8 (.A(clknet_4_13_0_clk),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _1315__9 (.A(clknet_4_13_0_clk),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _1316__10 (.A(clknet_4_13_0_clk),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _1317__11 (.A(clknet_4_15_0_clk),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _1318__12 (.A(clknet_4_15_0_clk),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _1319__13 (.A(clknet_4_15_0_clk),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _1320__14 (.A(clknet_4_15_0_clk),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _1321__15 (.A(clknet_4_15_0_clk),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _1322__16 (.A(clknet_4_14_0_clk),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _1323__17 (.A(clknet_4_14_0_clk),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _1324__18 (.A(clknet_4_14_0_clk),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _1325__19 (.A(clknet_4_14_0_clk),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _1326__20 (.A(clknet_4_14_0_clk),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _1327__21 (.A(clknet_4_12_0_clk),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _1328__22 (.A(clknet_4_13_0_clk),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _1329__23 (.A(clknet_4_5_0_clk),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _1330__24 (.A(clknet_4_3_0_clk),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _1331__25 (.A(clknet_4_5_0_clk),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _1332__26 (.A(clknet_4_6_0_clk),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _1333__27 (.A(clknet_4_7_0_clk),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _1334__28 (.A(clknet_4_5_0_clk),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _1335__29 (.A(clknet_4_7_0_clk),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _1336__30 (.A(clknet_4_5_0_clk),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _1337__31 (.A(clknet_4_5_0_clk),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _1338__32 (.A(clknet_4_5_0_clk),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _1339__33 (.A(clknet_4_4_0_clk),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _1340__34 (.A(clknet_4_4_0_clk),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _1341__35 (.A(clknet_4_4_0_clk),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _1342__36 (.A(clknet_4_4_0_clk),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _1343__37 (.A(clknet_4_9_0_clk),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _1344__38 (.A(clknet_4_11_0_clk),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _1345__39 (.A(clknet_4_11_0_clk),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _1346__40 (.A(clknet_4_11_0_clk),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _1347__41 (.A(clknet_4_14_0_clk),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _1348__42 (.A(clknet_4_14_0_clk),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _1349__43 (.A(clknet_4_14_0_clk),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _1350__44 (.A(clknet_4_14_0_clk),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _1351__45 (.A(clknet_4_7_0_clk),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _1352__46 (.A(clknet_4_7_0_clk),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _1353__47 (.A(clknet_4_7_0_clk),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _1354__48 (.A(clknet_4_7_0_clk),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _1355__49 (.A(clknet_4_5_0_clk),
    .Y(net115));
 sky130_fd_sc_hd__inv_2 _1356__50 (.A(clknet_4_5_0_clk),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _1357__51 (.A(clknet_4_5_0_clk),
    .Y(net117));
 sky130_fd_sc_hd__inv_2 _1358__52 (.A(clknet_4_5_0_clk),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _1359__53 (.A(clknet_4_5_0_clk),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _1360__54 (.A(clknet_4_4_0_clk),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _1361__55 (.A(clknet_4_4_0_clk),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _1362__56 (.A(clknet_4_4_0_clk),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _1363__57 (.A(clknet_4_4_0_clk),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _1364__58 (.A(clknet_4_9_0_clk),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _1365__59 (.A(clknet_4_11_0_clk),
    .Y(net125));
 sky130_fd_sc_hd__inv_2 _1366__60 (.A(clknet_4_11_0_clk),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _1367__61 (.A(clknet_4_9_0_clk),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _1368__62 (.A(clknet_4_12_0_clk),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _1369__63 (.A(clknet_4_9_0_clk),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _1370__64 (.A(clknet_4_12_0_clk),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _1371__65 (.A(clknet_4_12_0_clk),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _1372__66 (.A(clknet_4_13_0_clk),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _1373__67 (.A(clknet_4_6_0_clk),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _1374__68 (.A(clknet_4_6_0_clk),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _1375__69 (.A(clknet_4_13_0_clk),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _1376__70 (.A(clknet_4_6_0_clk),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _1377__71 (.A(clknet_4_6_0_clk),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _1378__72 (.A(clknet_4_6_0_clk),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _1379__73 (.A(clknet_4_6_0_clk),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _1380__74 (.A(clknet_4_12_0_clk),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _1381__75 (.A(clknet_4_11_0_clk),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _1382__76 (.A(clknet_4_11_0_clk),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _1383__77 (.A(clknet_4_11_0_clk),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _1384__78 (.A(clknet_4_11_0_clk),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _1385__79 (.A(clknet_4_10_0_clk),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _1386__80 (.A(clknet_4_10_0_clk),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _1387__81 (.A(clknet_4_10_0_clk),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _1388__82 (.A(clknet_4_10_0_clk),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _1389__83 (.A(clknet_4_10_0_clk),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _1390__84 (.A(clknet_4_10_0_clk),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _1391__85 (.A(clknet_4_10_0_clk),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _1392__86 (.A(clknet_4_10_0_clk),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _1393__87 (.A(clknet_4_8_0_clk),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _1394__88 (.A(clknet_4_8_0_clk),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _1395__89 (.A(clknet_4_8_0_clk),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _1396__90 (.A(clknet_4_8_0_clk),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _1397__91 (.A(clknet_4_8_0_clk),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _1398__92 (.A(clknet_4_8_0_clk),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _1399__93 (.A(clknet_4_8_0_clk),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _1400__94 (.A(clknet_4_8_0_clk),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _1401__95 (.A(clknet_4_2_0_clk),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _1402__96 (.A(clknet_4_2_0_clk),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _1403__97 (.A(clknet_4_2_0_clk),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _1404__98 (.A(clknet_4_2_0_clk),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _1405__99 (.A(clknet_4_2_0_clk),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _1406__100 (.A(clknet_4_2_0_clk),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _1407__101 (.A(clknet_4_0_0_clk),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _1408__102 (.A(clknet_4_0_0_clk),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _1409__103 (.A(clknet_4_0_0_clk),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _1410__104 (.A(clknet_4_0_0_clk),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _1411__105 (.A(clknet_4_0_0_clk),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _1412__106 (.A(clknet_4_0_0_clk),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _1413__107 (.A(clknet_4_11_0_clk),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _1414__108 (.A(clknet_4_10_0_clk),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _1415__109 (.A(clknet_4_10_0_clk),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _1416__110 (.A(clknet_4_8_0_clk),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _1417__111 (.A(clknet_4_12_0_clk),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _1418__112 (.A(clknet_4_9_0_clk),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _1419__113 (.A(clknet_4_9_0_clk),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _1420__114 (.A(clknet_4_8_0_clk),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _1421__115 (.A(clknet_4_3_0_clk),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _1422__116 (.A(clknet_4_9_0_clk),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _1423__117 (.A(clknet_4_9_0_clk),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _1424__118 (.A(clknet_4_9_0_clk),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _1425__119 (.A(clknet_4_2_0_clk),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _1426__120 (.A(clknet_4_8_0_clk),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _1427__121 (.A(clknet_4_2_0_clk),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _1428__122 (.A(clknet_4_2_0_clk),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _1429__123 (.A(clknet_4_3_0_clk),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _1430__124 (.A(clknet_4_3_0_clk),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _1431__125 (.A(clknet_4_3_0_clk),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _1432__126 (.A(clknet_4_3_0_clk),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _1433__127 (.A(clknet_4_12_0_clk),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _1434__128 (.A(clknet_4_3_0_clk),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _1435__129 (.A(clknet_4_3_0_clk),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _1436__130 (.A(clknet_4_1_0_clk),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _1437__131 (.A(clknet_4_1_0_clk),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _1438__132 (.A(clknet_4_1_0_clk),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _1439__133 (.A(clknet_4_1_0_clk),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _1440__134 (.A(clknet_4_1_0_clk),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _1441__135 (.A(clknet_4_1_0_clk),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _1442__136 (.A(clknet_4_1_0_clk),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _1443__137 (.A(clknet_4_0_0_clk),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _1444__138 (.A(clknet_4_0_0_clk),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _1445__139 (.A(clknet_4_0_0_clk),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _1446__140 (.A(clknet_4_0_0_clk),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _1447__141 (.A(clknet_4_1_0_clk),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _1448__142 (.A(clknet_4_1_0_clk),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _1449__143 (.A(clknet_4_1_0_clk),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _1450__144 (.A(clknet_4_1_0_clk),
    .Y(net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(net67),
    .D(_0143_),
    .Q(stack_out));
 sky130_fd_sc_hd__dfxtp_4 _1452_ (.CLK(net69),
    .D(_0144_),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_4 _1453_ (.CLK(net70),
    .D(_0145_),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_4 _1454_ (.CLK(net71),
    .D(_0146_),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_4 _1455_ (.CLK(net72),
    .D(_0147_),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_1 _1456_ (.CLK(net73),
    .D(_0148_),
    .Q(timer_mode));
 sky130_fd_sc_hd__dfxtp_1 _1457_ (.CLK(net74),
    .D(_0149_),
    .Q(\stack[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1458_ (.CLK(net75),
    .D(_0150_),
    .Q(\stack[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1459_ (.CLK(net76),
    .D(_0151_),
    .Q(\stack[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1460_ (.CLK(net77),
    .D(_0152_),
    .Q(\stack[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1461_ (.CLK(net78),
    .D(_0153_),
    .Q(\stack[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1462_ (.CLK(net79),
    .D(_0154_),
    .Q(\stack[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1463_ (.CLK(net80),
    .D(_0155_),
    .Q(\stack[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1464_ (.CLK(net81),
    .D(_0156_),
    .Q(\stack[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1465_ (.CLK(net82),
    .D(_0157_),
    .Q(\stack[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1466_ (.CLK(net83),
    .D(_0158_),
    .Q(\stack[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1467_ (.CLK(net84),
    .D(_0159_),
    .Q(\stack[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1468_ (.CLK(net85),
    .D(_0160_),
    .Q(\stack[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1469_ (.CLK(net86),
    .D(_0161_),
    .Q(\stack[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1470_ (.CLK(net87),
    .D(_0162_),
    .Q(\stack[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1471_ (.CLK(net88),
    .D(_0163_),
    .Q(\stack[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1472_ (.CLK(net89),
    .D(_0164_),
    .Q(eeprom_copi));
 sky130_fd_sc_hd__dfxtp_1 _1473_ (.CLK(net90),
    .D(_0165_),
    .Q(timer_out));
 sky130_fd_sc_hd__dfxtp_1 _1474_ (.CLK(net91),
    .D(_0166_),
    .Q(eeprom_cs));
 sky130_fd_sc_hd__dfxtp_1 _1475_ (.CLK(clknet_4_13_0_clk),
    .D(net10),
    .Q(\uio_in_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1476_ (.CLK(clknet_4_15_0_clk),
    .D(net2),
    .Q(\ui_in_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1477_ (.CLK(clknet_4_15_0_clk),
    .D(net3),
    .Q(\ui_in_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1478_ (.CLK(clknet_4_15_0_clk),
    .D(net4),
    .Q(\ui_in_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1479_ (.CLK(clknet_4_15_0_clk),
    .D(net5),
    .Q(\ui_in_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1480_ (.CLK(clknet_4_15_0_clk),
    .D(net6),
    .Q(\ui_in_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1481_ (.CLK(clknet_4_15_0_clk),
    .D(net7),
    .Q(\ui_in_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1482_ (.CLK(clknet_4_15_0_clk),
    .D(net8),
    .Q(\ui_in_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1483_ (.CLK(clknet_4_15_0_clk),
    .D(net9),
    .Q(\ui_in_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1484_ (.CLK(net92),
    .D(_0167_),
    .Q(\fetch_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1485_ (.CLK(net93),
    .D(_0168_),
    .Q(\fetch_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1486_ (.CLK(net94),
    .D(_0169_),
    .Q(\fetch_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1487_ (.CLK(net95),
    .D(_0170_),
    .Q(\fetch_state[3] ));
 sky130_fd_sc_hd__dfxtp_4 _1488_ (.CLK(net96),
    .D(_0171_),
    .Q(\fetch_count[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1489_ (.CLK(net97),
    .D(_0172_),
    .Q(\fetch_count[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1490_ (.CLK(net98),
    .D(_0173_),
    .Q(\fetch_count[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1491_ (.CLK(net99),
    .D(_0174_),
    .Q(\fetch_prev_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1492_ (.CLK(net100),
    .D(_0175_),
    .Q(\fetch_prev_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1493_ (.CLK(net101),
    .D(net214),
    .Q(\fetch_prev_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1494_ (.CLK(net102),
    .D(_0177_),
    .Q(\fetch_prev_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1495_ (.CLK(net103),
    .D(_0178_),
    .Q(\cur_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1496_ (.CLK(net104),
    .D(_0179_),
    .Q(\cur_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1497_ (.CLK(net105),
    .D(_0180_),
    .Q(\cur_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1498_ (.CLK(net106),
    .D(_0181_),
    .Q(\cur_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1499_ (.CLK(net107),
    .D(_0182_),
    .Q(\cur_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1500_ (.CLK(net108),
    .D(_0183_),
    .Q(\cur_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1501_ (.CLK(net109),
    .D(_0184_),
    .Q(\cur_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1502_ (.CLK(net110),
    .D(_0185_),
    .Q(\cur_addr[7] ));
 sky130_fd_sc_hd__dfxtp_4 _1503_ (.CLK(net111),
    .D(_0186_),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_4 _1504_ (.CLK(net112),
    .D(_0187_),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_4 _1505_ (.CLK(net113),
    .D(_0188_),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_4 _1506_ (.CLK(net114),
    .D(_0189_),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfxtp_1 _1507_ (.CLK(net115),
    .D(_0190_),
    .Q(eeprom_oe_copi));
 sky130_fd_sc_hd__dfxtp_1 _1508_ (.CLK(net116),
    .D(_0191_),
    .Q(\cycle_start_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1509_ (.CLK(net117),
    .D(_0192_),
    .Q(\cycle_start_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1510_ (.CLK(net118),
    .D(_0193_),
    .Q(\cycle_start_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1511_ (.CLK(net119),
    .D(_0194_),
    .Q(\cycle_start_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1512_ (.CLK(net120),
    .D(_0195_),
    .Q(\cycle_start_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1513_ (.CLK(net121),
    .D(_0196_),
    .Q(\cycle_start_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1514_ (.CLK(net122),
    .D(_0197_),
    .Q(\cycle_start_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1515_ (.CLK(net123),
    .D(_0198_),
    .Q(\cycle_start_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1516_ (.CLK(net124),
    .D(_0199_),
    .Q(\cycle_end_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1517_ (.CLK(net125),
    .D(_0200_),
    .Q(\cycle_end_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1518_ (.CLK(net126),
    .D(_0201_),
    .Q(\cycle_end_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1519_ (.CLK(net127),
    .D(_0202_),
    .Q(\cycle_end_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1520_ (.CLK(net128),
    .D(_0203_),
    .Q(\cycle_end_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1521_ (.CLK(net129),
    .D(_0204_),
    .Q(\cycle_end_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1522_ (.CLK(net130),
    .D(_0205_),
    .Q(\cycle_end_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1523_ (.CLK(net131),
    .D(_0206_),
    .Q(\cycle_end_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1524_ (.CLK(net132),
    .D(_0207_),
    .Q(\instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1525_ (.CLK(net133),
    .D(_0208_),
    .Q(\instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1526_ (.CLK(net134),
    .D(_0209_),
    .Q(\instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1527_ (.CLK(net135),
    .D(_0210_),
    .Q(\instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1528_ (.CLK(net136),
    .D(_0211_),
    .Q(\instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1529_ (.CLK(net137),
    .D(_0212_),
    .Q(\instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1530_ (.CLK(net138),
    .D(_0213_),
    .Q(\instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1531_ (.CLK(net139),
    .D(_0214_),
    .Q(\instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1532_ (.CLK(net140),
    .D(_0215_),
    .Q(\stack[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1533_ (.CLK(net141),
    .D(_0216_),
    .Q(\timer_clock_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1534_ (.CLK(net142),
    .D(net240),
    .Q(\timer_clock_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1535_ (.CLK(net143),
    .D(_0218_),
    .Q(\timer_clock_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1536_ (.CLK(net144),
    .D(_0219_),
    .Q(\timer_clock_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1537_ (.CLK(net145),
    .D(_0220_),
    .Q(\timer_clock_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1538_ (.CLK(net146),
    .D(_0221_),
    .Q(\timer_clock_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1539_ (.CLK(net147),
    .D(_0222_),
    .Q(\timer_clock_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1540_ (.CLK(net148),
    .D(_0223_),
    .Q(\timer_clock_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1541_ (.CLK(net149),
    .D(_0224_),
    .Q(\timer_clock_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1542_ (.CLK(net150),
    .D(_0225_),
    .Q(\timer_clock_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1543_ (.CLK(net151),
    .D(_0226_),
    .Q(\timer_clock_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1544_ (.CLK(net152),
    .D(_0227_),
    .Q(\timer_clock_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1545_ (.CLK(net153),
    .D(_0228_),
    .Q(\timer_clock_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1546_ (.CLK(net154),
    .D(_0229_),
    .Q(\timer_clock_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1547_ (.CLK(net155),
    .D(_0230_),
    .Q(\timer_clock_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1548_ (.CLK(net156),
    .D(_0231_),
    .Q(\timer_clock_counter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1549_ (.CLK(net157),
    .D(_0232_),
    .Q(\timer_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1550_ (.CLK(net158),
    .D(_0233_),
    .Q(\timer_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1551_ (.CLK(net159),
    .D(_0234_),
    .Q(\timer_counter[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1552_ (.CLK(net160),
    .D(_0235_),
    .Q(\timer_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1553_ (.CLK(net161),
    .D(_0236_),
    .Q(\timer_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1554_ (.CLK(net162),
    .D(_0237_),
    .Q(\timer_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1555_ (.CLK(net163),
    .D(_0238_),
    .Q(\timer_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1556_ (.CLK(net164),
    .D(_0239_),
    .Q(\timer_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1557_ (.CLK(net165),
    .D(_0240_),
    .Q(\timer_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1558_ (.CLK(net166),
    .D(_0241_),
    .Q(\timer_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1559_ (.CLK(net167),
    .D(_0242_),
    .Q(\timer_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1560_ (.CLK(net168),
    .D(_0243_),
    .Q(\timer_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1561_ (.CLK(net169),
    .D(_0244_),
    .Q(\timer_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1562_ (.CLK(net170),
    .D(_0245_),
    .Q(\timer_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1563_ (.CLK(net171),
    .D(_0246_),
    .Q(\timer_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1564_ (.CLK(net172),
    .D(_0247_),
    .Q(\timer_counter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1565_ (.CLK(net173),
    .D(_0248_),
    .Q(\timer_clock_divisor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1566_ (.CLK(net174),
    .D(_0249_),
    .Q(\timer_clock_divisor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1567_ (.CLK(net175),
    .D(_0250_),
    .Q(\timer_clock_divisor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1568_ (.CLK(net176),
    .D(_0251_),
    .Q(\timer_clock_divisor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1569_ (.CLK(net177),
    .D(_0252_),
    .Q(\timer_period_a[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1570_ (.CLK(net178),
    .D(_0253_),
    .Q(\timer_period_a[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1571_ (.CLK(net179),
    .D(_0254_),
    .Q(\timer_period_a[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1572_ (.CLK(net180),
    .D(_0255_),
    .Q(\timer_period_a[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1573_ (.CLK(net181),
    .D(_0256_),
    .Q(\timer_period_a[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1574_ (.CLK(net182),
    .D(_0257_),
    .Q(\timer_period_a[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1575_ (.CLK(net183),
    .D(_0258_),
    .Q(\timer_period_a[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1576_ (.CLK(net184),
    .D(_0259_),
    .Q(\timer_period_a[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1577_ (.CLK(net185),
    .D(_0260_),
    .Q(\timer_period_a[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1578_ (.CLK(net186),
    .D(_0261_),
    .Q(\timer_period_a[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1579_ (.CLK(net187),
    .D(_0262_),
    .Q(\timer_period_a[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1580_ (.CLK(net188),
    .D(_0263_),
    .Q(\timer_period_a[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1581_ (.CLK(net189),
    .D(_0264_),
    .Q(\timer_period_a[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1582_ (.CLK(net190),
    .D(_0265_),
    .Q(\timer_period_a[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1583_ (.CLK(net191),
    .D(_0266_),
    .Q(\timer_period_a[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1584_ (.CLK(net192),
    .D(_0267_),
    .Q(\timer_period_a[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1585_ (.CLK(net193),
    .D(_0268_),
    .Q(timer_enabled));
 sky130_fd_sc_hd__dfxtp_1 _1586_ (.CLK(net194),
    .D(_0269_),
    .Q(timer_phase));
 sky130_fd_sc_hd__dfxtp_1 _1587_ (.CLK(net195),
    .D(_0270_),
    .Q(\timer_period_b[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1588_ (.CLK(net196),
    .D(_0271_),
    .Q(\timer_period_b[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1589_ (.CLK(net197),
    .D(_0272_),
    .Q(\timer_period_b[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1590_ (.CLK(net198),
    .D(_0273_),
    .Q(\timer_period_b[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1591_ (.CLK(net199),
    .D(_0274_),
    .Q(\timer_period_b[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1592_ (.CLK(net200),
    .D(_0275_),
    .Q(\timer_period_b[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1593_ (.CLK(net201),
    .D(_0276_),
    .Q(\timer_period_b[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1594_ (.CLK(net202),
    .D(_0277_),
    .Q(\timer_period_b[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1595_ (.CLK(net203),
    .D(_0278_),
    .Q(\timer_period_b[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1596_ (.CLK(net204),
    .D(_0279_),
    .Q(\timer_period_b[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1597_ (.CLK(net205),
    .D(_0280_),
    .Q(\timer_period_b[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1598_ (.CLK(net206),
    .D(_0281_),
    .Q(\timer_period_b[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1599_ (.CLK(net207),
    .D(_0282_),
    .Q(\timer_period_b[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1600_ (.CLK(net208),
    .D(_0283_),
    .Q(\timer_period_b[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1601_ (.CLK(net209),
    .D(_0284_),
    .Q(\timer_period_b[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1602_ (.CLK(net210),
    .D(_0285_),
    .Q(\timer_period_b[15] ));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_66 (.LO(net66));
 sky130_fd_sc_hd__inv_2 _0753__1 (.A(clknet_4_7_0_clk),
    .Y(net67));
 sky130_fd_sc_hd__buf_2 _1609_ (.A(eeprom_oe_copi),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__buf_2 _1610_ (.A(eeprom_oe_copi),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__buf_2 _1611_ (.A(eeprom_oe_copi),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__buf_2 _1612_ (.A(eeprom_oe_copi),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__buf_2 _1613_ (.A(eeprom_oe_copi),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__buf_2 _1614_ (.A(eeprom_sck),
    .X(uio_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _1615_ (.A(eeprom_cs),
    .X(uio_out[1]));
 sky130_fd_sc_hd__clkbuf_4 _1616_ (.A(eeprom_copi),
    .X(uio_out[2]));
 sky130_fd_sc_hd__clkbuf_4 _1617_ (.A(stack_out),
    .X(uio_out[6]));
 sky130_fd_sc_hd__buf_2 _1618_ (.A(timer_out),
    .X(uio_out[7]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(_0468_),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout12 (.A(_0468_),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(_0672_),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(_0671_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(_0496_),
    .X(net15));
 sky130_fd_sc_hd__buf_1 fanout16 (.A(_0496_),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 max_cap17 (.A(_0366_),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(_0520_),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(_0418_),
    .X(net20));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(_0562_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(_0561_),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(_0423_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(_0422_),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(timer_enabled),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 fanout30 (.A(timer_enabled),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(net33),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(\instr[7] ),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(\instr[6] ),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(\instr[5] ),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(\instr[4] ),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net41),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(\instr[3] ),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 fanout44 (.A(\instr[2] ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(\instr[1] ),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(\instr[0] ),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(\fetch_state[3] ),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__buf_1 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net54),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(net1),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net57),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net1),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net60),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 fanout60 (.A(net1),
    .X(net60));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_61 (.LO(net61));
 sky130_fd_sc_hd__inv_2 _0753__2 (.A(clknet_4_7_0_clk),
    .Y(net68));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__inv_2 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_4 clkload1 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_2 clkload5 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__inv_4 clkload6 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__inv_2 clkload7 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__inv_2 clkload8 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_8 clkload9 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload10 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__inv_4 clkload11 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\timer_clock_counter[15] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(eeprom_copi),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\fetch_prev_state[2] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0176_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\timer_clock_counter[13] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\timer_clock_counter[10] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\fetch_prev_state[3] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\timer_clock_counter[8] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\timer_clock_counter[6] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\timer_counter[3] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\timer_clock_counter[4] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(eeprom_cs),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\cur_addr[7] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(eeprom_oe_copi),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\timer_period_a[4] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\timer_period_a[12] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\timer_clock_counter[7] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\timer_period_b[12] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\cur_addr[3] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0587_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(timer_phase),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\cur_addr[4] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\timer_clock_counter[9] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\cur_addr[6] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0585_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\timer_clock_counter[12] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\stack[14] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\cycle_end_addr[0] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\timer_clock_counter[0] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0217_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\timer_period_b[4] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\cur_addr[5] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\cur_addr[2] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(timer_mode),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\stack[8] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\cur_addr[0] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\stack[9] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\fetch_state[1] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\stack[13] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\timer_counter[12] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\stack[10] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\stack[11] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\cycle_end_addr[1] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\cycle_start_addr[0] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\cycle_start_addr[2] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\cycle_start_addr[4] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\cycle_start_addr[7] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\fetch_prev_state[0] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\stack[12] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\cycle_start_addr[6] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\cycle_end_addr[6] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\cycle_start_addr[5] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\cycle_start_addr[1] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\stack[4] ),
    .X(net264));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_331 ();
 assign uio_oe[3] = net61;
 assign uio_oe[4] = net62;
 assign uio_oe[5] = net63;
 assign uio_out[3] = net64;
 assign uio_out[4] = net65;
 assign uio_out[5] = net66;
endmodule
