VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.150 BY 17.150 ;
  OBS
      LAYER met1 ;
        RECT 0.000 16.800 17.150 17.150 ;
        RECT 0.000 16.100 2.100 16.800 ;
      LAYER met1 ;
        RECT 2.100 16.100 3.850 16.800 ;
      LAYER met1 ;
        RECT 3.850 16.100 5.600 16.800 ;
      LAYER met1 ;
        RECT 5.600 16.100 6.650 16.800 ;
      LAYER met1 ;
        RECT 6.650 16.100 8.400 16.800 ;
      LAYER met1 ;
        RECT 8.400 16.100 10.150 16.800 ;
      LAYER met1 ;
        RECT 10.150 16.100 11.200 16.800 ;
        RECT 0.000 15.400 1.750 16.100 ;
      LAYER met1 ;
        RECT 1.750 15.750 4.200 16.100 ;
        RECT 1.750 15.400 2.450 15.750 ;
      LAYER met1 ;
        RECT 2.450 15.400 3.150 15.750 ;
        RECT 0.000 14.700 3.150 15.400 ;
      LAYER met1 ;
        RECT 3.150 14.700 4.200 15.750 ;
      LAYER met1 ;
        RECT 4.200 15.400 5.250 16.100 ;
      LAYER met1 ;
        RECT 5.250 15.750 7.000 16.100 ;
      LAYER met1 ;
        RECT 7.000 15.750 8.050 16.100 ;
      LAYER met1 ;
        RECT 8.050 15.750 10.500 16.100 ;
        RECT 5.250 15.400 5.950 15.750 ;
      LAYER met1 ;
        RECT 4.200 14.700 4.900 15.400 ;
        RECT 0.000 14.350 2.800 14.700 ;
      LAYER met1 ;
        RECT 2.800 14.350 3.850 14.700 ;
      LAYER met1 ;
        RECT 0.000 13.650 2.450 14.350 ;
      LAYER met1 ;
        RECT 2.450 14.000 3.850 14.350 ;
      LAYER met1 ;
        RECT 3.850 14.000 4.900 14.700 ;
      LAYER met1 ;
        RECT 2.450 13.650 3.500 14.000 ;
      LAYER met1 ;
        RECT 3.500 13.650 4.900 14.000 ;
      LAYER met1 ;
        RECT 4.900 13.650 5.950 15.400 ;
      LAYER met1 ;
        RECT 0.000 12.950 2.100 13.650 ;
      LAYER met1 ;
        RECT 2.100 12.950 3.150 13.650 ;
      LAYER met1 ;
        RECT 3.150 13.300 5.250 13.650 ;
      LAYER met1 ;
        RECT 5.250 13.300 5.950 13.650 ;
      LAYER met1 ;
        RECT 5.950 13.300 6.300 15.750 ;
      LAYER met1 ;
        RECT 6.300 13.300 7.350 15.750 ;
      LAYER met1 ;
        RECT 7.350 15.400 8.050 15.750 ;
      LAYER met1 ;
        RECT 8.050 15.400 8.750 15.750 ;
      LAYER met1 ;
        RECT 8.750 15.400 9.450 15.750 ;
        RECT 7.350 14.700 9.450 15.400 ;
      LAYER met1 ;
        RECT 9.450 14.700 10.500 15.750 ;
      LAYER met1 ;
        RECT 10.500 14.700 11.200 16.100 ;
      LAYER met1 ;
        RECT 11.200 15.750 13.650 16.800 ;
      LAYER met1 ;
        RECT 13.650 15.750 17.150 16.800 ;
      LAYER met1 ;
        RECT 11.200 15.400 12.250 15.750 ;
      LAYER met1 ;
        RECT 12.250 15.400 17.150 15.750 ;
      LAYER met1 ;
        RECT 11.200 15.050 13.300 15.400 ;
      LAYER met1 ;
        RECT 13.300 15.050 17.150 15.400 ;
        RECT 7.350 14.350 9.100 14.700 ;
      LAYER met1 ;
        RECT 9.100 14.350 10.150 14.700 ;
      LAYER met1 ;
        RECT 7.350 13.650 8.750 14.350 ;
      LAYER met1 ;
        RECT 8.750 14.000 10.150 14.350 ;
      LAYER met1 ;
        RECT 10.150 14.000 11.200 14.700 ;
      LAYER met1 ;
        RECT 11.200 14.350 13.650 15.050 ;
        RECT 11.200 14.000 12.250 14.350 ;
      LAYER met1 ;
        RECT 12.250 14.000 12.600 14.350 ;
      LAYER met1 ;
        RECT 12.600 14.000 13.650 14.350 ;
        RECT 8.750 13.650 9.800 14.000 ;
      LAYER met1 ;
        RECT 9.800 13.650 12.950 14.000 ;
      LAYER met1 ;
        RECT 12.950 13.650 13.650 14.000 ;
      LAYER met1 ;
        RECT 7.350 13.300 8.400 13.650 ;
        RECT 3.150 12.950 3.500 13.300 ;
      LAYER met1 ;
        RECT 3.500 12.950 4.200 13.300 ;
      LAYER met1 ;
        RECT 4.200 12.950 5.250 13.300 ;
      LAYER met1 ;
        RECT 5.250 12.950 7.000 13.300 ;
      LAYER met1 ;
        RECT 7.000 12.950 8.400 13.300 ;
      LAYER met1 ;
        RECT 8.400 12.950 9.450 13.650 ;
      LAYER met1 ;
        RECT 9.450 13.300 11.200 13.650 ;
      LAYER met1 ;
        RECT 11.200 13.300 11.900 13.650 ;
      LAYER met1 ;
        RECT 11.900 13.300 12.600 13.650 ;
        RECT 9.450 12.950 9.800 13.300 ;
      LAYER met1 ;
        RECT 9.800 12.950 10.500 13.300 ;
      LAYER met1 ;
        RECT 10.500 12.950 11.200 13.300 ;
      LAYER met1 ;
        RECT 11.200 12.950 12.250 13.300 ;
      LAYER met1 ;
        RECT 12.250 12.950 12.600 13.300 ;
      LAYER met1 ;
        RECT 12.600 12.950 13.650 13.650 ;
      LAYER met1 ;
        RECT 13.650 12.950 17.150 15.050 ;
        RECT 0.000 12.250 1.750 12.950 ;
      LAYER met1 ;
        RECT 1.750 12.250 4.200 12.950 ;
      LAYER met1 ;
        RECT 4.200 12.250 5.600 12.950 ;
      LAYER met1 ;
        RECT 5.600 12.600 7.000 12.950 ;
      LAYER met1 ;
        RECT 7.000 12.600 8.050 12.950 ;
      LAYER met1 ;
        RECT 5.600 12.250 6.650 12.600 ;
      LAYER met1 ;
        RECT 6.650 12.250 8.050 12.600 ;
      LAYER met1 ;
        RECT 8.050 12.250 10.500 12.950 ;
      LAYER met1 ;
        RECT 10.500 12.250 11.550 12.950 ;
      LAYER met1 ;
        RECT 11.550 12.250 13.300 12.950 ;
      LAYER met1 ;
        RECT 13.300 12.250 17.150 12.950 ;
        RECT 0.000 11.900 17.150 12.250 ;
        RECT 0.000 10.850 1.400 11.900 ;
      LAYER met1 ;
        RECT 1.400 10.850 4.200 11.900 ;
      LAYER met1 ;
        RECT 4.200 11.550 5.600 11.900 ;
      LAYER met1 ;
        RECT 5.600 11.550 8.750 11.900 ;
      LAYER met1 ;
        RECT 4.200 10.850 5.250 11.550 ;
      LAYER met1 ;
        RECT 5.250 10.850 8.750 11.550 ;
      LAYER met1 ;
        RECT 8.750 10.850 9.450 11.900 ;
        RECT 0.000 10.500 1.750 10.850 ;
      LAYER met1 ;
        RECT 1.750 10.500 4.200 10.850 ;
      LAYER met1 ;
        RECT 4.200 10.500 4.900 10.850 ;
      LAYER met1 ;
        RECT 4.900 10.500 6.650 10.850 ;
      LAYER met1 ;
        RECT 6.650 10.500 7.700 10.850 ;
        RECT 0.000 7.350 2.100 10.500 ;
        RECT 0.000 6.300 0.350 7.350 ;
      LAYER met1 ;
        RECT 0.350 6.650 1.750 7.350 ;
      LAYER met1 ;
        RECT 1.750 6.650 2.100 7.350 ;
      LAYER met1 ;
        RECT 2.100 6.650 3.500 10.500 ;
      LAYER met1 ;
        RECT 3.500 9.100 4.900 10.500 ;
      LAYER met1 ;
        RECT 4.900 9.450 6.300 10.500 ;
      LAYER met1 ;
        RECT 6.300 9.800 7.700 10.500 ;
      LAYER met1 ;
        RECT 7.700 9.800 9.100 10.850 ;
      LAYER met1 ;
        RECT 9.100 9.800 9.450 10.850 ;
        RECT 6.300 9.450 9.450 9.800 ;
      LAYER met1 ;
        RECT 4.900 9.100 6.650 9.450 ;
      LAYER met1 ;
        RECT 6.650 9.100 7.700 9.450 ;
      LAYER met1 ;
        RECT 7.700 9.100 8.400 9.450 ;
      LAYER met1 ;
        RECT 8.400 9.100 9.450 9.450 ;
      LAYER met1 ;
        RECT 9.450 9.100 10.850 11.900 ;
      LAYER met1 ;
        RECT 10.850 11.200 12.250 11.900 ;
      LAYER met1 ;
        RECT 12.250 11.200 13.650 11.900 ;
      LAYER met1 ;
        RECT 10.850 10.150 11.900 11.200 ;
      LAYER met1 ;
        RECT 11.900 10.850 13.650 11.200 ;
      LAYER met1 ;
        RECT 13.650 10.850 17.150 11.900 ;
      LAYER met1 ;
        RECT 11.900 10.150 13.300 10.850 ;
      LAYER met1 ;
        RECT 10.850 9.100 11.200 10.150 ;
      LAYER met1 ;
        RECT 11.200 9.800 13.300 10.150 ;
      LAYER met1 ;
        RECT 13.300 9.800 17.150 10.850 ;
      LAYER met1 ;
        RECT 11.200 9.100 12.600 9.800 ;
      LAYER met1 ;
        RECT 3.500 8.400 5.250 9.100 ;
      LAYER met1 ;
        RECT 5.250 8.400 8.750 9.100 ;
      LAYER met1 ;
        RECT 8.750 8.400 9.450 9.100 ;
      LAYER met1 ;
        RECT 9.450 8.750 12.600 9.100 ;
      LAYER met1 ;
        RECT 12.600 8.750 17.150 9.800 ;
      LAYER met1 ;
        RECT 9.450 8.400 11.900 8.750 ;
      LAYER met1 ;
        RECT 11.900 8.400 17.150 8.750 ;
        RECT 3.500 8.050 5.600 8.400 ;
      LAYER met1 ;
        RECT 5.600 8.050 9.100 8.400 ;
      LAYER met1 ;
        RECT 3.500 7.350 7.700 8.050 ;
      LAYER met1 ;
        RECT 0.350 6.300 3.500 6.650 ;
      LAYER met1 ;
        RECT 3.500 6.300 4.900 7.350 ;
      LAYER met1 ;
        RECT 4.900 6.650 6.300 7.350 ;
      LAYER met1 ;
        RECT 6.300 6.650 7.700 7.350 ;
      LAYER met1 ;
        RECT 7.700 6.650 9.100 8.050 ;
        RECT 4.900 6.300 9.100 6.650 ;
      LAYER met1 ;
        RECT 9.100 6.300 9.450 8.400 ;
      LAYER met1 ;
        RECT 9.450 8.050 12.600 8.400 ;
      LAYER met1 ;
        RECT 0.000 5.600 0.700 6.300 ;
      LAYER met1 ;
        RECT 0.700 5.600 3.150 6.300 ;
      LAYER met1 ;
        RECT 3.150 5.600 5.250 6.300 ;
      LAYER met1 ;
        RECT 5.250 5.600 8.750 6.300 ;
      LAYER met1 ;
        RECT 0.000 5.250 1.050 5.600 ;
      LAYER met1 ;
        RECT 1.050 5.250 3.150 5.600 ;
      LAYER met1 ;
        RECT 3.150 5.250 5.600 5.600 ;
      LAYER met1 ;
        RECT 5.600 5.250 8.750 5.600 ;
      LAYER met1 ;
        RECT 8.750 5.250 9.450 6.300 ;
      LAYER met1 ;
        RECT 9.450 5.250 10.850 8.050 ;
      LAYER met1 ;
        RECT 10.850 7.000 11.200 8.050 ;
      LAYER met1 ;
        RECT 11.200 7.350 12.600 8.050 ;
      LAYER met1 ;
        RECT 12.600 7.350 17.150 8.400 ;
      LAYER met1 ;
        RECT 11.200 7.000 13.300 7.350 ;
      LAYER met1 ;
        RECT 10.850 6.300 11.900 7.000 ;
      LAYER met1 ;
        RECT 11.900 6.650 13.300 7.000 ;
      LAYER met1 ;
        RECT 13.300 6.650 17.150 7.350 ;
      LAYER met1 ;
        RECT 11.900 6.300 13.650 6.650 ;
      LAYER met1 ;
        RECT 10.850 5.250 12.250 6.300 ;
      LAYER met1 ;
        RECT 12.250 5.250 13.650 6.300 ;
      LAYER met1 ;
        RECT 13.650 5.250 17.150 6.650 ;
        RECT 0.000 4.900 17.150 5.250 ;
        RECT 0.000 3.850 1.400 4.900 ;
      LAYER met1 ;
        RECT 1.400 4.550 3.850 4.900 ;
      LAYER met1 ;
        RECT 3.850 4.550 4.550 4.900 ;
      LAYER met1 ;
        RECT 4.550 4.550 7.000 4.900 ;
      LAYER met1 ;
        RECT 7.000 4.550 8.750 4.900 ;
      LAYER met1 ;
        RECT 8.750 4.550 9.450 4.900 ;
        RECT 1.400 4.200 4.200 4.550 ;
      LAYER met1 ;
        RECT 4.200 4.200 4.550 4.550 ;
      LAYER met1 ;
        RECT 4.550 4.200 7.350 4.550 ;
      LAYER met1 ;
        RECT 7.350 4.200 8.400 4.550 ;
      LAYER met1 ;
        RECT 8.400 4.200 9.450 4.550 ;
      LAYER met1 ;
        RECT 9.450 4.200 11.550 4.900 ;
      LAYER met1 ;
        RECT 11.550 4.200 12.600 4.900 ;
      LAYER met1 ;
        RECT 12.600 4.200 17.150 4.900 ;
      LAYER met1 ;
        RECT 1.400 3.850 3.850 4.200 ;
      LAYER met1 ;
        RECT 3.850 3.850 4.550 4.200 ;
      LAYER met1 ;
        RECT 4.550 3.850 7.000 4.200 ;
      LAYER met1 ;
        RECT 7.000 3.850 8.050 4.200 ;
        RECT 0.000 0.350 2.100 3.850 ;
      LAYER met1 ;
        RECT 2.100 0.350 3.150 3.850 ;
      LAYER met1 ;
        RECT 3.150 0.350 5.250 3.850 ;
      LAYER met1 ;
        RECT 5.250 0.350 6.300 3.850 ;
      LAYER met1 ;
        RECT 6.300 3.500 8.050 3.850 ;
      LAYER met1 ;
        RECT 8.050 3.500 9.450 4.200 ;
      LAYER met1 ;
        RECT 9.450 3.500 11.200 4.200 ;
      LAYER met1 ;
        RECT 11.200 3.850 12.950 4.200 ;
      LAYER met1 ;
        RECT 12.950 3.850 17.150 4.200 ;
      LAYER met1 ;
        RECT 11.200 3.500 11.900 3.850 ;
      LAYER met1 ;
        RECT 6.300 1.400 8.400 3.500 ;
      LAYER met1 ;
        RECT 8.400 1.400 9.450 3.500 ;
      LAYER met1 ;
        RECT 9.450 1.750 10.850 3.500 ;
      LAYER met1 ;
        RECT 10.850 1.750 11.900 3.500 ;
      LAYER met1 ;
        RECT 9.450 1.400 11.200 1.750 ;
      LAYER met1 ;
        RECT 11.200 1.400 11.900 1.750 ;
      LAYER met1 ;
        RECT 11.900 1.400 12.250 3.850 ;
      LAYER met1 ;
        RECT 12.250 1.400 13.300 3.850 ;
      LAYER met1 ;
        RECT 13.300 1.400 17.150 3.850 ;
        RECT 6.300 0.350 8.050 1.400 ;
      LAYER met1 ;
        RECT 8.050 1.050 9.800 1.400 ;
      LAYER met1 ;
        RECT 9.800 1.050 11.200 1.400 ;
      LAYER met1 ;
        RECT 11.200 1.050 12.950 1.400 ;
        RECT 8.050 0.350 10.150 1.050 ;
      LAYER met1 ;
        RECT 10.150 0.350 11.550 1.050 ;
      LAYER met1 ;
        RECT 11.550 0.700 12.950 1.050 ;
      LAYER met1 ;
        RECT 12.950 0.700 17.150 1.400 ;
      LAYER met1 ;
        RECT 11.550 0.350 12.600 0.700 ;
      LAYER met1 ;
        RECT 12.600 0.350 17.150 0.700 ;
        RECT 0.000 0.000 17.150 0.350 ;
      LAYER met2 ;
        RECT 2.100 16.100 3.850 16.800 ;
        RECT 5.600 16.100 6.650 16.800 ;
        RECT 8.400 16.100 10.150 16.800 ;
        RECT 1.750 15.750 4.200 16.100 ;
        RECT 1.750 15.400 2.450 15.750 ;
        RECT 3.150 14.700 4.200 15.750 ;
        RECT 5.250 15.750 7.000 16.100 ;
        RECT 8.050 15.750 10.500 16.100 ;
        RECT 5.250 15.400 5.950 15.750 ;
        RECT 2.800 14.350 3.850 14.700 ;
        RECT 2.450 14.000 3.850 14.350 ;
        RECT 2.450 13.650 3.500 14.000 ;
        RECT 4.900 13.650 5.950 15.400 ;
        RECT 2.100 12.950 3.150 13.650 ;
        RECT 5.250 13.300 5.950 13.650 ;
        RECT 6.300 13.300 7.350 15.750 ;
        RECT 8.050 15.400 8.750 15.750 ;
        RECT 9.450 14.700 10.500 15.750 ;
        RECT 11.200 15.750 13.650 16.800 ;
        RECT 11.200 15.400 12.250 15.750 ;
        RECT 11.200 15.050 13.300 15.400 ;
        RECT 9.100 14.350 10.150 14.700 ;
        RECT 8.750 14.000 10.150 14.350 ;
        RECT 11.200 14.350 13.650 15.050 ;
        RECT 11.200 14.000 12.250 14.350 ;
        RECT 12.600 14.000 13.650 14.350 ;
        RECT 8.750 13.650 9.800 14.000 ;
        RECT 12.950 13.650 13.650 14.000 ;
        RECT 3.500 12.950 4.200 13.300 ;
        RECT 5.250 12.950 7.000 13.300 ;
        RECT 8.400 12.950 9.450 13.650 ;
        RECT 11.200 13.300 11.900 13.650 ;
        RECT 9.800 12.950 10.500 13.300 ;
        RECT 11.200 12.950 12.250 13.300 ;
        RECT 12.600 12.950 13.650 13.650 ;
        RECT 1.750 12.250 4.200 12.950 ;
        RECT 5.600 12.600 7.000 12.950 ;
        RECT 5.600 12.250 6.650 12.600 ;
        RECT 8.050 12.250 10.500 12.950 ;
        RECT 11.550 12.250 13.300 12.950 ;
        RECT 1.400 10.850 4.200 11.900 ;
        RECT 5.600 11.550 8.750 11.900 ;
        RECT 5.250 10.850 8.750 11.550 ;
        RECT 1.750 10.500 4.200 10.850 ;
        RECT 4.900 10.500 6.650 10.850 ;
        RECT 0.350 6.650 1.750 7.350 ;
        RECT 2.100 6.650 3.500 10.500 ;
        RECT 4.900 9.450 6.300 10.500 ;
        RECT 7.700 9.800 9.100 10.850 ;
        RECT 4.900 9.100 6.650 9.450 ;
        RECT 7.700 9.100 8.400 9.450 ;
        RECT 9.450 9.100 10.850 11.900 ;
        RECT 12.250 11.200 13.650 11.900 ;
        RECT 11.900 10.850 13.650 11.200 ;
        RECT 11.900 10.150 13.300 10.850 ;
        RECT 11.200 9.800 13.300 10.150 ;
        RECT 11.200 9.100 12.600 9.800 ;
        RECT 5.250 8.400 8.750 9.100 ;
        RECT 9.450 8.750 12.600 9.100 ;
        RECT 9.450 8.400 11.900 8.750 ;
        RECT 5.600 8.050 9.100 8.400 ;
        RECT 0.350 6.300 3.500 6.650 ;
        RECT 4.900 6.650 6.300 7.350 ;
        RECT 7.700 6.650 9.100 8.050 ;
        RECT 4.900 6.300 9.100 6.650 ;
        RECT 9.450 8.050 12.600 8.400 ;
        RECT 0.700 5.600 3.150 6.300 ;
        RECT 5.250 5.600 8.750 6.300 ;
        RECT 1.050 5.250 3.150 5.600 ;
        RECT 5.600 5.250 8.750 5.600 ;
        RECT 9.450 5.250 10.850 8.050 ;
        RECT 11.200 7.350 12.600 8.050 ;
        RECT 11.200 7.000 13.300 7.350 ;
        RECT 11.900 6.650 13.300 7.000 ;
        RECT 11.900 6.300 13.650 6.650 ;
        RECT 12.250 5.250 13.650 6.300 ;
        RECT 1.400 4.550 3.850 4.900 ;
        RECT 4.550 4.550 7.000 4.900 ;
        RECT 8.750 4.550 9.450 4.900 ;
        RECT 1.400 4.200 4.200 4.550 ;
        RECT 4.550 4.200 7.350 4.550 ;
        RECT 8.400 4.200 9.450 4.550 ;
        RECT 11.550 4.200 12.600 4.900 ;
        RECT 1.400 3.850 3.850 4.200 ;
        RECT 4.550 3.850 7.000 4.200 ;
        RECT 2.100 0.350 3.150 3.850 ;
        RECT 5.250 0.350 6.300 3.850 ;
        RECT 8.050 3.500 9.450 4.200 ;
        RECT 11.200 3.850 12.950 4.200 ;
        RECT 11.200 3.500 11.900 3.850 ;
        RECT 8.400 1.400 9.450 3.500 ;
        RECT 10.850 1.750 11.900 3.500 ;
        RECT 11.200 1.400 11.900 1.750 ;
        RECT 12.250 1.400 13.300 3.850 ;
        RECT 8.050 1.050 9.800 1.400 ;
        RECT 11.200 1.050 12.950 1.400 ;
        RECT 8.050 0.350 10.150 1.050 ;
        RECT 11.550 0.700 12.950 1.050 ;
        RECT 11.550 0.350 12.600 0.700 ;
  END
END my_logo
END LIBRARY

