magic
tech sky130A
magscale 1 2
timestamp 1738297850
<< viali >>
rect 7205 44489 7239 44523
rect 7665 44489 7699 44523
rect 7941 44489 7975 44523
rect 8769 44489 8803 44523
rect 9321 44489 9355 44523
rect 11713 44489 11747 44523
rect 12817 44489 12851 44523
rect 13093 44489 13127 44523
rect 26433 44421 26467 44455
rect 29009 44353 29043 44387
rect 8033 44285 8067 44319
rect 8585 44285 8619 44319
rect 9137 44285 9171 44319
rect 12357 44285 12391 44319
rect 12449 44285 12483 44319
rect 13737 44285 13771 44319
rect 13829 44285 13863 44319
rect 14013 44285 14047 44319
rect 14105 44285 14139 44319
rect 14565 44285 14599 44319
rect 15209 44285 15243 44319
rect 17049 44285 17083 44319
rect 19349 44285 19383 44319
rect 21649 44285 21683 44319
rect 24041 44285 24075 44319
rect 24409 44285 24443 44319
rect 24961 44285 24995 44319
rect 25513 44285 25547 44319
rect 25789 44285 25823 44319
rect 26065 44285 26099 44319
rect 27813 44285 27847 44319
rect 27905 44285 27939 44319
rect 28181 44285 28215 44319
rect 29285 44285 29319 44319
rect 27546 44217 27580 44251
rect 8125 44149 8159 44183
rect 12265 44149 12299 44183
rect 12541 44149 12575 44183
rect 13553 44149 13587 44183
rect 14473 44149 14507 44183
rect 15025 44149 15059 44183
rect 16957 44149 16991 44183
rect 19441 44149 19475 44183
rect 21833 44149 21867 44183
rect 23857 44149 23891 44183
rect 24593 44149 24627 44183
rect 25145 44149 25179 44183
rect 25697 44149 25731 44183
rect 25973 44149 26007 44183
rect 26249 44149 26283 44183
rect 28089 44149 28123 44183
rect 28365 44149 28399 44183
rect 6561 43945 6595 43979
rect 6929 43945 6963 43979
rect 9689 43945 9723 43979
rect 10701 43945 10735 43979
rect 13277 43945 13311 43979
rect 13553 43945 13587 43979
rect 18153 43945 18187 43979
rect 26433 43945 26467 43979
rect 27905 43945 27939 43979
rect 15945 43877 15979 43911
rect 22394 43877 22428 43911
rect 23213 43877 23247 43911
rect 25154 43877 25188 43911
rect 27546 43877 27580 43911
rect 6745 43809 6779 43843
rect 7113 43809 7147 43843
rect 8309 43809 8343 43843
rect 8576 43809 8610 43843
rect 10333 43809 10367 43843
rect 10517 43809 10551 43843
rect 12090 43809 12124 43843
rect 12357 43809 12391 43843
rect 12817 43809 12851 43843
rect 13369 43809 13403 43843
rect 14289 43809 14323 43843
rect 16313 43809 16347 43843
rect 16773 43809 16807 43843
rect 19257 43809 19291 43843
rect 23121 43809 23155 43843
rect 23305 43809 23339 43843
rect 23489 43809 23523 43843
rect 29018 43809 29052 43843
rect 29285 43809 29319 43843
rect 14197 43741 14231 43775
rect 14565 43741 14599 43775
rect 17049 43741 17083 43775
rect 19533 43741 19567 43775
rect 22661 43741 22695 43775
rect 25421 43741 25455 43775
rect 27813 43741 27847 43775
rect 16129 43673 16163 43707
rect 9781 43605 9815 43639
rect 10977 43605 11011 43639
rect 12725 43605 12759 43639
rect 20637 43605 20671 43639
rect 21281 43605 21315 43639
rect 22937 43605 22971 43639
rect 24041 43605 24075 43639
rect 8861 43401 8895 43435
rect 11621 43401 11655 43435
rect 13645 43401 13679 43435
rect 15301 43401 15335 43435
rect 13369 43333 13403 43367
rect 15117 43265 15151 43299
rect 18797 43265 18831 43299
rect 9229 43197 9263 43231
rect 9597 43197 9631 43231
rect 9689 43197 9723 43231
rect 9781 43197 9815 43231
rect 11437 43197 11471 43231
rect 11989 43197 12023 43231
rect 12256 43197 12290 43231
rect 13829 43197 13863 43231
rect 14105 43197 14139 43231
rect 14841 43197 14875 43231
rect 15025 43197 15059 43231
rect 15577 43197 15611 43231
rect 15669 43197 15703 43231
rect 15761 43197 15795 43231
rect 15945 43197 15979 43231
rect 16037 43197 16071 43231
rect 16313 43197 16347 43231
rect 16773 43197 16807 43231
rect 17049 43197 17083 43231
rect 17417 43197 17451 43231
rect 17693 43197 17727 43231
rect 17923 43197 17957 43231
rect 18281 43197 18315 43231
rect 18429 43197 18463 43231
rect 18705 43197 18739 43231
rect 19257 43197 19291 43231
rect 19625 43197 19659 43231
rect 19717 43197 19751 43231
rect 19993 43197 20027 43231
rect 20545 43197 20579 43231
rect 21281 43197 21315 43231
rect 21557 43197 21591 43231
rect 21741 43197 21775 43231
rect 24970 43197 25004 43231
rect 25237 43197 25271 43231
rect 26709 43197 26743 43231
rect 28181 43197 28215 43231
rect 9045 43129 9079 43163
rect 16129 43129 16163 43163
rect 16957 43129 16991 43163
rect 18061 43129 18095 43163
rect 18153 43129 18187 43163
rect 19349 43129 19383 43163
rect 19441 43129 19475 43163
rect 22008 43129 22042 43163
rect 23305 43129 23339 43163
rect 26442 43129 26476 43163
rect 27936 43129 27970 43163
rect 9873 43061 9907 43095
rect 14749 43061 14783 43095
rect 16497 43061 16531 43095
rect 16589 43061 16623 43095
rect 17233 43061 17267 43095
rect 17601 43061 17635 43095
rect 17785 43061 17819 43095
rect 19073 43061 19107 43095
rect 19809 43061 19843 43095
rect 20177 43061 20211 43095
rect 20361 43061 20395 43095
rect 21097 43061 21131 43095
rect 21465 43061 21499 43095
rect 23121 43061 23155 43095
rect 23581 43061 23615 43095
rect 23857 43061 23891 43095
rect 25329 43061 25363 43095
rect 26801 43061 26835 43095
rect 12173 42857 12207 42891
rect 13921 42857 13955 42891
rect 14105 42857 14139 42891
rect 15669 42857 15703 42891
rect 19717 42857 19751 42891
rect 22661 42857 22695 42891
rect 17509 42789 17543 42823
rect 9413 42721 9447 42755
rect 9680 42721 9714 42755
rect 12265 42721 12299 42755
rect 12541 42721 12575 42755
rect 12808 42721 12842 42755
rect 14013 42721 14047 42755
rect 16405 42721 16439 42755
rect 16498 42721 16532 42755
rect 16681 42721 16715 42755
rect 16773 42721 16807 42755
rect 16909 42721 16943 42755
rect 17417 42721 17451 42755
rect 17693 42721 17727 42755
rect 17969 42721 18003 42755
rect 19625 42721 19659 42755
rect 19993 42721 20027 42755
rect 20085 42721 20119 42755
rect 20177 42721 20211 42755
rect 20361 42721 20395 42755
rect 21281 42721 21315 42755
rect 21537 42721 21571 42755
rect 22937 42721 22971 42755
rect 23029 42721 23063 42755
rect 23213 42721 23247 42755
rect 23305 42721 23339 42755
rect 23581 42721 23615 42755
rect 23673 42721 23707 42755
rect 23857 42721 23891 42755
rect 23949 42721 23983 42755
rect 24225 42721 24259 42755
rect 24317 42721 24351 42755
rect 24501 42721 24535 42755
rect 24593 42721 24627 42755
rect 29653 42721 29687 42755
rect 11529 42653 11563 42687
rect 14289 42653 14323 42687
rect 14565 42653 14599 42687
rect 19349 42653 19383 42687
rect 23397 42653 23431 42687
rect 10793 42585 10827 42619
rect 10977 42517 11011 42551
rect 17049 42517 17083 42551
rect 17877 42517 17911 42551
rect 22753 42517 22787 42551
rect 24041 42517 24075 42551
rect 29561 42517 29595 42551
rect 13553 42313 13587 42347
rect 14749 42313 14783 42347
rect 15025 42313 15059 42347
rect 17141 42313 17175 42347
rect 17325 42313 17359 42347
rect 21005 42313 21039 42347
rect 23857 42313 23891 42347
rect 18429 42245 18463 42279
rect 19533 42245 19567 42279
rect 15393 42177 15427 42211
rect 21281 42177 21315 42211
rect 13737 42109 13771 42143
rect 14013 42109 14047 42143
rect 14197 42109 14231 42143
rect 14657 42109 14691 42143
rect 15209 42109 15243 42143
rect 15485 42109 15519 42143
rect 15577 42109 15611 42143
rect 15761 42109 15795 42143
rect 16313 42109 16347 42143
rect 16405 42109 16439 42143
rect 16497 42109 16531 42143
rect 16681 42109 16715 42143
rect 16773 42109 16807 42143
rect 16957 42109 16991 42143
rect 18337 42099 18371 42133
rect 18496 42109 18530 42143
rect 18705 42109 18739 42143
rect 18889 42109 18923 42143
rect 18981 42109 19015 42143
rect 19073 42109 19107 42143
rect 19441 42109 19475 42143
rect 19625 42109 19659 42143
rect 20085 42109 20119 42143
rect 20269 42109 20303 42143
rect 20361 42109 20395 42143
rect 20545 42109 20579 42143
rect 20637 42109 20671 42143
rect 20729 42109 20763 42143
rect 21557 42109 21591 42143
rect 22385 42109 22419 42143
rect 23029 42109 23063 42143
rect 23121 42109 23155 42143
rect 23305 42109 23339 42143
rect 23397 42109 23431 42143
rect 24041 42109 24075 42143
rect 24133 42109 24167 42143
rect 24409 42109 24443 42143
rect 26709 42109 26743 42143
rect 28181 42109 28215 42143
rect 29561 42109 29595 42143
rect 30389 42109 30423 42143
rect 16037 42041 16071 42075
rect 16865 42041 16899 42075
rect 17293 42041 17327 42075
rect 17509 42041 17543 42075
rect 19349 42041 19383 42075
rect 20177 42041 20211 42075
rect 24225 42041 24259 42075
rect 21097 41973 21131 42007
rect 22293 41973 22327 42007
rect 22845 41973 22879 42007
rect 26617 41973 26651 42007
rect 28089 41973 28123 42007
rect 29009 41973 29043 42007
rect 29745 41973 29779 42007
rect 9689 41769 9723 41803
rect 13829 41769 13863 41803
rect 18061 41769 18095 41803
rect 29285 41769 29319 41803
rect 30757 41769 30791 41803
rect 9965 41633 9999 41667
rect 10057 41633 10091 41667
rect 10149 41633 10183 41667
rect 10333 41633 10367 41667
rect 13737 41633 13771 41667
rect 13921 41633 13955 41667
rect 17877 41633 17911 41667
rect 21281 41633 21315 41667
rect 21537 41633 21571 41667
rect 22753 41633 22787 41667
rect 23213 41633 23247 41667
rect 23949 41633 23983 41667
rect 26433 41633 26467 41667
rect 26700 41633 26734 41667
rect 27905 41633 27939 41667
rect 28172 41633 28206 41667
rect 29377 41633 29411 41667
rect 29633 41633 29667 41667
rect 13001 41565 13035 41599
rect 22661 41497 22695 41531
rect 22937 41497 22971 41531
rect 12449 41429 12483 41463
rect 23489 41429 23523 41463
rect 23765 41429 23799 41463
rect 27813 41429 27847 41463
rect 10609 41225 10643 41259
rect 15577 41225 15611 41259
rect 17969 41225 18003 41259
rect 18153 41225 18187 41259
rect 19533 41225 19567 41259
rect 20821 41225 20855 41259
rect 22845 41225 22879 41259
rect 26801 41225 26835 41259
rect 28181 41225 28215 41259
rect 28825 41225 28859 41259
rect 26249 41157 26283 41191
rect 9873 41089 9907 41123
rect 26617 41089 26651 41123
rect 27721 41089 27755 41123
rect 28273 41089 28307 41123
rect 29009 41089 29043 41123
rect 8585 41021 8619 41055
rect 8861 41021 8895 41055
rect 8953 41021 8987 41055
rect 9137 41021 9171 41055
rect 9229 41021 9263 41055
rect 10057 41021 10091 41055
rect 10149 41021 10183 41055
rect 10333 41021 10367 41055
rect 10425 41021 10459 41055
rect 11069 41021 11103 41055
rect 11161 41021 11195 41055
rect 11345 41021 11379 41055
rect 14381 41021 14415 41055
rect 15117 41021 15151 41055
rect 15209 41021 15243 41055
rect 15301 41021 15335 41055
rect 15485 41021 15519 41055
rect 15761 41021 15795 41055
rect 15853 41021 15887 41055
rect 16037 41021 16071 41055
rect 16129 41021 16163 41055
rect 16589 41021 16623 41055
rect 16773 41021 16807 41055
rect 17325 41021 17359 41055
rect 17693 41021 17727 41055
rect 18153 41021 18187 41055
rect 18521 41021 18555 41055
rect 19441 41021 19475 41055
rect 19625 41021 19659 41055
rect 19809 41021 19843 41055
rect 19993 41021 20027 41055
rect 20177 41021 20211 41055
rect 20361 41021 20395 41055
rect 20453 41021 20487 41055
rect 20545 41021 20579 41055
rect 22201 41021 22235 41055
rect 22753 41021 22787 41055
rect 23949 41021 23983 41055
rect 24216 41021 24250 41055
rect 26065 41021 26099 41055
rect 26525 41021 26559 41055
rect 26893 41021 26927 41055
rect 27169 41021 27203 41055
rect 27905 41021 27939 41055
rect 27997 41021 28031 41055
rect 28457 41021 28491 41055
rect 28549 41021 28583 41055
rect 28641 41021 28675 41055
rect 28825 41021 28859 41055
rect 29193 41021 29227 41055
rect 29285 41021 29319 41055
rect 30849 41021 30883 41055
rect 11612 40953 11646 40987
rect 12817 40953 12851 40987
rect 13001 40953 13035 40987
rect 16221 40953 16255 40987
rect 16405 40953 16439 40987
rect 17509 40953 17543 40987
rect 17601 40953 17635 40987
rect 23397 40953 23431 40987
rect 26249 40953 26283 40987
rect 28181 40953 28215 40987
rect 28273 40953 28307 40987
rect 29009 40953 29043 40987
rect 30604 40953 30638 40987
rect 8493 40885 8527 40919
rect 8677 40885 8711 40919
rect 9321 40885 9355 40919
rect 12725 40885 12759 40919
rect 13185 40885 13219 40919
rect 14289 40885 14323 40919
rect 14841 40885 14875 40919
rect 16681 40885 16715 40919
rect 17877 40885 17911 40919
rect 19993 40885 20027 40919
rect 22109 40885 22143 40919
rect 23305 40885 23339 40919
rect 25329 40885 25363 40919
rect 25513 40885 25547 40919
rect 26433 40885 26467 40919
rect 26617 40885 26651 40919
rect 29469 40885 29503 40919
rect 10793 40681 10827 40715
rect 10977 40681 11011 40715
rect 11805 40681 11839 40715
rect 15485 40681 15519 40715
rect 23305 40681 23339 40715
rect 24133 40681 24167 40715
rect 24869 40681 24903 40715
rect 25973 40681 26007 40715
rect 30849 40681 30883 40715
rect 31125 40681 31159 40715
rect 18061 40613 18095 40647
rect 19073 40613 19107 40647
rect 21465 40613 21499 40647
rect 30665 40613 30699 40647
rect 8125 40545 8159 40579
rect 8392 40545 8426 40579
rect 9689 40545 9723 40579
rect 9873 40545 9907 40579
rect 10057 40545 10091 40579
rect 10149 40545 10183 40579
rect 10333 40545 10367 40579
rect 10425 40545 10459 40579
rect 10517 40545 10551 40579
rect 11345 40545 11379 40579
rect 12081 40545 12115 40579
rect 12173 40545 12207 40579
rect 12265 40545 12299 40579
rect 12443 40545 12477 40579
rect 12909 40545 12943 40579
rect 13001 40545 13035 40579
rect 13093 40545 13127 40579
rect 13277 40545 13311 40579
rect 14105 40545 14139 40579
rect 14381 40545 14415 40579
rect 16497 40545 16531 40579
rect 16773 40545 16807 40579
rect 16957 40545 16991 40579
rect 17509 40545 17543 40579
rect 17693 40545 17727 40579
rect 18889 40545 18923 40579
rect 19165 40545 19199 40579
rect 21281 40545 21315 40579
rect 21925 40545 21959 40579
rect 22192 40545 22226 40579
rect 23489 40545 23523 40579
rect 24225 40545 24259 40579
rect 25145 40545 25179 40579
rect 25881 40545 25915 40579
rect 26065 40545 26099 40579
rect 26617 40545 26651 40579
rect 28365 40545 28399 40579
rect 28457 40545 28491 40579
rect 29653 40545 29687 40579
rect 30297 40545 30331 40579
rect 30389 40545 30423 40579
rect 30757 40545 30791 40579
rect 30941 40545 30975 40579
rect 31033 40545 31067 40579
rect 11437 40477 11471 40511
rect 11529 40477 11563 40511
rect 16589 40477 16623 40511
rect 17049 40477 17083 40511
rect 17233 40477 17267 40511
rect 17325 40477 17359 40511
rect 17417 40477 17451 40511
rect 17877 40477 17911 40511
rect 24869 40477 24903 40511
rect 25053 40477 25087 40511
rect 26433 40477 26467 40511
rect 26801 40477 26835 40511
rect 30665 40477 30699 40511
rect 16681 40409 16715 40443
rect 17991 40409 18025 40443
rect 9505 40341 9539 40375
rect 12633 40341 12667 40375
rect 16313 40341 16347 40375
rect 17785 40341 17819 40375
rect 18705 40341 18739 40375
rect 21649 40341 21683 40375
rect 23581 40341 23615 40375
rect 28641 40341 28675 40375
rect 30481 40341 30515 40375
rect 8861 40137 8895 40171
rect 9689 40137 9723 40171
rect 11161 40137 11195 40171
rect 15393 40137 15427 40171
rect 16129 40137 16163 40171
rect 17233 40137 17267 40171
rect 25145 40137 25179 40171
rect 27445 40137 27479 40171
rect 28641 40137 28675 40171
rect 22937 40069 22971 40103
rect 26157 40069 26191 40103
rect 10241 40001 10275 40035
rect 11713 40001 11747 40035
rect 11805 40001 11839 40035
rect 13093 40001 13127 40035
rect 13185 40001 13219 40035
rect 20085 40001 20119 40035
rect 21925 40001 21959 40035
rect 27997 40001 28031 40035
rect 28181 40001 28215 40035
rect 30941 40001 30975 40035
rect 9137 39933 9171 39967
rect 9229 39933 9263 39967
rect 9321 39933 9355 39967
rect 9505 39933 9539 39967
rect 10057 39933 10091 39967
rect 10609 39933 10643 39967
rect 10701 39933 10735 39967
rect 10885 39933 10919 39967
rect 10977 39933 11011 39967
rect 12265 39933 12299 39967
rect 13553 39933 13587 39967
rect 15577 39933 15611 39967
rect 15669 39933 15703 39967
rect 15853 39933 15887 39967
rect 15945 39933 15979 39967
rect 16405 39933 16439 39967
rect 16497 39933 16531 39967
rect 16589 39933 16623 39967
rect 16773 39933 16807 39967
rect 17141 39933 17175 39967
rect 17325 39933 17359 39967
rect 18337 39933 18371 39967
rect 18429 39933 18463 39967
rect 18705 39933 18739 39967
rect 18981 39933 19015 39967
rect 20453 39933 20487 39967
rect 20637 39933 20671 39967
rect 21281 39933 21315 39967
rect 21465 39933 21499 39967
rect 21557 39933 21591 39967
rect 21649 39933 21683 39967
rect 22201 39933 22235 39967
rect 22385 39933 22419 39967
rect 23305 39933 23339 39967
rect 23489 39933 23523 39967
rect 23673 39933 23707 39967
rect 24317 39933 24351 39967
rect 25973 39933 26007 39967
rect 26341 39933 26375 39967
rect 27077 39933 27111 39967
rect 28089 39933 28123 39967
rect 28273 39933 28307 39967
rect 30389 39933 30423 39967
rect 30757 39933 30791 39967
rect 31033 39933 31067 39967
rect 8585 39865 8619 39899
rect 8769 39865 8803 39899
rect 12449 39865 12483 39899
rect 13798 39865 13832 39899
rect 22661 39865 22695 39899
rect 25113 39865 25147 39899
rect 25329 39865 25363 39899
rect 27445 39865 27479 39899
rect 28825 39865 28859 39899
rect 8401 39797 8435 39831
rect 10149 39797 10183 39831
rect 11253 39797 11287 39831
rect 11621 39797 11655 39831
rect 12081 39797 12115 39831
rect 12633 39797 12667 39831
rect 13001 39797 13035 39831
rect 14933 39797 14967 39831
rect 20545 39797 20579 39831
rect 22109 39797 22143 39831
rect 22477 39797 22511 39831
rect 23121 39797 23155 39831
rect 24409 39797 24443 39831
rect 24961 39797 24995 39831
rect 25421 39797 25455 39831
rect 27629 39797 27663 39831
rect 27813 39797 27847 39831
rect 28457 39797 28491 39831
rect 28625 39797 28659 39831
rect 29837 39797 29871 39831
rect 30573 39797 30607 39831
rect 31125 39797 31159 39831
rect 10241 39593 10275 39627
rect 11253 39593 11287 39627
rect 13461 39593 13495 39627
rect 13737 39593 13771 39627
rect 15301 39593 15335 39627
rect 15669 39593 15703 39627
rect 19165 39593 19199 39627
rect 22661 39593 22695 39627
rect 25605 39593 25639 39627
rect 26065 39593 26099 39627
rect 26433 39593 26467 39627
rect 9597 39457 9631 39491
rect 9781 39457 9815 39491
rect 9873 39457 9907 39491
rect 9965 39457 9999 39491
rect 11529 39457 11563 39491
rect 11621 39457 11655 39491
rect 11713 39457 11747 39491
rect 11897 39457 11931 39491
rect 12357 39457 12391 39491
rect 12449 39457 12483 39491
rect 12633 39457 12667 39491
rect 12725 39457 12759 39491
rect 12817 39457 12851 39491
rect 13001 39457 13035 39491
rect 13093 39457 13127 39491
rect 13185 39457 13219 39491
rect 13829 39457 13863 39491
rect 15485 39457 15519 39491
rect 15761 39457 15795 39491
rect 18521 39457 18555 39491
rect 18705 39457 18739 39491
rect 18797 39457 18831 39491
rect 18889 39457 18923 39491
rect 19257 39457 19291 39491
rect 19441 39457 19475 39491
rect 19809 39457 19843 39491
rect 20177 39457 20211 39491
rect 20361 39457 20395 39491
rect 20453 39457 20487 39491
rect 20637 39457 20671 39491
rect 20729 39457 20763 39491
rect 20821 39457 20855 39491
rect 21281 39457 21315 39491
rect 21537 39457 21571 39491
rect 22753 39457 22787 39491
rect 23020 39457 23054 39491
rect 24225 39457 24259 39491
rect 24492 39457 24526 39491
rect 25697 39457 25731 39491
rect 27353 39457 27387 39491
rect 28411 39457 28445 39491
rect 29285 39457 29319 39491
rect 29837 39457 29871 39491
rect 31042 39457 31076 39491
rect 31309 39457 31343 39491
rect 14013 39389 14047 39423
rect 14565 39389 14599 39423
rect 19349 39389 19383 39423
rect 20269 39389 20303 39423
rect 21097 39389 21131 39423
rect 26617 39389 26651 39423
rect 26709 39389 26743 39423
rect 26801 39389 26835 39423
rect 26893 39389 26927 39423
rect 28273 39389 28307 39423
rect 28549 39389 28583 39423
rect 29469 39389 29503 39423
rect 29561 39389 29595 39423
rect 28825 39321 28859 39355
rect 29929 39321 29963 39355
rect 12173 39253 12207 39287
rect 19901 39253 19935 39287
rect 24133 39253 24167 39287
rect 26065 39253 26099 39287
rect 26249 39253 26283 39287
rect 27261 39253 27295 39287
rect 27629 39253 27663 39287
rect 29653 39253 29687 39287
rect 29745 39253 29779 39287
rect 24685 39049 24719 39083
rect 25053 39049 25087 39083
rect 27169 39049 27203 39083
rect 29561 39049 29595 39083
rect 30205 39049 30239 39083
rect 16405 38981 16439 39015
rect 17417 38981 17451 39015
rect 29745 38981 29779 39015
rect 10241 38913 10275 38947
rect 16957 38913 16991 38947
rect 25145 38913 25179 38947
rect 25881 38913 25915 38947
rect 26157 38913 26191 38947
rect 26295 38913 26329 38947
rect 8585 38845 8619 38879
rect 9045 38845 9079 38879
rect 9137 38845 9171 38879
rect 9321 38845 9355 38879
rect 9413 38845 9447 38879
rect 12357 38845 12391 38879
rect 15577 38845 15611 38879
rect 15761 38845 15795 38879
rect 16313 38845 16347 38879
rect 17233 38845 17267 38879
rect 19993 38845 20027 38879
rect 24869 38845 24903 38879
rect 25237 38845 25271 38879
rect 25421 38845 25455 38879
rect 26433 38845 26467 38879
rect 28282 38845 28316 38879
rect 28549 38845 28583 38879
rect 28733 38845 28767 38879
rect 28825 38845 28859 38879
rect 30205 38845 30239 38879
rect 30389 38845 30423 38879
rect 9597 38777 9631 38811
rect 12173 38777 12207 38811
rect 20453 38777 20487 38811
rect 29377 38777 29411 38811
rect 8493 38709 8527 38743
rect 9689 38709 9723 38743
rect 12541 38709 12575 38743
rect 15945 38709 15979 38743
rect 16221 38709 16255 38743
rect 16773 38709 16807 38743
rect 16865 38709 16899 38743
rect 19901 38709 19935 38743
rect 20177 38709 20211 38743
rect 27077 38709 27111 38743
rect 29582 38709 29616 38743
rect 9505 38505 9539 38539
rect 14365 38505 14399 38539
rect 14657 38505 14691 38539
rect 15025 38505 15059 38539
rect 15301 38505 15335 38539
rect 17509 38505 17543 38539
rect 23581 38505 23615 38539
rect 28457 38505 28491 38539
rect 13093 38437 13127 38471
rect 14565 38437 14599 38471
rect 23489 38437 23523 38471
rect 27344 38437 27378 38471
rect 8125 38369 8159 38403
rect 8392 38369 8426 38403
rect 9873 38369 9907 38403
rect 9965 38369 9999 38403
rect 10057 38369 10091 38403
rect 10241 38369 10275 38403
rect 11437 38369 11471 38403
rect 11529 38369 11563 38403
rect 11621 38369 11655 38403
rect 11805 38369 11839 38403
rect 12449 38369 12483 38403
rect 13001 38369 13035 38403
rect 13737 38369 13771 38403
rect 13829 38369 13863 38403
rect 13921 38369 13955 38403
rect 14105 38369 14139 38403
rect 14841 38369 14875 38403
rect 15117 38369 15151 38403
rect 15485 38369 15519 38403
rect 16129 38369 16163 38403
rect 17877 38369 17911 38403
rect 18061 38369 18095 38403
rect 18797 38369 18831 38403
rect 19165 38369 19199 38403
rect 19349 38369 19383 38403
rect 19717 38369 19751 38403
rect 19984 38369 20018 38403
rect 22477 38369 22511 38403
rect 22661 38369 22695 38403
rect 23765 38369 23799 38403
rect 27077 38369 27111 38403
rect 29377 38369 29411 38403
rect 9597 38301 9631 38335
rect 11897 38301 11931 38335
rect 13277 38301 13311 38335
rect 15761 38301 15795 38335
rect 16405 38301 16439 38335
rect 18705 38301 18739 38335
rect 18889 38301 18923 38335
rect 18981 38301 19015 38335
rect 23949 38301 23983 38335
rect 12633 38233 12667 38267
rect 18521 38233 18555 38267
rect 19257 38233 19291 38267
rect 11161 38165 11195 38199
rect 13461 38165 13495 38199
rect 14197 38165 14231 38199
rect 14381 38165 14415 38199
rect 15669 38165 15703 38199
rect 17969 38165 18003 38199
rect 21097 38165 21131 38199
rect 22385 38165 22419 38199
rect 29285 38165 29319 38199
rect 9689 37961 9723 37995
rect 12541 37961 12575 37995
rect 13185 37961 13219 37995
rect 15209 37961 15243 37995
rect 15945 37961 15979 37995
rect 17233 37961 17267 37995
rect 18429 37961 18463 37995
rect 19809 37961 19843 37995
rect 23581 37961 23615 37995
rect 10149 37825 10183 37859
rect 10333 37825 10367 37859
rect 13645 37825 13679 37859
rect 13829 37825 13863 37859
rect 17877 37825 17911 37859
rect 19349 37825 19383 37859
rect 21925 37825 21959 37859
rect 22201 37825 22235 37859
rect 29101 37825 29135 37859
rect 10057 37757 10091 37791
rect 10885 37757 10919 37791
rect 10977 37757 11011 37791
rect 11161 37757 11195 37791
rect 11417 37757 11451 37791
rect 12633 37757 12667 37791
rect 12725 37757 12759 37791
rect 12909 37757 12943 37791
rect 13001 37757 13035 37791
rect 13737 37757 13771 37791
rect 15301 37757 15335 37791
rect 15485 37757 15519 37791
rect 15577 37757 15611 37791
rect 15669 37757 15703 37791
rect 16957 37757 16991 37791
rect 18245 37757 18279 37791
rect 18981 37757 19015 37791
rect 19533 37757 19567 37791
rect 20085 37757 20119 37791
rect 20177 37757 20211 37791
rect 20269 37757 20303 37791
rect 20453 37757 20487 37791
rect 20913 37757 20947 37791
rect 22017 37757 22051 37791
rect 24961 37757 24995 37791
rect 29368 37757 29402 37791
rect 30665 37757 30699 37791
rect 9413 37689 9447 37723
rect 9597 37689 9631 37723
rect 14096 37689 14130 37723
rect 17693 37689 17727 37723
rect 18797 37689 18831 37723
rect 18889 37689 18923 37723
rect 21649 37689 21683 37723
rect 22468 37689 22502 37723
rect 9229 37621 9263 37655
rect 17601 37621 17635 37655
rect 20637 37621 20671 37655
rect 21557 37621 21591 37655
rect 30481 37621 30515 37655
rect 31309 37621 31343 37655
rect 8861 37417 8895 37451
rect 14105 37417 14139 37451
rect 15945 37417 15979 37451
rect 20361 37417 20395 37451
rect 20453 37417 20487 37451
rect 22661 37417 22695 37451
rect 23397 37417 23431 37451
rect 30389 37417 30423 37451
rect 14289 37349 14323 37383
rect 16129 37349 16163 37383
rect 19165 37349 19199 37383
rect 24271 37349 24305 37383
rect 24501 37349 24535 37383
rect 25605 37349 25639 37383
rect 27629 37349 27663 37383
rect 30113 37349 30147 37383
rect 30757 37349 30791 37383
rect 9137 37281 9171 37315
rect 9229 37281 9263 37315
rect 9321 37281 9355 37315
rect 9505 37281 9539 37315
rect 10149 37281 10183 37315
rect 10333 37281 10367 37315
rect 10517 37281 10551 37315
rect 13553 37281 13587 37315
rect 15117 37281 15151 37315
rect 15761 37281 15795 37315
rect 16957 37281 16991 37315
rect 18245 37281 18279 37315
rect 19625 37281 19659 37315
rect 19717 37281 19751 37315
rect 19993 37281 20027 37315
rect 20177 37281 20211 37315
rect 20729 37281 20763 37315
rect 20821 37281 20855 37315
rect 20913 37281 20947 37315
rect 21097 37281 21131 37315
rect 21281 37281 21315 37315
rect 21537 37281 21571 37315
rect 22753 37281 22787 37315
rect 23581 37281 23615 37315
rect 24409 37281 24443 37315
rect 24593 37281 24627 37315
rect 24869 37281 24903 37315
rect 26157 37281 26191 37315
rect 26801 37281 26835 37315
rect 26893 37281 26927 37315
rect 28984 37281 29018 37315
rect 29101 37281 29135 37315
rect 30297 37281 30331 37315
rect 30481 37281 30515 37315
rect 31033 37281 31067 37315
rect 31125 37281 31159 37315
rect 31309 37281 31343 37315
rect 13829 37213 13863 37247
rect 15485 37213 15519 37247
rect 18337 37213 18371 37247
rect 23765 37213 23799 37247
rect 24133 37213 24167 37247
rect 26433 37213 26467 37247
rect 28825 37213 28859 37247
rect 29837 37213 29871 37247
rect 30021 37213 30055 37247
rect 30757 37213 30791 37247
rect 19165 37145 19199 37179
rect 27169 37145 27203 37179
rect 27353 37145 27387 37179
rect 29377 37145 29411 37179
rect 30665 37145 30699 37179
rect 31125 37145 31159 37179
rect 9597 37077 9631 37111
rect 10701 37077 10735 37111
rect 13737 37077 13771 37111
rect 15577 37077 15611 37111
rect 18429 37077 18463 37111
rect 18613 37077 18647 37111
rect 19901 37077 19935 37111
rect 24777 37077 24811 37111
rect 26065 37077 26099 37111
rect 27077 37077 27111 37111
rect 28181 37077 28215 37111
rect 30941 37077 30975 37111
rect 9781 36873 9815 36907
rect 15117 36873 15151 36907
rect 16221 36873 16255 36907
rect 17877 36873 17911 36907
rect 18981 36873 19015 36907
rect 21005 36873 21039 36907
rect 23673 36873 23707 36907
rect 27261 36873 27295 36907
rect 29653 36873 29687 36907
rect 13093 36805 13127 36839
rect 13829 36805 13863 36839
rect 21925 36805 21959 36839
rect 10333 36737 10367 36771
rect 13737 36737 13771 36771
rect 14565 36737 14599 36771
rect 16405 36737 16439 36771
rect 18041 36737 18075 36771
rect 23949 36737 23983 36771
rect 25881 36737 25915 36771
rect 27813 36737 27847 36771
rect 27905 36737 27939 36771
rect 8033 36669 8067 36703
rect 8125 36669 8159 36703
rect 8401 36669 8435 36703
rect 10517 36669 10551 36703
rect 11161 36669 11195 36703
rect 11253 36669 11287 36703
rect 11437 36669 11471 36703
rect 11529 36669 11563 36703
rect 14013 36669 14047 36703
rect 14749 36669 14783 36703
rect 15025 36669 15059 36703
rect 15117 36669 15151 36703
rect 15301 36669 15335 36703
rect 16129 36669 16163 36703
rect 16497 36669 16531 36703
rect 18153 36669 18187 36703
rect 18889 36669 18923 36703
rect 19257 36669 19291 36703
rect 19349 36669 19383 36703
rect 21097 36669 21131 36703
rect 21741 36669 21775 36703
rect 22109 36669 22143 36703
rect 23029 36669 23063 36703
rect 23305 36669 23339 36703
rect 23489 36669 23523 36703
rect 24133 36669 24167 36703
rect 24409 36669 24443 36703
rect 29193 36669 29227 36703
rect 29285 36669 29319 36703
rect 29929 36669 29963 36703
rect 8668 36601 8702 36635
rect 10425 36601 10459 36635
rect 13369 36601 13403 36635
rect 14381 36601 14415 36635
rect 18429 36601 18463 36635
rect 18521 36601 18555 36635
rect 20361 36601 20395 36635
rect 20545 36601 20579 36635
rect 20637 36601 20671 36635
rect 20821 36601 20855 36635
rect 23187 36601 23221 36635
rect 23397 36601 23431 36635
rect 24317 36601 24351 36635
rect 24654 36601 24688 36635
rect 26126 36601 26160 36635
rect 29469 36601 29503 36635
rect 30174 36601 30208 36635
rect 10885 36533 10919 36567
rect 10977 36533 11011 36567
rect 12909 36533 12943 36567
rect 18705 36533 18739 36567
rect 21281 36533 21315 36567
rect 21557 36533 21591 36567
rect 25789 36533 25823 36567
rect 27353 36533 27387 36567
rect 27721 36533 27755 36567
rect 29669 36533 29703 36567
rect 29837 36533 29871 36567
rect 31309 36533 31343 36567
rect 9045 36329 9079 36363
rect 10057 36329 10091 36363
rect 13185 36329 13219 36363
rect 14565 36329 14599 36363
rect 16221 36329 16255 36363
rect 23857 36329 23891 36363
rect 25329 36329 25363 36363
rect 30021 36329 30055 36363
rect 31033 36329 31067 36363
rect 16773 36261 16807 36295
rect 19533 36261 19567 36295
rect 19901 36261 19935 36295
rect 23371 36261 23405 36295
rect 24685 36261 24719 36295
rect 25145 36261 25179 36295
rect 30205 36261 30239 36295
rect 30665 36261 30699 36295
rect 9321 36193 9355 36227
rect 9413 36193 9447 36227
rect 9505 36193 9539 36227
rect 9689 36193 9723 36227
rect 10333 36193 10367 36227
rect 10425 36193 10459 36227
rect 10517 36193 10551 36227
rect 10701 36193 10735 36227
rect 11989 36193 12023 36227
rect 12081 36193 12115 36227
rect 12265 36193 12299 36227
rect 12357 36193 12391 36227
rect 12909 36193 12943 36227
rect 13369 36193 13403 36227
rect 13921 36193 13955 36227
rect 14381 36193 14415 36227
rect 14657 36193 14691 36227
rect 16129 36193 16163 36227
rect 16313 36193 16347 36227
rect 16589 36193 16623 36227
rect 16865 36193 16899 36227
rect 17969 36193 18003 36227
rect 18429 36193 18463 36227
rect 19717 36193 19751 36227
rect 19993 36193 20027 36227
rect 20177 36193 20211 36227
rect 20269 36193 20303 36227
rect 20361 36193 20395 36227
rect 21557 36193 21591 36227
rect 22109 36193 22143 36227
rect 22569 36193 22603 36227
rect 23489 36193 23523 36227
rect 23581 36193 23615 36227
rect 23673 36193 23707 36227
rect 24179 36193 24213 36227
rect 24317 36193 24351 36227
rect 24409 36193 24443 36227
rect 24501 36193 24535 36227
rect 24777 36193 24811 36227
rect 24961 36193 24995 36227
rect 25421 36193 25455 36227
rect 25881 36193 25915 36227
rect 25973 36193 26007 36227
rect 26249 36193 26283 36227
rect 26433 36193 26467 36227
rect 26616 36193 26650 36227
rect 26709 36193 26743 36227
rect 26801 36193 26835 36227
rect 26985 36193 27019 36227
rect 30573 36193 30607 36227
rect 30849 36193 30883 36227
rect 31125 36193 31159 36227
rect 13553 36125 13587 36159
rect 14105 36125 14139 36159
rect 18245 36125 18279 36159
rect 23213 36125 23247 36159
rect 24041 36125 24075 36159
rect 13645 36057 13679 36091
rect 22293 36057 22327 36091
rect 26157 36057 26191 36091
rect 11805 35989 11839 36023
rect 12633 35989 12667 36023
rect 14197 35989 14231 36023
rect 16405 35989 16439 36023
rect 17049 35989 17083 36023
rect 18429 35989 18463 36023
rect 18613 35989 18647 36023
rect 20637 35989 20671 36023
rect 21373 35989 21407 36023
rect 22017 35989 22051 36023
rect 25697 35989 25731 36023
rect 27077 35989 27111 36023
rect 30205 35989 30239 36023
rect 12725 35785 12759 35819
rect 21741 35785 21775 35819
rect 23213 35785 23247 35819
rect 24041 35785 24075 35819
rect 28365 35785 28399 35819
rect 16313 35649 16347 35683
rect 21833 35649 21867 35683
rect 9505 35581 9539 35615
rect 9689 35581 9723 35615
rect 9781 35581 9815 35615
rect 9873 35581 9907 35615
rect 10977 35581 11011 35615
rect 11069 35581 11103 35615
rect 11253 35581 11287 35615
rect 13001 35581 13035 35615
rect 13093 35581 13127 35615
rect 13185 35581 13219 35615
rect 13369 35581 13403 35615
rect 13921 35581 13955 35615
rect 15209 35581 15243 35615
rect 15393 35581 15427 35615
rect 15485 35581 15519 35615
rect 15577 35581 15611 35615
rect 15945 35581 15979 35615
rect 16129 35581 16163 35615
rect 16221 35581 16255 35615
rect 16497 35581 16531 35615
rect 16773 35581 16807 35615
rect 19073 35581 19107 35615
rect 20085 35581 20119 35615
rect 20177 35581 20211 35615
rect 20361 35581 20395 35615
rect 20628 35581 20662 35615
rect 23857 35581 23891 35615
rect 24041 35581 24075 35615
rect 27813 35581 27847 35615
rect 28089 35581 28123 35615
rect 11520 35513 11554 35547
rect 13553 35513 13587 35547
rect 13737 35513 13771 35547
rect 15853 35513 15887 35547
rect 16681 35513 16715 35547
rect 17018 35513 17052 35547
rect 22100 35513 22134 35547
rect 28273 35513 28307 35547
rect 10149 35445 10183 35479
rect 12633 35445 12667 35479
rect 18153 35445 18187 35479
rect 18981 35445 19015 35479
rect 27629 35445 27663 35479
rect 27997 35445 28031 35479
rect 9965 35241 9999 35275
rect 11437 35241 11471 35275
rect 12173 35241 12207 35275
rect 16589 35241 16623 35275
rect 16957 35241 16991 35275
rect 19073 35241 19107 35275
rect 22201 35241 22235 35275
rect 22477 35241 22511 35275
rect 22845 35241 22879 35275
rect 25329 35241 25363 35275
rect 26985 35241 27019 35275
rect 27277 35241 27311 35275
rect 27537 35241 27571 35275
rect 30021 35241 30055 35275
rect 14105 35173 14139 35207
rect 18429 35173 18463 35207
rect 21833 35173 21867 35207
rect 22049 35173 22083 35207
rect 26709 35173 26743 35207
rect 26893 35173 26927 35207
rect 27077 35173 27111 35207
rect 29837 35173 29871 35207
rect 30757 35173 30791 35207
rect 30849 35173 30883 35207
rect 11713 35105 11747 35139
rect 11805 35105 11839 35139
rect 11897 35105 11931 35139
rect 12081 35105 12115 35139
rect 12541 35105 12575 35139
rect 13277 35105 13311 35139
rect 13369 35105 13403 35139
rect 13553 35105 13587 35139
rect 13645 35105 13679 35139
rect 13737 35105 13771 35139
rect 14289 35105 14323 35139
rect 14381 35105 14415 35139
rect 14565 35105 14599 35139
rect 14657 35105 14691 35139
rect 14749 35105 14783 35139
rect 16129 35105 16163 35139
rect 16221 35105 16255 35139
rect 16405 35105 16439 35139
rect 17049 35105 17083 35139
rect 18797 35105 18831 35139
rect 18889 35105 18923 35139
rect 19533 35105 19567 35139
rect 19717 35105 19751 35139
rect 19809 35105 19843 35139
rect 24593 35105 24627 35139
rect 24777 35105 24811 35139
rect 25237 35105 25271 35139
rect 25421 35105 25455 35139
rect 26985 35105 27019 35139
rect 28181 35105 28215 35139
rect 28319 35105 28353 35139
rect 29653 35105 29687 35139
rect 29745 35105 29779 35139
rect 30113 35105 30147 35139
rect 30481 35105 30515 35139
rect 30573 35105 30607 35139
rect 31125 35105 31159 35139
rect 9689 35037 9723 35071
rect 9873 35037 9907 35071
rect 12633 35037 12667 35071
rect 12817 35037 12851 35071
rect 22937 35037 22971 35071
rect 23121 35037 23155 35071
rect 28457 35037 28491 35071
rect 29193 35037 29227 35071
rect 29377 35037 29411 35071
rect 30849 35037 30883 35071
rect 14933 34969 14967 35003
rect 19625 34969 19659 35003
rect 24777 34969 24811 35003
rect 28733 34969 28767 35003
rect 29469 34969 29503 35003
rect 30205 34969 30239 35003
rect 31033 34969 31067 35003
rect 10333 34901 10367 34935
rect 13093 34901 13127 34935
rect 14013 34901 14047 34935
rect 18797 34901 18831 34935
rect 19349 34901 19383 34935
rect 22017 34901 22051 34935
rect 27261 34901 27295 34935
rect 27445 34901 27479 34935
rect 30757 34901 30791 34935
rect 9781 34697 9815 34731
rect 13369 34697 13403 34731
rect 20729 34697 20763 34731
rect 22569 34697 22603 34731
rect 23949 34697 23983 34731
rect 24133 34697 24167 34731
rect 28365 34697 28399 34731
rect 30389 34697 30423 34731
rect 30665 34697 30699 34731
rect 15025 34629 15059 34663
rect 16313 34629 16347 34663
rect 18429 34629 18463 34663
rect 25053 34629 25087 34663
rect 8125 34561 8159 34595
rect 8401 34561 8435 34595
rect 12541 34561 12575 34595
rect 13645 34561 13679 34595
rect 15761 34561 15795 34595
rect 15920 34561 15954 34595
rect 16957 34561 16991 34595
rect 18797 34561 18831 34595
rect 18981 34561 19015 34595
rect 19073 34561 19107 34595
rect 21189 34561 21223 34595
rect 25973 34561 26007 34595
rect 8217 34493 8251 34527
rect 10057 34493 10091 34527
rect 10149 34493 10183 34527
rect 10333 34493 10367 34527
rect 10425 34493 10459 34527
rect 12449 34493 12483 34527
rect 12725 34493 12759 34527
rect 12909 34493 12943 34527
rect 13001 34493 13035 34527
rect 13093 34493 13127 34527
rect 13912 34493 13946 34527
rect 15117 34493 15151 34527
rect 16037 34493 16071 34527
rect 16773 34493 16807 34527
rect 18337 34493 18371 34527
rect 18705 34493 18739 34527
rect 19329 34493 19363 34527
rect 20637 34493 20671 34527
rect 20821 34493 20855 34527
rect 20913 34493 20947 34527
rect 22109 34493 22143 34527
rect 22293 34493 22327 34527
rect 23305 34493 23339 34527
rect 23673 34493 23707 34527
rect 24685 34493 24719 34527
rect 24777 34493 24811 34527
rect 25053 34493 25087 34527
rect 26709 34493 26743 34527
rect 26801 34493 26835 34527
rect 26985 34493 27019 34527
rect 28641 34493 28675 34527
rect 28733 34493 28767 34527
rect 29009 34493 29043 34527
rect 31309 34493 31343 34527
rect 8668 34425 8702 34459
rect 18981 34425 19015 34459
rect 22569 34425 22603 34459
rect 24133 34425 24167 34459
rect 24317 34425 24351 34459
rect 25145 34425 25179 34459
rect 27252 34425 27286 34459
rect 29276 34425 29310 34459
rect 9873 34357 9907 34391
rect 20453 34357 20487 34391
rect 21925 34357 21959 34391
rect 22385 34357 22419 34391
rect 23581 34357 23615 34391
rect 24593 34357 24627 34391
rect 24869 34357 24903 34391
rect 8861 34153 8895 34187
rect 9597 34153 9631 34187
rect 14473 34153 14507 34187
rect 18153 34153 18187 34187
rect 18245 34153 18279 34187
rect 19257 34153 19291 34187
rect 21649 34153 21683 34187
rect 29193 34153 29227 34187
rect 31309 34153 31343 34187
rect 9965 34085 9999 34119
rect 11161 34085 11195 34119
rect 13185 34085 13219 34119
rect 13277 34085 13311 34119
rect 13645 34085 13679 34119
rect 15393 34085 15427 34119
rect 16865 34085 16899 34119
rect 27353 34085 27387 34119
rect 27721 34085 27755 34119
rect 29009 34085 29043 34119
rect 30196 34085 30230 34119
rect 9137 34017 9171 34051
rect 9229 34017 9263 34051
rect 9321 34017 9355 34051
rect 9505 34017 9539 34051
rect 9781 34017 9815 34051
rect 11345 34017 11379 34051
rect 13001 34017 13035 34051
rect 13461 34017 13495 34051
rect 14105 34017 14139 34051
rect 14841 34017 14875 34051
rect 15485 34017 15519 34051
rect 15699 34017 15733 34051
rect 15853 34017 15887 34051
rect 16497 34017 16531 34051
rect 16589 34017 16623 34051
rect 18337 34017 18371 34051
rect 18429 34017 18463 34051
rect 18521 34017 18555 34051
rect 18889 34017 18923 34051
rect 19073 34017 19107 34051
rect 19533 34017 19567 34051
rect 19809 34017 19843 34051
rect 22477 34017 22511 34051
rect 22733 34017 22767 34051
rect 24593 34017 24627 34051
rect 24860 34017 24894 34051
rect 26249 34017 26283 34051
rect 27169 34017 27203 34051
rect 28641 34017 28675 34051
rect 29469 34017 29503 34051
rect 29745 34017 29779 34051
rect 29929 34017 29963 34051
rect 13921 33949 13955 33983
rect 14013 33949 14047 33983
rect 17601 33949 17635 33983
rect 18061 33949 18095 33983
rect 18981 33949 19015 33983
rect 21741 33949 21775 33983
rect 21833 33949 21867 33983
rect 26985 33949 27019 33983
rect 29285 33949 29319 33983
rect 29561 33949 29595 33983
rect 29653 33949 29687 33983
rect 15117 33881 15151 33915
rect 25973 33881 26007 33915
rect 27905 33881 27939 33915
rect 11529 33813 11563 33847
rect 14657 33813 14691 33847
rect 14933 33813 14967 33847
rect 16313 33813 16347 33847
rect 16681 33813 16715 33847
rect 18705 33813 18739 33847
rect 19717 33813 19751 33847
rect 21281 33813 21315 33847
rect 23857 33813 23891 33847
rect 26157 33813 26191 33847
rect 26433 33813 26467 33847
rect 27537 33813 27571 33847
rect 29009 33813 29043 33847
rect 13829 33609 13863 33643
rect 16129 33609 16163 33643
rect 18889 33609 18923 33643
rect 21741 33609 21775 33643
rect 23857 33609 23891 33643
rect 27353 33609 27387 33643
rect 18797 33541 18831 33575
rect 21649 33541 21683 33575
rect 28365 33541 28399 33575
rect 16865 33473 16899 33507
rect 20085 33473 20119 33507
rect 20269 33473 20303 33507
rect 25973 33473 26007 33507
rect 28457 33473 28491 33507
rect 9229 33405 9263 33439
rect 10609 33405 10643 33439
rect 10701 33405 10735 33439
rect 10793 33405 10827 33439
rect 10977 33405 11011 33439
rect 11345 33405 11379 33439
rect 11437 33405 11471 33439
rect 11529 33405 11563 33439
rect 11713 33405 11747 33439
rect 11989 33405 12023 33439
rect 12173 33405 12207 33439
rect 12265 33405 12299 33439
rect 12449 33402 12483 33436
rect 12541 33405 12575 33439
rect 12633 33405 12667 33439
rect 14013 33405 14047 33439
rect 14197 33405 14231 33439
rect 16405 33405 16439 33439
rect 16497 33405 16531 33439
rect 16589 33405 16623 33439
rect 16773 33405 16807 33439
rect 18705 33405 18739 33439
rect 20177 33405 20211 33439
rect 22385 33405 22419 33439
rect 23489 33405 23523 33439
rect 24133 33405 24167 33439
rect 24225 33405 24259 33439
rect 24317 33405 24351 33439
rect 24409 33405 24443 33439
rect 24593 33405 24627 33439
rect 25789 33405 25823 33439
rect 28089 33405 28123 33439
rect 28641 33405 28675 33439
rect 28733 33405 28767 33439
rect 9413 33337 9447 33371
rect 11805 33337 11839 33371
rect 17132 33337 17166 33371
rect 19073 33337 19107 33371
rect 20536 33337 20570 33371
rect 22661 33337 22695 33371
rect 26240 33337 26274 33371
rect 28365 33337 28399 33371
rect 28457 33337 28491 33371
rect 9597 33269 9631 33303
rect 10333 33269 10367 33303
rect 11069 33269 11103 33303
rect 12909 33269 12943 33303
rect 18245 33269 18279 33303
rect 18981 33269 19015 33303
rect 28181 33269 28215 33303
rect 10425 33065 10459 33099
rect 13093 33065 13127 33099
rect 16773 33065 16807 33099
rect 18889 33065 18923 33099
rect 20085 33065 20119 33099
rect 22569 33065 22603 33099
rect 24225 33065 24259 33099
rect 24777 33065 24811 33099
rect 26433 33065 26467 33099
rect 26617 33065 26651 33099
rect 29101 33065 29135 33099
rect 9321 32997 9355 33031
rect 10517 32997 10551 33031
rect 12725 32997 12759 33031
rect 14197 32997 14231 33031
rect 15025 32997 15059 33031
rect 19625 32997 19659 33031
rect 27997 32997 28031 33031
rect 8861 32929 8895 32963
rect 8953 32929 8987 32963
rect 9137 32929 9171 32963
rect 9229 32929 9263 32963
rect 9597 32929 9631 32963
rect 9689 32929 9723 32963
rect 9781 32929 9815 32963
rect 9965 32929 9999 32963
rect 11529 32929 11563 32963
rect 11621 32929 11655 32963
rect 13369 32929 13403 32963
rect 13461 32929 13495 32963
rect 13645 32929 13679 32963
rect 13737 32929 13771 32963
rect 15393 32929 15427 32963
rect 16865 32929 16899 32963
rect 19103 32929 19137 32963
rect 19257 32929 19291 32963
rect 19901 32929 19935 32963
rect 22201 32929 22235 32963
rect 22385 32929 22419 32963
rect 24225 32929 24259 32963
rect 24409 32929 24443 32963
rect 24961 32929 24995 32963
rect 25237 32929 25271 32963
rect 25605 32929 25639 32963
rect 26157 32929 26191 32963
rect 26985 32929 27019 32963
rect 28365 32929 28399 32963
rect 29653 32929 29687 32963
rect 10609 32861 10643 32895
rect 11713 32861 11747 32895
rect 12449 32861 12483 32895
rect 12633 32861 12667 32895
rect 16313 32861 16347 32895
rect 16405 32861 16439 32895
rect 16497 32861 16531 32895
rect 16589 32861 16623 32895
rect 19717 32861 19751 32895
rect 25145 32861 25179 32895
rect 25421 32861 25455 32895
rect 25881 32861 25915 32895
rect 15209 32793 15243 32827
rect 25973 32793 26007 32827
rect 27629 32793 27663 32827
rect 8677 32725 8711 32759
rect 10057 32725 10091 32759
rect 11161 32725 11195 32759
rect 13185 32725 13219 32759
rect 19809 32725 19843 32759
rect 25789 32725 25823 32759
rect 26617 32725 26651 32759
rect 27537 32725 27571 32759
rect 29009 32725 29043 32759
rect 9413 32521 9447 32555
rect 15853 32521 15887 32555
rect 17141 32521 17175 32555
rect 17693 32521 17727 32555
rect 22477 32521 22511 32555
rect 28825 32521 28859 32555
rect 20913 32453 20947 32487
rect 10057 32385 10091 32419
rect 14289 32385 14323 32419
rect 14473 32385 14507 32419
rect 16129 32385 16163 32419
rect 16221 32385 16255 32419
rect 16405 32385 16439 32419
rect 20637 32385 20671 32419
rect 22017 32385 22051 32419
rect 9781 32317 9815 32351
rect 10425 32317 10459 32351
rect 10517 32317 10551 32351
rect 10701 32317 10735 32351
rect 10793 32317 10827 32351
rect 10977 32317 11011 32351
rect 11069 32317 11103 32351
rect 11253 32317 11287 32351
rect 11345 32317 11379 32351
rect 12357 32317 12391 32351
rect 12541 32317 12575 32351
rect 12633 32317 12667 32351
rect 12725 32317 12759 32351
rect 14381 32317 14415 32351
rect 16313 32317 16347 32351
rect 17417 32317 17451 32351
rect 17601 32317 17635 32351
rect 17877 32317 17911 32351
rect 19625 32317 19659 32351
rect 20177 32317 20211 32351
rect 20270 32317 20304 32351
rect 20717 32317 20751 32351
rect 21189 32317 21223 32351
rect 21281 32317 21315 32351
rect 21741 32317 21775 32351
rect 22201 32317 22235 32351
rect 22661 32317 22695 32351
rect 22753 32317 22787 32351
rect 22845 32317 22879 32351
rect 22983 32317 23017 32351
rect 23121 32317 23155 32351
rect 23397 32317 23431 32351
rect 25237 32317 25271 32351
rect 27169 32317 27203 32351
rect 27261 32317 27295 32351
rect 27445 32317 27479 32351
rect 29009 32317 29043 32351
rect 14740 32249 14774 32283
rect 16957 32249 16991 32283
rect 17173 32249 17207 32283
rect 19993 32249 20027 32283
rect 20361 32249 20395 32283
rect 20499 32249 20533 32283
rect 27712 32249 27746 32283
rect 9873 32181 9907 32215
rect 10241 32181 10275 32215
rect 11529 32181 11563 32215
rect 13001 32181 13035 32215
rect 15945 32181 15979 32215
rect 17325 32181 17359 32215
rect 17509 32181 17543 32215
rect 19717 32181 19751 32215
rect 21465 32181 21499 32215
rect 21649 32181 21683 32215
rect 22385 32181 22419 32215
rect 23305 32181 23339 32215
rect 25329 32181 25363 32215
rect 29101 32181 29135 32215
rect 10793 31977 10827 32011
rect 14933 31977 14967 32011
rect 15669 31977 15703 32011
rect 16497 31977 16531 32011
rect 20913 31977 20947 32011
rect 24225 31977 24259 32011
rect 27997 31977 28031 32011
rect 10425 31909 10459 31943
rect 10609 31909 10643 31943
rect 16665 31909 16699 31943
rect 16865 31909 16899 31943
rect 16957 31909 16991 31943
rect 19073 31909 19107 31943
rect 19778 31909 19812 31943
rect 24685 31909 24719 31943
rect 29110 31909 29144 31943
rect 9137 31841 9171 31875
rect 12633 31841 12667 31875
rect 13553 31841 13587 31875
rect 13691 31841 13725 31875
rect 15209 31841 15243 31875
rect 15301 31841 15335 31875
rect 15393 31841 15427 31875
rect 15577 31841 15611 31875
rect 15853 31841 15887 31875
rect 17141 31841 17175 31875
rect 17509 31841 17543 31875
rect 17877 31841 17911 31875
rect 17969 31841 18003 31875
rect 18981 31841 19015 31875
rect 19165 31841 19199 31875
rect 19533 31841 19567 31875
rect 21281 31841 21315 31875
rect 21548 31841 21582 31875
rect 22753 31841 22787 31875
rect 23009 31841 23043 31875
rect 24409 31841 24443 31875
rect 26433 31841 26467 31875
rect 26617 31841 26651 31875
rect 29377 31841 29411 31875
rect 12817 31773 12851 31807
rect 13277 31773 13311 31807
rect 13829 31773 13863 31807
rect 17325 31773 17359 31807
rect 24501 31773 24535 31807
rect 24133 31705 24167 31739
rect 9045 31637 9079 31671
rect 14473 31637 14507 31671
rect 16681 31637 16715 31671
rect 17693 31637 17727 31671
rect 22661 31637 22695 31671
rect 24685 31637 24719 31671
rect 26525 31637 26559 31671
rect 11713 31433 11747 31467
rect 14933 31433 14967 31467
rect 21281 31433 21315 31467
rect 22385 31433 22419 31467
rect 17049 31365 17083 31399
rect 15301 31297 15335 31331
rect 15485 31297 15519 31331
rect 16313 31297 16347 31331
rect 17877 31297 17911 31331
rect 21465 31297 21499 31331
rect 22109 31297 22143 31331
rect 23581 31297 23615 31331
rect 24225 31297 24259 31331
rect 25973 31297 26007 31331
rect 26433 31297 26467 31331
rect 8953 31229 8987 31263
rect 9045 31229 9079 31263
rect 9137 31229 9171 31263
rect 9321 31229 9355 31263
rect 9689 31229 9723 31263
rect 9781 31229 9815 31263
rect 9873 31229 9907 31263
rect 10057 31229 10091 31263
rect 10793 31229 10827 31263
rect 10977 31229 11011 31263
rect 11069 31229 11103 31263
rect 11161 31229 11195 31263
rect 11989 31229 12023 31263
rect 12081 31229 12115 31263
rect 12173 31229 12207 31263
rect 12357 31229 12391 31263
rect 13185 31229 13219 31263
rect 13277 31229 13311 31263
rect 13553 31229 13587 31263
rect 13820 31229 13854 31263
rect 15393 31229 15427 31263
rect 15761 31229 15795 31263
rect 15853 31229 15887 31263
rect 16037 31229 16071 31263
rect 16129 31229 16163 31263
rect 17601 31229 17635 31263
rect 17785 31229 17819 31263
rect 17969 31229 18003 31263
rect 18153 31229 18187 31263
rect 18705 31229 18739 31263
rect 20821 31229 20855 31263
rect 21005 31229 21039 31263
rect 21373 31229 21407 31263
rect 21649 31229 21683 31263
rect 21741 31229 21775 31263
rect 22569 31229 22603 31263
rect 22753 31229 22787 31263
rect 23029 31229 23063 31263
rect 23489 31229 23523 31263
rect 23949 31229 23983 31263
rect 26065 31229 26099 31263
rect 27353 31229 27387 31263
rect 27445 31229 27479 31263
rect 27629 31229 27663 31263
rect 17325 31161 17359 31195
rect 18337 31161 18371 31195
rect 18950 31161 18984 31195
rect 21097 31161 21131 31195
rect 21833 31161 21867 31195
rect 21951 31161 21985 31195
rect 22661 31161 22695 31195
rect 22891 31161 22925 31195
rect 24470 31161 24504 31195
rect 26525 31161 26559 31195
rect 26709 31161 26743 31195
rect 27169 31161 27203 31195
rect 8677 31093 8711 31127
rect 9413 31093 9447 31127
rect 11437 31093 11471 31127
rect 15669 31093 15703 31127
rect 16865 31093 16899 31127
rect 20085 31093 20119 31127
rect 24041 31093 24075 31127
rect 25605 31093 25639 31127
rect 26893 31093 26927 31127
rect 26985 31093 27019 31127
rect 27537 31093 27571 31127
rect 10241 30889 10275 30923
rect 12817 30889 12851 30923
rect 13553 30889 13587 30923
rect 15853 30889 15887 30923
rect 16221 30889 16255 30923
rect 18245 30889 18279 30923
rect 19073 30889 19107 30923
rect 23673 30889 23707 30923
rect 9106 30821 9140 30855
rect 13921 30821 13955 30855
rect 15393 30821 15427 30855
rect 24133 30821 24167 30855
rect 24470 30821 24504 30855
rect 26709 30821 26743 30855
rect 26801 30821 26835 30855
rect 28089 30821 28123 30855
rect 8861 30753 8895 30787
rect 11161 30753 11195 30787
rect 11897 30753 11931 30787
rect 13277 30753 13311 30787
rect 13369 30753 13403 30787
rect 13737 30753 13771 30787
rect 14197 30753 14231 30787
rect 14565 30753 14599 30787
rect 14933 30753 14967 30787
rect 15577 30753 15611 30787
rect 15761 30753 15795 30787
rect 16497 30753 16531 30787
rect 16773 30753 16807 30787
rect 16957 30753 16991 30787
rect 18797 30753 18831 30787
rect 19165 30753 19199 30787
rect 23305 30753 23339 30787
rect 23489 30753 23523 30787
rect 23765 30753 23799 30787
rect 23949 30753 23983 30787
rect 24225 30753 24259 30787
rect 26433 30753 26467 30787
rect 26526 30753 26560 30787
rect 26939 30753 26973 30787
rect 27905 30753 27939 30787
rect 10977 30685 11011 30719
rect 11621 30685 11655 30719
rect 12035 30685 12069 30719
rect 12173 30685 12207 30719
rect 17141 30685 17175 30719
rect 17601 30685 17635 30719
rect 17233 30617 17267 30651
rect 16589 30549 16623 30583
rect 16681 30549 16715 30583
rect 25605 30549 25639 30583
rect 27077 30549 27111 30583
rect 27721 30549 27755 30583
rect 10701 30345 10735 30379
rect 15577 30345 15611 30379
rect 15945 30345 15979 30379
rect 16681 30345 16715 30379
rect 23857 30345 23891 30379
rect 12449 30277 12483 30311
rect 16221 30277 16255 30311
rect 16589 30277 16623 30311
rect 17049 30277 17083 30311
rect 25237 30277 25271 30311
rect 15853 30209 15887 30243
rect 17785 30209 17819 30243
rect 24501 30209 24535 30243
rect 24593 30209 24627 30243
rect 9045 30141 9079 30175
rect 9137 30141 9171 30175
rect 9321 30141 9355 30175
rect 10793 30141 10827 30175
rect 10885 30141 10919 30175
rect 11069 30141 11103 30175
rect 11336 30141 11370 30175
rect 14381 30141 14415 30175
rect 15945 30141 15979 30175
rect 16497 30141 16531 30175
rect 16773 30141 16807 30175
rect 16957 30141 16991 30175
rect 17233 30141 17267 30175
rect 17325 30141 17359 30175
rect 17509 30141 17543 30175
rect 17601 30141 17635 30175
rect 17877 30141 17911 30175
rect 19257 30141 19291 30175
rect 24041 30141 24075 30175
rect 24869 30141 24903 30175
rect 25053 30141 25087 30175
rect 27169 30141 27203 30175
rect 27261 30141 27295 30175
rect 27445 30141 27479 30175
rect 9588 30073 9622 30107
rect 24133 30073 24167 30107
rect 24225 30073 24259 30107
rect 24343 30073 24377 30107
rect 24731 30073 24765 30107
rect 24961 30073 24995 30107
rect 27690 30073 27724 30107
rect 14289 30005 14323 30039
rect 19165 30005 19199 30039
rect 28825 30005 28859 30039
rect 16773 29801 16807 29835
rect 17601 29801 17635 29835
rect 18613 29801 18647 29835
rect 20361 29801 20395 29835
rect 27629 29801 27663 29835
rect 27813 29801 27847 29835
rect 17233 29733 17267 29767
rect 17433 29733 17467 29767
rect 17785 29733 17819 29767
rect 26433 29733 26467 29767
rect 14105 29665 14139 29699
rect 14372 29665 14406 29699
rect 16405 29665 16439 29699
rect 16865 29665 16899 29699
rect 17693 29665 17727 29699
rect 17969 29665 18003 29699
rect 18245 29665 18279 29699
rect 18613 29665 18647 29699
rect 18981 29665 19015 29699
rect 19248 29665 19282 29699
rect 20729 29665 20763 29699
rect 21741 29665 21775 29699
rect 21833 29665 21867 29699
rect 22017 29665 22051 29699
rect 22293 29665 22327 29699
rect 22385 29665 22419 29699
rect 22753 29665 22787 29699
rect 23581 29665 23615 29699
rect 23857 29665 23891 29699
rect 25237 29665 25271 29699
rect 25330 29665 25364 29699
rect 26709 29665 26743 29699
rect 28457 29665 28491 29699
rect 16589 29597 16623 29631
rect 18797 29597 18831 29631
rect 26617 29597 26651 29631
rect 26801 29597 26835 29631
rect 26893 29597 26927 29631
rect 28641 29597 28675 29631
rect 15485 29529 15519 29563
rect 23765 29529 23799 29563
rect 25605 29529 25639 29563
rect 28181 29529 28215 29563
rect 28273 29529 28307 29563
rect 16129 29461 16163 29495
rect 16497 29461 16531 29495
rect 17417 29461 17451 29495
rect 18153 29461 18187 29495
rect 20637 29461 20671 29495
rect 22109 29461 22143 29495
rect 22661 29461 22695 29495
rect 23397 29461 23431 29495
rect 27813 29461 27847 29495
rect 14749 29257 14783 29291
rect 17509 29257 17543 29291
rect 18153 29257 18187 29291
rect 19625 29257 19659 29291
rect 26065 29257 26099 29291
rect 11437 29189 11471 29223
rect 17325 29189 17359 29223
rect 25881 29189 25915 29223
rect 14657 29121 14691 29155
rect 20453 29121 20487 29155
rect 23673 29121 23707 29155
rect 24225 29121 24259 29155
rect 25789 29121 25823 29155
rect 27813 29121 27847 29155
rect 11253 29053 11287 29087
rect 11437 29053 11471 29087
rect 11713 29053 11747 29087
rect 12357 29053 12391 29087
rect 12817 29053 12851 29087
rect 13093 29053 13127 29087
rect 13185 29053 13219 29087
rect 13369 29053 13403 29087
rect 14197 29053 14231 29087
rect 14289 29053 14323 29087
rect 15025 29053 15059 29087
rect 15117 29053 15151 29087
rect 15209 29053 15243 29087
rect 15393 29053 15427 29087
rect 18337 29053 18371 29087
rect 19349 29053 19383 29087
rect 19533 29053 19567 29087
rect 19901 29053 19935 29087
rect 20177 29053 20211 29087
rect 21925 29053 21959 29087
rect 23857 29053 23891 29087
rect 24041 29053 24075 29087
rect 25145 29053 25179 29087
rect 25238 29053 25272 29087
rect 25513 29053 25547 29087
rect 25697 29053 25731 29087
rect 25881 29053 25915 29087
rect 26157 29053 26191 29087
rect 28457 29053 28491 29087
rect 11621 28985 11655 29019
rect 13001 28985 13035 29019
rect 13553 28985 13587 29019
rect 14473 28985 14507 29019
rect 17049 28985 17083 29019
rect 18521 28985 18555 29019
rect 19809 28985 19843 29019
rect 20085 28985 20119 29019
rect 20698 28985 20732 29019
rect 22192 28985 22226 29019
rect 23489 28985 23523 29019
rect 27997 28985 28031 29019
rect 28181 28985 28215 29019
rect 28365 28985 28399 29019
rect 11161 28917 11195 28951
rect 12449 28917 12483 28951
rect 12633 28917 12667 28951
rect 13185 28917 13219 28951
rect 21833 28917 21867 28951
rect 23305 28917 23339 28951
rect 12357 28713 12391 28747
rect 14289 28713 14323 28747
rect 14933 28713 14967 28747
rect 15577 28713 15611 28747
rect 15745 28713 15779 28747
rect 16865 28713 16899 28747
rect 17417 28713 17451 28747
rect 20545 28713 20579 28747
rect 22753 28713 22787 28747
rect 27169 28713 27203 28747
rect 14197 28645 14231 28679
rect 15117 28645 15151 28679
rect 15945 28645 15979 28679
rect 21649 28645 21683 28679
rect 23388 28645 23422 28679
rect 25605 28645 25639 28679
rect 10977 28577 11011 28611
rect 11244 28577 11278 28611
rect 12541 28577 12575 28611
rect 12817 28577 12851 28611
rect 14657 28577 14691 28611
rect 15301 28577 15335 28611
rect 16773 28577 16807 28611
rect 16957 28577 16991 28611
rect 17325 28577 17359 28611
rect 17509 28577 17543 28611
rect 17877 28577 17911 28611
rect 18061 28577 18095 28611
rect 20177 28577 20211 28611
rect 20729 28577 20763 28611
rect 21281 28577 21315 28611
rect 21465 28577 21499 28611
rect 21557 28577 21591 28611
rect 21767 28577 21801 28611
rect 21925 28577 21959 28611
rect 22109 28577 22143 28611
rect 22247 28577 22281 28611
rect 22385 28577 22419 28611
rect 22477 28577 22511 28611
rect 22569 28577 22603 28611
rect 23121 28577 23155 28611
rect 25329 28577 25363 28611
rect 25421 28577 25455 28611
rect 25973 28577 26007 28611
rect 26433 28577 26467 28611
rect 26617 28577 26651 28611
rect 26893 28577 26927 28611
rect 28834 28577 28868 28611
rect 29101 28577 29135 28611
rect 14473 28509 14507 28543
rect 14565 28509 14599 28543
rect 14749 28509 14783 28543
rect 20361 28509 20395 28543
rect 20913 28509 20947 28543
rect 25697 28509 25731 28543
rect 26065 28509 26099 28543
rect 15761 28373 15795 28407
rect 17969 28373 18003 28407
rect 19993 28373 20027 28407
rect 24501 28373 24535 28407
rect 26249 28373 26283 28407
rect 26709 28373 26743 28407
rect 26801 28373 26835 28407
rect 27721 28373 27755 28407
rect 11437 28169 11471 28203
rect 13737 28169 13771 28203
rect 15853 28169 15887 28203
rect 17509 28169 17543 28203
rect 19625 28169 19659 28203
rect 23857 28169 23891 28203
rect 24777 28169 24811 28203
rect 25789 28169 25823 28203
rect 28089 28169 28123 28203
rect 28273 28169 28307 28203
rect 15945 28101 15979 28135
rect 17325 28101 17359 28135
rect 17693 28101 17727 28135
rect 16865 28033 16899 28067
rect 17969 28033 18003 28067
rect 24777 28033 24811 28067
rect 11345 27965 11379 27999
rect 11529 27965 11563 27999
rect 11713 27965 11747 27999
rect 12081 27965 12115 27999
rect 13553 27965 13587 27999
rect 13645 27965 13679 27999
rect 15301 27965 15335 27999
rect 15669 27965 15703 27999
rect 16129 27965 16163 27999
rect 16221 27965 16255 27999
rect 16313 27965 16347 27999
rect 16405 27965 16439 27999
rect 16589 27965 16623 27999
rect 18981 27965 19015 27999
rect 20913 27965 20947 27999
rect 22293 27965 22327 27999
rect 24041 27965 24075 27999
rect 24133 27965 24167 27999
rect 24225 27965 24259 27999
rect 24501 27965 24535 27999
rect 24869 27965 24903 27999
rect 25605 27965 25639 27999
rect 25759 27965 25793 27999
rect 27721 27965 27755 27999
rect 11897 27897 11931 27931
rect 13829 27897 13863 27931
rect 15485 27897 15519 27931
rect 15577 27897 15611 27931
rect 17325 27897 17359 27931
rect 24343 27897 24377 27931
rect 24593 27897 24627 27931
rect 28089 27897 28123 27931
rect 16773 27829 16807 27863
rect 18889 27829 18923 27863
rect 22201 27829 22235 27863
rect 25053 27829 25087 27863
rect 14381 27625 14415 27659
rect 25053 27625 25087 27659
rect 27530 27625 27564 27659
rect 11897 27557 11931 27591
rect 16773 27557 16807 27591
rect 18245 27557 18279 27591
rect 21649 27557 21683 27591
rect 21741 27557 21775 27591
rect 22201 27557 22235 27591
rect 25329 27557 25363 27591
rect 27445 27557 27479 27591
rect 27721 27557 27755 27591
rect 11713 27489 11747 27523
rect 11989 27489 12023 27523
rect 12081 27489 12115 27523
rect 13737 27489 13771 27523
rect 13830 27489 13864 27523
rect 14013 27489 14047 27523
rect 14105 27489 14139 27523
rect 14243 27489 14277 27523
rect 14473 27489 14507 27523
rect 14657 27489 14691 27523
rect 16681 27489 16715 27523
rect 16865 27489 16899 27523
rect 18705 27489 18739 27523
rect 18961 27489 18995 27523
rect 20453 27489 20487 27523
rect 20545 27489 20579 27523
rect 21005 27489 21039 27523
rect 21557 27489 21591 27523
rect 21879 27489 21913 27523
rect 23857 27489 23891 27523
rect 24041 27489 24075 27523
rect 24501 27489 24535 27523
rect 24777 27489 24811 27523
rect 25053 27489 25087 27523
rect 25145 27489 25179 27523
rect 26985 27489 27019 27523
rect 27353 27489 27387 27523
rect 27629 27489 27663 27523
rect 28549 27489 28583 27523
rect 12357 27421 12391 27455
rect 14565 27421 14599 27455
rect 15393 27421 15427 27455
rect 15853 27421 15887 27455
rect 17969 27421 18003 27455
rect 18153 27421 18187 27455
rect 22017 27421 22051 27455
rect 22845 27421 22879 27455
rect 23765 27421 23799 27455
rect 24593 27421 24627 27455
rect 25789 27421 25823 27455
rect 26893 27421 26927 27455
rect 28273 27421 28307 27455
rect 12173 27353 12207 27387
rect 12265 27353 12299 27387
rect 15669 27353 15703 27387
rect 18613 27353 18647 27387
rect 24961 27353 24995 27387
rect 26065 27353 26099 27387
rect 26525 27353 26559 27387
rect 11529 27285 11563 27319
rect 20085 27285 20119 27319
rect 20269 27285 20303 27319
rect 20821 27285 20855 27319
rect 21373 27285 21407 27319
rect 23121 27285 23155 27319
rect 24225 27285 24259 27319
rect 24593 27285 24627 27319
rect 26249 27285 26283 27319
rect 26433 27285 26467 27319
rect 27077 27285 27111 27319
rect 29101 27285 29135 27319
rect 12541 27081 12575 27115
rect 14565 27081 14599 27115
rect 21097 27081 21131 27115
rect 26341 27081 26375 27115
rect 26433 27081 26467 27115
rect 26801 27081 26835 27115
rect 14381 27013 14415 27047
rect 25881 27013 25915 27047
rect 10977 26945 11011 26979
rect 11161 26945 11195 26979
rect 19533 26945 19567 26979
rect 19717 26945 19751 26979
rect 25973 26945 26007 26979
rect 26525 26945 26559 26979
rect 28825 26945 28859 26979
rect 29101 26945 29135 26979
rect 11069 26877 11103 26911
rect 11428 26877 11462 26911
rect 14197 26877 14231 26911
rect 14289 26877 14323 26911
rect 14565 26877 14599 26911
rect 14749 26877 14783 26911
rect 17509 26877 17543 26911
rect 18245 26877 18279 26911
rect 19257 26877 19291 26911
rect 19625 26877 19659 26911
rect 19984 26877 20018 26911
rect 21189 26877 21223 26911
rect 21456 26877 21490 26911
rect 22845 26877 22879 26911
rect 22937 26877 22971 26911
rect 23029 26877 23063 26911
rect 23305 26877 23339 26911
rect 23489 26877 23523 26911
rect 23581 26877 23615 26911
rect 23857 26877 23891 26911
rect 24124 26877 24158 26911
rect 26065 26877 26099 26911
rect 26249 26877 26283 26911
rect 26893 26877 26927 26911
rect 29009 26877 29043 26911
rect 14473 26809 14507 26843
rect 23147 26809 23181 26843
rect 25513 26809 25547 26843
rect 28580 26809 28614 26843
rect 16957 26741 16991 26775
rect 17693 26741 17727 26775
rect 18705 26741 18739 26775
rect 22569 26741 22603 26775
rect 22661 26741 22695 26775
rect 25237 26741 25271 26775
rect 26985 26741 27019 26775
rect 27445 26741 27479 26775
rect 14473 26537 14507 26571
rect 14749 26537 14783 26571
rect 17049 26537 17083 26571
rect 17417 26537 17451 26571
rect 17509 26537 17543 26571
rect 18245 26537 18279 26571
rect 18337 26537 18371 26571
rect 19073 26537 19107 26571
rect 19717 26537 19751 26571
rect 20269 26537 20303 26571
rect 21373 26537 21407 26571
rect 24133 26537 24167 26571
rect 27077 26537 27111 26571
rect 28365 26537 28399 26571
rect 15117 26469 15151 26503
rect 23627 26469 23661 26503
rect 23857 26469 23891 26503
rect 26709 26469 26743 26503
rect 26801 26469 26835 26503
rect 27629 26469 27663 26503
rect 27845 26469 27879 26503
rect 16773 26401 16807 26435
rect 20453 26401 20487 26435
rect 20545 26401 20579 26435
rect 20637 26401 20671 26435
rect 20775 26401 20809 26435
rect 21465 26401 21499 26435
rect 21741 26401 21775 26435
rect 22008 26401 22042 26435
rect 23765 26401 23799 26435
rect 23949 26401 23983 26435
rect 26433 26401 26467 26435
rect 26526 26401 26560 26435
rect 26898 26401 26932 26435
rect 28089 26401 28123 26435
rect 28181 26401 28215 26435
rect 12633 26333 12667 26367
rect 12817 26333 12851 26367
rect 13553 26333 13587 26367
rect 13670 26333 13704 26367
rect 13829 26333 13863 26367
rect 15209 26333 15243 26367
rect 15301 26333 15335 26367
rect 17693 26333 17727 26367
rect 18429 26333 18463 26367
rect 19165 26333 19199 26367
rect 19257 26333 19291 26367
rect 19533 26333 19567 26367
rect 19901 26333 19935 26367
rect 20913 26333 20947 26367
rect 23489 26333 23523 26367
rect 28365 26333 28399 26367
rect 13277 26265 13311 26299
rect 27997 26265 28031 26299
rect 16681 26197 16715 26231
rect 17877 26197 17911 26231
rect 18705 26197 18739 26231
rect 19901 26197 19935 26231
rect 23121 26197 23155 26231
rect 27813 26197 27847 26231
rect 13001 25993 13035 26027
rect 14473 25993 14507 26027
rect 15301 25993 15335 26027
rect 15853 25993 15887 26027
rect 18521 25993 18555 26027
rect 20361 25993 20395 26027
rect 13369 25925 13403 25959
rect 13001 25857 13035 25891
rect 13553 25857 13587 25891
rect 15025 25857 15059 25891
rect 15393 25857 15427 25891
rect 17969 25857 18003 25891
rect 12173 25789 12207 25823
rect 12909 25789 12943 25823
rect 13185 25789 13219 25823
rect 15577 25789 15611 25823
rect 15853 25789 15887 25823
rect 16037 25789 16071 25823
rect 16221 25789 16255 25823
rect 16497 25789 16531 25823
rect 16764 25789 16798 25823
rect 18337 25789 18371 25823
rect 18889 25789 18923 25823
rect 19073 25789 19107 25823
rect 19257 25789 19291 25823
rect 19809 25789 19843 25823
rect 27905 25789 27939 25823
rect 28181 25789 28215 25823
rect 14841 25721 14875 25755
rect 15301 25721 15335 25755
rect 27721 25721 27755 25755
rect 12081 25653 12115 25687
rect 14197 25653 14231 25687
rect 14933 25653 14967 25687
rect 15761 25653 15795 25687
rect 16313 25653 16347 25687
rect 17877 25653 17911 25687
rect 18153 25653 18187 25687
rect 18797 25653 18831 25687
rect 28089 25653 28123 25687
rect 13277 25449 13311 25483
rect 17877 25449 17911 25483
rect 24225 25449 24259 25483
rect 25697 25449 25731 25483
rect 14565 25381 14599 25415
rect 14749 25381 14783 25415
rect 14841 25381 14875 25415
rect 16764 25381 16798 25415
rect 18604 25381 18638 25415
rect 22753 25381 22787 25415
rect 23397 25381 23431 25415
rect 24593 25381 24627 25415
rect 25329 25381 25363 25415
rect 25421 25381 25455 25415
rect 11897 25313 11931 25347
rect 12164 25313 12198 25347
rect 13645 25313 13679 25347
rect 15025 25313 15059 25347
rect 15301 25313 15335 25347
rect 16405 25313 16439 25347
rect 16497 25313 16531 25347
rect 18337 25313 18371 25347
rect 20545 25313 20579 25347
rect 22201 25313 22235 25347
rect 22569 25313 22603 25347
rect 22661 25313 22695 25347
rect 22871 25313 22905 25347
rect 23259 25313 23293 25347
rect 23489 25313 23523 25347
rect 23581 25313 23615 25347
rect 23857 25313 23891 25347
rect 24501 25313 24535 25347
rect 25145 25313 25179 25347
rect 25513 25313 25547 25347
rect 27721 25313 27755 25347
rect 15945 25245 15979 25279
rect 23029 25245 23063 25279
rect 23121 25245 23155 25279
rect 23949 25245 23983 25279
rect 14381 25177 14415 25211
rect 14289 25109 14323 25143
rect 15209 25109 15243 25143
rect 16221 25109 16255 25143
rect 19717 25109 19751 25143
rect 20453 25109 20487 25143
rect 22109 25109 22143 25143
rect 22385 25109 22419 25143
rect 23765 25109 23799 25143
rect 24041 25109 24075 25143
rect 27629 25109 27663 25143
rect 13001 24905 13035 24939
rect 16037 24905 16071 24939
rect 23305 24905 23339 24939
rect 27261 24905 27295 24939
rect 28825 24905 28859 24939
rect 24869 24837 24903 24871
rect 17693 24769 17727 24803
rect 17785 24769 17819 24803
rect 18061 24769 18095 24803
rect 18245 24769 18279 24803
rect 20269 24769 20303 24803
rect 24501 24769 24535 24803
rect 25789 24769 25823 24803
rect 11345 24701 11379 24735
rect 11437 24701 11471 24735
rect 11621 24701 11655 24735
rect 13829 24701 13863 24735
rect 13921 24701 13955 24735
rect 14013 24701 14047 24735
rect 14197 24701 14231 24735
rect 14381 24701 14415 24735
rect 14473 24701 14507 24735
rect 14657 24701 14691 24735
rect 19073 24701 19107 24735
rect 19257 24701 19291 24735
rect 19809 24701 19843 24735
rect 21925 24701 21959 24735
rect 23397 24701 23431 24735
rect 24041 24701 24075 24735
rect 24225 24701 24259 24735
rect 25053 24701 25087 24735
rect 25237 24701 25271 24735
rect 25329 24701 25363 24735
rect 25421 24701 25455 24735
rect 25605 24701 25639 24735
rect 25881 24701 25915 24735
rect 26065 24701 26099 24735
rect 26157 24701 26191 24735
rect 26249 24701 26283 24735
rect 26433 24701 26467 24735
rect 26893 24701 26927 24735
rect 27445 24701 27479 24735
rect 11888 24633 11922 24667
rect 13553 24633 13587 24667
rect 14924 24633 14958 24667
rect 20514 24633 20548 24667
rect 22192 24633 22226 24667
rect 26709 24633 26743 24667
rect 27690 24633 27724 24667
rect 19993 24565 20027 24599
rect 21649 24565 21683 24599
rect 23489 24565 23523 24599
rect 23857 24565 23891 24599
rect 24961 24565 24995 24599
rect 26617 24565 26651 24599
rect 26985 24565 27019 24599
rect 27077 24565 27111 24599
rect 13093 24361 13127 24395
rect 20361 24361 20395 24395
rect 22017 24361 22051 24395
rect 22661 24361 22695 24395
rect 24685 24361 24719 24395
rect 25329 24361 25363 24395
rect 27537 24361 27571 24395
rect 27721 24361 27755 24395
rect 14473 24293 14507 24327
rect 14657 24293 14691 24327
rect 21557 24293 21591 24327
rect 21767 24293 21801 24327
rect 25697 24293 25731 24327
rect 26525 24293 26559 24327
rect 13369 24225 13403 24259
rect 13461 24225 13495 24259
rect 13553 24225 13587 24259
rect 13737 24225 13771 24259
rect 14197 24225 14231 24259
rect 14381 24225 14415 24259
rect 14841 24225 14875 24259
rect 15393 24225 15427 24259
rect 15485 24225 15519 24259
rect 15577 24225 15611 24259
rect 15761 24225 15795 24259
rect 16405 24225 16439 24259
rect 16589 24225 16623 24259
rect 20545 24225 20579 24259
rect 21281 24225 21315 24259
rect 21465 24225 21499 24259
rect 21649 24225 21683 24259
rect 22201 24225 22235 24259
rect 23774 24225 23808 24259
rect 24041 24225 24075 24259
rect 24317 24225 24351 24259
rect 24961 24225 24995 24259
rect 25421 24225 25455 24259
rect 25513 24225 25547 24259
rect 25789 24225 25823 24259
rect 25881 24225 25915 24259
rect 26249 24225 26283 24259
rect 26617 24225 26651 24259
rect 28181 24225 28215 24259
rect 28365 24225 28399 24259
rect 20729 24157 20763 24191
rect 21925 24157 21959 24191
rect 22385 24157 22419 24191
rect 24225 24157 24259 24191
rect 24869 24157 24903 24191
rect 26157 24157 26191 24191
rect 28089 24089 28123 24123
rect 14013 24021 14047 24055
rect 15117 24021 15151 24055
rect 16221 24021 16255 24055
rect 25421 24021 25455 24055
rect 27721 24021 27755 24055
rect 28549 24021 28583 24055
rect 16405 23817 16439 23851
rect 20361 23817 20395 23851
rect 26985 23817 27019 23851
rect 27905 23817 27939 23851
rect 28365 23817 28399 23851
rect 30389 23817 30423 23851
rect 13369 23681 13403 23715
rect 14289 23681 14323 23715
rect 27537 23681 27571 23715
rect 27997 23681 28031 23715
rect 12541 23613 12575 23647
rect 15393 23613 15427 23647
rect 15761 23613 15795 23647
rect 15853 23613 15887 23647
rect 15945 23613 15979 23647
rect 16129 23613 16163 23647
rect 16957 23613 16991 23647
rect 17141 23613 17175 23647
rect 18949 23613 18983 23647
rect 19073 23613 19107 23647
rect 19165 23613 19199 23647
rect 19349 23613 19383 23647
rect 20269 23613 20303 23647
rect 27077 23613 27111 23647
rect 27721 23613 27755 23647
rect 28641 23613 28675 23647
rect 28733 23613 28767 23647
rect 29009 23613 29043 23647
rect 13001 23545 13035 23579
rect 13185 23545 13219 23579
rect 14657 23545 14691 23579
rect 17693 23545 17727 23579
rect 17877 23545 17911 23579
rect 18061 23545 18095 23579
rect 29254 23545 29288 23579
rect 12449 23477 12483 23511
rect 13737 23477 13771 23511
rect 15485 23477 15519 23511
rect 17233 23477 17267 23511
rect 18705 23477 18739 23511
rect 19165 23477 19199 23511
rect 28365 23477 28399 23511
rect 28549 23477 28583 23511
rect 13645 23273 13679 23307
rect 16221 23273 16255 23307
rect 27537 23273 27571 23307
rect 12532 23205 12566 23239
rect 13737 23205 13771 23239
rect 22293 23205 22327 23239
rect 23121 23205 23155 23239
rect 25053 23205 25087 23239
rect 28149 23205 28183 23239
rect 28365 23205 28399 23239
rect 28549 23205 28583 23239
rect 12265 23137 12299 23171
rect 14013 23137 14047 23171
rect 14105 23137 14139 23171
rect 14197 23137 14231 23171
rect 14381 23137 14415 23171
rect 14657 23137 14691 23171
rect 17334 23137 17368 23171
rect 17601 23137 17635 23171
rect 17877 23137 17911 23171
rect 18889 23137 18923 23171
rect 19165 23137 19199 23171
rect 19533 23137 19567 23171
rect 19625 23137 19659 23171
rect 19901 23137 19935 23171
rect 20085 23137 20119 23171
rect 20729 23137 20763 23171
rect 21005 23137 21039 23171
rect 21281 23137 21315 23171
rect 21741 23137 21775 23171
rect 21925 23137 21959 23171
rect 22109 23137 22143 23171
rect 23489 23137 23523 23171
rect 24041 23137 24075 23171
rect 24133 23137 24167 23171
rect 24225 23137 24259 23171
rect 24363 23137 24397 23171
rect 26617 23137 26651 23171
rect 26985 23137 27019 23171
rect 27629 23137 27663 23171
rect 27721 23137 27755 23171
rect 19257 23069 19291 23103
rect 24501 23069 24535 23103
rect 25881 23069 25915 23103
rect 27353 23069 27387 23103
rect 20729 23001 20763 23035
rect 23857 23001 23891 23035
rect 27997 23001 28031 23035
rect 28733 23001 28767 23035
rect 19441 22933 19475 22967
rect 19717 22933 19751 22967
rect 19993 22933 20027 22967
rect 21373 22933 21407 22967
rect 23397 22933 23431 22967
rect 26525 22933 26559 22967
rect 27077 22933 27111 22967
rect 27905 22933 27939 22967
rect 28181 22933 28215 22967
rect 16865 22729 16899 22763
rect 20729 22729 20763 22763
rect 21465 22729 21499 22763
rect 13369 22661 13403 22695
rect 17877 22593 17911 22627
rect 19349 22593 19383 22627
rect 23857 22593 23891 22627
rect 12633 22525 12667 22559
rect 13553 22525 13587 22559
rect 13829 22525 13863 22559
rect 14013 22525 14047 22559
rect 14105 22525 14139 22559
rect 14197 22525 14231 22559
rect 14565 22525 14599 22559
rect 14832 22525 14866 22559
rect 16221 22525 16255 22559
rect 16405 22525 16439 22559
rect 16497 22525 16531 22559
rect 16589 22525 16623 22559
rect 17141 22525 17175 22559
rect 18153 22525 18187 22559
rect 18337 22525 18371 22559
rect 18705 22525 18739 22559
rect 18889 22525 18923 22559
rect 19616 22525 19650 22559
rect 20821 22525 20855 22559
rect 21097 22525 21131 22559
rect 21189 22525 21223 22559
rect 21281 22525 21315 22559
rect 21741 22525 21775 22559
rect 21833 22525 21867 22559
rect 21925 22525 21959 22559
rect 22043 22525 22077 22559
rect 22201 22525 22235 22559
rect 22937 22525 22971 22559
rect 24409 22525 24443 22559
rect 24593 22525 24627 22559
rect 24777 22525 24811 22559
rect 27261 22525 27295 22559
rect 27354 22525 27388 22559
rect 27491 22525 27525 22559
rect 27626 22525 27660 22559
rect 27726 22525 27760 22559
rect 28733 22525 28767 22559
rect 13001 22457 13035 22491
rect 13185 22457 13219 22491
rect 20959 22457 20993 22491
rect 23489 22457 23523 22491
rect 12725 22389 12759 22423
rect 13645 22389 13679 22423
rect 14473 22389 14507 22423
rect 15945 22389 15979 22423
rect 18245 22389 18279 22423
rect 18981 22389 19015 22423
rect 21557 22389 21591 22423
rect 23397 22389 23431 22423
rect 24685 22389 24719 22423
rect 27905 22389 27939 22423
rect 28641 22389 28675 22423
rect 12541 22185 12575 22219
rect 20177 22185 20211 22219
rect 25145 22185 25179 22219
rect 25329 22185 25363 22219
rect 14280 22117 14314 22151
rect 15485 22117 15519 22151
rect 18613 22117 18647 22151
rect 20545 22117 20579 22151
rect 21548 22117 21582 22151
rect 23366 22117 23400 22151
rect 25973 22117 26007 22151
rect 26433 22117 26467 22151
rect 27813 22117 27847 22151
rect 28043 22083 28077 22117
rect 13654 22049 13688 22083
rect 13921 22049 13955 22083
rect 14013 22049 14047 22083
rect 15669 22049 15703 22083
rect 16129 22049 16163 22083
rect 16681 22049 16715 22083
rect 17325 22049 17359 22083
rect 17417 22049 17451 22083
rect 17509 22049 17543 22083
rect 17693 22049 17727 22083
rect 17969 22049 18003 22083
rect 18153 22049 18187 22083
rect 18429 22049 18463 22083
rect 18797 22049 18831 22083
rect 19064 22049 19098 22083
rect 20453 22049 20487 22083
rect 20637 22049 20671 22083
rect 20755 22049 20789 22083
rect 23121 22049 23155 22083
rect 25237 22049 25271 22083
rect 26065 22049 26099 22083
rect 26249 22049 26283 22083
rect 26801 22049 26835 22083
rect 26893 22049 26927 22083
rect 27353 22049 27387 22083
rect 27629 22049 27663 22083
rect 28457 22049 28491 22083
rect 28724 22049 28758 22083
rect 15853 21981 15887 22015
rect 18245 21981 18279 22015
rect 20913 21981 20947 22015
rect 21281 21981 21315 22015
rect 24685 21981 24719 22015
rect 26525 21981 26559 22015
rect 27445 21981 27479 22015
rect 17877 21913 17911 21947
rect 22661 21913 22695 21947
rect 25053 21913 25087 21947
rect 25513 21913 25547 21947
rect 26065 21913 26099 21947
rect 27077 21913 27111 21947
rect 15393 21845 15427 21879
rect 17049 21845 17083 21879
rect 20269 21845 20303 21879
rect 24501 21845 24535 21879
rect 25605 21845 25639 21879
rect 25697 21845 25731 21879
rect 27169 21845 27203 21879
rect 27353 21845 27387 21879
rect 27997 21845 28031 21879
rect 28181 21845 28215 21879
rect 29837 21845 29871 21879
rect 13553 21641 13587 21675
rect 14749 21641 14783 21675
rect 19441 21641 19475 21675
rect 20453 21641 20487 21675
rect 21465 21641 21499 21675
rect 23213 21641 23247 21675
rect 24501 21641 24535 21675
rect 26341 21641 26375 21675
rect 28733 21641 28767 21675
rect 23121 21573 23155 21607
rect 26433 21573 26467 21607
rect 27997 21573 28031 21607
rect 23581 21505 23615 21539
rect 23857 21505 23891 21539
rect 24593 21505 24627 21539
rect 25697 21505 25731 21539
rect 25789 21505 25823 21539
rect 26249 21505 26283 21539
rect 27261 21505 27295 21539
rect 13829 21437 13863 21471
rect 13921 21437 13955 21471
rect 14013 21437 14047 21471
rect 14197 21437 14231 21471
rect 14841 21437 14875 21471
rect 16405 21437 16439 21471
rect 16589 21437 16623 21471
rect 16681 21437 16715 21471
rect 16865 21437 16899 21471
rect 17132 21437 17166 21471
rect 19257 21437 19291 21471
rect 19625 21437 19659 21471
rect 19809 21437 19843 21471
rect 20269 21437 20303 21471
rect 21557 21437 21591 21471
rect 21741 21437 21775 21471
rect 22008 21437 22042 21471
rect 23397 21437 23431 21471
rect 24869 21437 24903 21471
rect 24961 21437 24995 21471
rect 25053 21437 25087 21471
rect 25421 21437 25455 21471
rect 25605 21437 25639 21471
rect 25973 21437 26007 21471
rect 26525 21437 26559 21471
rect 27169 21437 27203 21471
rect 27445 21437 27479 21471
rect 27813 21437 27847 21471
rect 28089 21437 28123 21471
rect 28273 21437 28307 21471
rect 28365 21437 28399 21471
rect 28457 21437 28491 21471
rect 29009 21437 29043 21471
rect 19993 21369 20027 21403
rect 24731 21369 24765 21403
rect 27629 21369 27663 21403
rect 16313 21301 16347 21335
rect 18245 21301 18279 21335
rect 18705 21301 18739 21335
rect 20085 21301 20119 21335
rect 25237 21301 25271 21335
rect 26157 21301 26191 21335
rect 27721 21301 27755 21335
rect 29101 21301 29135 21335
rect 17601 21097 17635 21131
rect 21925 21097 21959 21131
rect 25145 21097 25179 21131
rect 27721 21097 27755 21131
rect 27997 21097 28031 21131
rect 30205 21097 30239 21131
rect 15945 21029 15979 21063
rect 16374 21029 16408 21063
rect 17785 21029 17819 21063
rect 28733 21029 28767 21063
rect 29070 21029 29104 21063
rect 15301 20961 15335 20995
rect 15485 20961 15519 20995
rect 15577 20961 15611 20995
rect 15669 20961 15703 20995
rect 16129 20961 16163 20995
rect 17969 20961 18003 20995
rect 22017 20961 22051 20995
rect 24777 20961 24811 20995
rect 27445 20961 27479 20995
rect 27629 20961 27663 20995
rect 27813 20961 27847 20995
rect 28089 20961 28123 20995
rect 28273 20961 28307 20995
rect 28365 20961 28399 20995
rect 28457 20961 28491 20995
rect 28825 20961 28859 20995
rect 24869 20893 24903 20927
rect 17509 20757 17543 20791
rect 15853 20553 15887 20587
rect 25697 20553 25731 20587
rect 26157 20553 26191 20587
rect 28181 20553 28215 20587
rect 20361 20417 20395 20451
rect 22937 20417 22971 20451
rect 16037 20349 16071 20383
rect 17785 20349 17819 20383
rect 18429 20349 18463 20383
rect 19257 20349 19291 20383
rect 19625 20349 19659 20383
rect 19901 20349 19935 20383
rect 20085 20349 20119 20383
rect 22017 20349 22051 20383
rect 22477 20349 22511 20383
rect 22569 20349 22603 20383
rect 22661 20349 22695 20383
rect 22799 20349 22833 20383
rect 25053 20349 25087 20383
rect 25201 20349 25235 20383
rect 25329 20349 25363 20383
rect 25518 20349 25552 20383
rect 26065 20349 26099 20383
rect 28273 20349 28307 20383
rect 16221 20281 16255 20315
rect 17969 20281 18003 20315
rect 18705 20281 18739 20315
rect 19993 20281 20027 20315
rect 20223 20281 20257 20315
rect 25421 20281 25455 20315
rect 18153 20213 18187 20247
rect 18337 20213 18371 20247
rect 19533 20213 19567 20247
rect 19717 20213 19751 20247
rect 22109 20213 22143 20247
rect 22293 20213 22327 20247
rect 19073 20009 19107 20043
rect 19432 19941 19466 19975
rect 21557 19941 21591 19975
rect 23121 19941 23155 19975
rect 26157 19941 26191 19975
rect 14841 19873 14875 19907
rect 14933 19873 14967 19907
rect 15025 19873 15059 19907
rect 15209 19873 15243 19907
rect 17693 19873 17727 19907
rect 17960 19873 17994 19907
rect 19165 19873 19199 19907
rect 20821 19873 20855 19907
rect 21281 19873 21315 19907
rect 21465 19873 21499 19907
rect 21649 19873 21683 19907
rect 21767 19873 21801 19907
rect 21925 19873 21959 19907
rect 23857 19873 23891 19907
rect 24961 19873 24995 19907
rect 25789 19873 25823 19907
rect 25881 19873 25915 19907
rect 26433 19873 26467 19907
rect 26617 19873 26651 19907
rect 26801 19873 26835 19907
rect 26985 19873 27019 19907
rect 27629 19873 27663 19907
rect 21005 19805 21039 19839
rect 22293 19805 22327 19839
rect 23765 19805 23799 19839
rect 24225 19805 24259 19839
rect 24869 19805 24903 19839
rect 26249 19805 26283 19839
rect 26709 19805 26743 19839
rect 27537 19805 27571 19839
rect 20545 19737 20579 19771
rect 25329 19737 25363 19771
rect 14565 19669 14599 19703
rect 20637 19669 20671 19703
rect 25605 19669 25639 19703
rect 27169 19669 27203 19703
rect 27261 19669 27295 19703
rect 19257 19465 19291 19499
rect 21741 19465 21775 19499
rect 23213 19465 23247 19499
rect 26433 19465 26467 19499
rect 28273 19465 28307 19499
rect 25237 19397 25271 19431
rect 23305 19329 23339 19363
rect 26709 19329 26743 19363
rect 14105 19261 14139 19295
rect 14197 19261 14231 19295
rect 14381 19261 14415 19295
rect 14648 19261 14682 19295
rect 15853 19261 15887 19295
rect 16221 19261 16255 19295
rect 16773 19261 16807 19295
rect 16865 19261 16899 19295
rect 16957 19261 16991 19295
rect 17141 19261 17175 19295
rect 17233 19261 17267 19295
rect 17877 19261 17911 19295
rect 17969 19261 18003 19295
rect 18061 19261 18095 19295
rect 18245 19261 18279 19295
rect 19441 19261 19475 19295
rect 19625 19261 19659 19295
rect 20269 19261 20303 19295
rect 20361 19261 20395 19295
rect 21833 19261 21867 19295
rect 23489 19261 23523 19295
rect 23857 19261 23891 19295
rect 25329 19261 25363 19295
rect 26341 19261 26375 19295
rect 26985 19261 27019 19295
rect 27169 19261 27203 19295
rect 16037 19193 16071 19227
rect 20177 19193 20211 19227
rect 20628 19193 20662 19227
rect 22100 19193 22134 19227
rect 23673 19193 23707 19227
rect 24102 19193 24136 19227
rect 26065 19193 26099 19227
rect 26433 19193 26467 19227
rect 27077 19193 27111 19227
rect 28089 19193 28123 19227
rect 28289 19193 28323 19227
rect 15761 19125 15795 19159
rect 16497 19125 16531 19159
rect 17325 19125 17359 19159
rect 17601 19125 17635 19159
rect 26525 19125 26559 19159
rect 28457 19125 28491 19159
rect 21557 18921 21591 18955
rect 22109 18921 22143 18955
rect 23581 18921 23615 18955
rect 24409 18921 24443 18955
rect 25881 18921 25915 18955
rect 27813 18921 27847 18955
rect 16742 18853 16776 18887
rect 18061 18853 18095 18887
rect 23857 18853 23891 18887
rect 27445 18853 27479 18887
rect 28273 18853 28307 18887
rect 29377 18853 29411 18887
rect 29653 18853 29687 18887
rect 15577 18785 15611 18819
rect 15761 18785 15795 18819
rect 16497 18785 16531 18819
rect 19625 18785 19659 18819
rect 21465 18783 21499 18817
rect 21925 18785 21959 18819
rect 22385 18785 22419 18819
rect 23765 18785 23799 18819
rect 23949 18785 23983 18819
rect 24067 18785 24101 18819
rect 24501 18785 24535 18819
rect 25053 18785 25087 18819
rect 25973 18785 26007 18819
rect 26617 18785 26651 18819
rect 27169 18785 27203 18819
rect 27353 18785 27387 18819
rect 27721 18785 27755 18819
rect 27997 18785 28031 18819
rect 29009 18785 29043 18819
rect 29837 18785 29871 18819
rect 18889 18717 18923 18751
rect 21741 18717 21775 18751
rect 24225 18717 24259 18751
rect 26525 18717 26559 18751
rect 26985 18717 27019 18751
rect 27445 18717 27479 18751
rect 27629 18717 27663 18751
rect 28181 18717 28215 18751
rect 28825 18717 28859 18751
rect 30021 18649 30055 18683
rect 15945 18581 15979 18615
rect 17877 18581 17911 18615
rect 19533 18581 19567 18615
rect 27353 18581 27387 18615
rect 29377 18581 29411 18615
rect 29561 18581 29595 18615
rect 16773 18377 16807 18411
rect 30389 18377 30423 18411
rect 20821 18241 20855 18275
rect 14565 18173 14599 18207
rect 14657 18173 14691 18207
rect 15393 18173 15427 18207
rect 17785 18173 17819 18207
rect 18153 18173 18187 18207
rect 18245 18173 18279 18207
rect 18337 18173 18371 18207
rect 18521 18173 18555 18207
rect 18889 18173 18923 18207
rect 20361 18173 20395 18207
rect 27077 18173 27111 18207
rect 27169 18173 27203 18207
rect 27353 18173 27387 18207
rect 27609 18173 27643 18207
rect 29009 18173 29043 18207
rect 29276 18173 29310 18207
rect 15025 18105 15059 18139
rect 15209 18105 15243 18139
rect 15638 18105 15672 18139
rect 16957 18105 16991 18139
rect 20453 18105 20487 18139
rect 20545 18105 20579 18139
rect 20683 18105 20717 18139
rect 14841 18037 14875 18071
rect 17877 18037 17911 18071
rect 20177 18037 20211 18071
rect 28733 18037 28767 18071
rect 15209 17833 15243 17867
rect 17325 17833 17359 17867
rect 20729 17833 20763 17867
rect 29193 17833 29227 17867
rect 17509 17765 17543 17799
rect 21557 17765 21591 17799
rect 21649 17765 21683 17799
rect 22477 17765 22511 17799
rect 22569 17765 22603 17799
rect 24777 17765 24811 17799
rect 14657 17697 14691 17731
rect 14749 17697 14783 17731
rect 14841 17697 14875 17731
rect 15025 17697 15059 17731
rect 16589 17697 16623 17731
rect 17693 17697 17727 17731
rect 18052 17697 18086 17731
rect 19349 17697 19383 17731
rect 19616 17697 19650 17731
rect 21465 17697 21499 17731
rect 21767 17697 21801 17731
rect 22201 17697 22235 17731
rect 22359 17697 22393 17731
rect 22661 17697 22695 17731
rect 23121 17697 23155 17731
rect 24501 17697 24535 17731
rect 24685 17697 24719 17731
rect 25237 17697 25271 17731
rect 25911 17697 25945 17731
rect 26065 17697 26099 17731
rect 29101 17697 29135 17731
rect 15761 17629 15795 17663
rect 17785 17629 17819 17663
rect 21925 17629 21959 17663
rect 23305 17629 23339 17663
rect 25145 17629 25179 17663
rect 25697 17561 25731 17595
rect 14381 17493 14415 17527
rect 19165 17493 19199 17527
rect 21281 17493 21315 17527
rect 22845 17493 22879 17527
rect 22937 17493 22971 17527
rect 24409 17493 24443 17527
rect 25605 17493 25639 17527
rect 15301 17289 15335 17323
rect 15393 17289 15427 17323
rect 17969 17289 18003 17323
rect 19441 17289 19475 17323
rect 21833 17289 21867 17323
rect 23581 17289 23615 17323
rect 26249 17289 26283 17323
rect 26985 17289 27019 17323
rect 17693 17221 17727 17255
rect 20269 17153 20303 17187
rect 20453 17153 20487 17187
rect 24501 17153 24535 17187
rect 24593 17153 24627 17187
rect 25881 17153 25915 17187
rect 13645 17085 13679 17119
rect 13737 17085 13771 17119
rect 13921 17085 13955 17119
rect 14188 17085 14222 17119
rect 15669 17085 15703 17119
rect 15761 17085 15795 17119
rect 15853 17085 15887 17119
rect 16037 17085 16071 17119
rect 17325 17085 17359 17119
rect 18061 17085 18095 17119
rect 19625 17085 19659 17119
rect 19809 17085 19843 17119
rect 20361 17085 20395 17119
rect 21925 17085 21959 17119
rect 22017 17085 22051 17119
rect 22201 17085 22235 17119
rect 22468 17085 22502 17119
rect 24041 17085 24075 17119
rect 24225 17085 24259 17119
rect 24363 17085 24397 17119
rect 24869 17085 24903 17119
rect 24961 17085 24995 17119
rect 25053 17085 25087 17119
rect 25513 17085 25547 17119
rect 25697 17085 25731 17119
rect 25789 17085 25823 17119
rect 26065 17085 26099 17119
rect 26341 17085 26375 17119
rect 26434 17085 26468 17119
rect 26806 17085 26840 17119
rect 27261 17085 27295 17119
rect 17509 17017 17543 17051
rect 20698 17017 20732 17051
rect 24134 17017 24168 17051
rect 24751 17017 24785 17051
rect 26617 17017 26651 17051
rect 26709 17017 26743 17051
rect 27169 17017 27203 17051
rect 23857 16949 23891 16983
rect 25237 16949 25271 16983
rect 17325 16745 17359 16779
rect 20545 16745 20579 16779
rect 23121 16745 23155 16779
rect 25605 16745 25639 16779
rect 17969 16677 18003 16711
rect 21557 16677 21591 16711
rect 21649 16677 21683 16711
rect 21787 16677 21821 16711
rect 22615 16677 22649 16711
rect 22845 16677 22879 16711
rect 15301 16609 15335 16643
rect 15455 16609 15489 16643
rect 16129 16609 16163 16643
rect 16405 16609 16439 16643
rect 16497 16609 16531 16643
rect 17141 16609 17175 16643
rect 17417 16609 17451 16643
rect 18521 16609 18555 16643
rect 18614 16609 18648 16643
rect 20729 16609 20763 16643
rect 21465 16609 21499 16643
rect 21925 16609 21959 16643
rect 22477 16609 22511 16643
rect 22753 16609 22787 16643
rect 22937 16609 22971 16643
rect 23581 16609 23615 16643
rect 23673 16609 23707 16643
rect 24225 16609 24259 16643
rect 24492 16609 24526 16643
rect 25697 16609 25731 16643
rect 25881 16609 25915 16643
rect 25973 16609 26007 16643
rect 26893 16609 26927 16643
rect 27261 16609 27295 16643
rect 27445 16609 27479 16643
rect 27537 16609 27571 16643
rect 27629 16609 27663 16643
rect 27997 16609 28031 16643
rect 20913 16541 20947 16575
rect 15669 16473 15703 16507
rect 18337 16473 18371 16507
rect 18889 16473 18923 16507
rect 16221 16405 16255 16439
rect 16681 16405 16715 16439
rect 16957 16405 16991 16439
rect 18429 16405 18463 16439
rect 21281 16405 21315 16439
rect 23857 16405 23891 16439
rect 26985 16405 27019 16439
rect 27905 16405 27939 16439
rect 28089 16405 28123 16439
rect 16773 16201 16807 16235
rect 17417 16201 17451 16235
rect 19349 16201 19383 16235
rect 19533 16201 19567 16235
rect 25237 16201 25271 16235
rect 27261 16201 27295 16235
rect 27077 16133 27111 16167
rect 17877 16065 17911 16099
rect 18429 16065 18463 16099
rect 20729 16065 20763 16099
rect 28825 16065 28859 16099
rect 29101 16065 29135 16099
rect 15393 15997 15427 16031
rect 15485 15997 15519 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 15946 15997 15980 16031
rect 16129 15997 16163 16031
rect 16359 15997 16393 16031
rect 16957 15997 16991 16031
rect 17049 15997 17083 16031
rect 17141 15997 17175 16031
rect 17325 15997 17359 16031
rect 17601 15997 17635 16031
rect 17693 15997 17727 16031
rect 17969 15997 18003 16031
rect 18061 15997 18095 16031
rect 18154 15997 18188 16031
rect 18705 15997 18739 16031
rect 18798 15997 18832 16031
rect 18981 15997 19015 16031
rect 19170 15997 19204 16031
rect 19441 15997 19475 16031
rect 19625 15997 19659 16031
rect 20913 15997 20947 16031
rect 21557 15997 21591 16031
rect 23489 15997 23523 16031
rect 23581 15997 23615 16031
rect 23857 15997 23891 16031
rect 24113 15997 24147 16031
rect 26709 15997 26743 16031
rect 27169 15997 27203 16031
rect 27353 15997 27387 16031
rect 28558 15997 28592 16031
rect 29009 15997 29043 16031
rect 15577 15929 15611 15963
rect 16221 15929 16255 15963
rect 19073 15929 19107 15963
rect 26893 15929 26927 15963
rect 15209 15861 15243 15895
rect 16497 15861 16531 15895
rect 21097 15861 21131 15895
rect 21465 15861 21499 15895
rect 26525 15861 26559 15895
rect 26801 15861 26835 15895
rect 27445 15861 27479 15895
rect 15669 15657 15703 15691
rect 16405 15657 16439 15691
rect 17785 15657 17819 15691
rect 22661 15657 22695 15691
rect 27261 15657 27295 15691
rect 15209 15589 15243 15623
rect 20269 15589 20303 15623
rect 21526 15589 21560 15623
rect 27077 15589 27111 15623
rect 28466 15589 28500 15623
rect 16497 15521 16531 15555
rect 17877 15521 17911 15555
rect 19441 15521 19475 15555
rect 19901 15521 19935 15555
rect 21281 15521 21315 15555
rect 26433 15521 26467 15555
rect 26617 15521 26651 15555
rect 28733 15521 28767 15555
rect 19533 15453 19567 15487
rect 20913 15453 20947 15487
rect 15485 15385 15519 15419
rect 19993 15385 20027 15419
rect 26709 15385 26743 15419
rect 27353 15385 27387 15419
rect 19717 15317 19751 15351
rect 26617 15317 26651 15351
rect 27077 15317 27111 15351
rect 16957 15113 16991 15147
rect 21005 15113 21039 15147
rect 23489 15113 23523 15147
rect 27077 15113 27111 15147
rect 27261 15113 27295 15147
rect 17877 15045 17911 15079
rect 16497 14977 16531 15011
rect 19257 14977 19291 15011
rect 19625 14977 19659 15011
rect 21649 14977 21683 15011
rect 14933 14909 14967 14943
rect 15945 14909 15979 14943
rect 16405 14909 16439 14943
rect 16681 14909 16715 14943
rect 16773 14909 16807 14943
rect 18061 14909 18095 14943
rect 18981 14909 19015 14943
rect 19073 14909 19107 14943
rect 19165 14909 19199 14943
rect 19881 14909 19915 14943
rect 21833 14909 21867 14943
rect 22109 14909 22143 14943
rect 24961 14909 24995 14943
rect 25145 14909 25179 14943
rect 25237 14909 25271 14943
rect 25329 14909 25363 14943
rect 25697 14909 25731 14943
rect 27169 14909 27203 14943
rect 27353 14909 27387 14943
rect 18153 14841 18187 14875
rect 22017 14841 22051 14875
rect 22354 14841 22388 14875
rect 25605 14841 25639 14875
rect 25942 14841 25976 14875
rect 14841 14773 14875 14807
rect 15853 14773 15887 14807
rect 18245 14773 18279 14807
rect 18429 14773 18463 14807
rect 18797 14773 18831 14807
rect 15101 14569 15135 14603
rect 16129 14569 16163 14603
rect 17325 14569 17359 14603
rect 17877 14569 17911 14603
rect 22293 14569 22327 14603
rect 25129 14569 25163 14603
rect 25881 14569 25915 14603
rect 26157 14569 26191 14603
rect 15301 14501 15335 14535
rect 18337 14501 18371 14535
rect 24685 14501 24719 14535
rect 25329 14501 25363 14535
rect 14473 14433 14507 14467
rect 15577 14433 15611 14467
rect 16865 14433 16899 14467
rect 17141 14433 17175 14467
rect 18061 14433 18095 14467
rect 19726 14433 19760 14467
rect 20269 14433 20303 14467
rect 22385 14433 22419 14467
rect 23949 14433 23983 14467
rect 24133 14433 24167 14467
rect 24317 14433 24351 14467
rect 25973 14433 26007 14467
rect 26249 14433 26283 14467
rect 14381 14365 14415 14399
rect 15485 14365 15519 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 18245 14365 18279 14399
rect 19993 14365 20027 14399
rect 20177 14365 20211 14399
rect 18613 14297 18647 14331
rect 24961 14297 24995 14331
rect 14197 14229 14231 14263
rect 14933 14229 14967 14263
rect 15117 14229 15151 14263
rect 15853 14229 15887 14263
rect 17049 14229 17083 14263
rect 18245 14229 18279 14263
rect 24041 14229 24075 14263
rect 24685 14229 24719 14263
rect 24869 14229 24903 14263
rect 25145 14229 25179 14263
rect 15301 14025 15335 14059
rect 17509 14025 17543 14059
rect 19165 14025 19199 14059
rect 23489 14025 23523 14059
rect 25329 14025 25363 14059
rect 18981 13957 19015 13991
rect 25237 13957 25271 13991
rect 15485 13889 15519 13923
rect 18153 13889 18187 13923
rect 18705 13889 18739 13923
rect 23121 13889 23155 13923
rect 23857 13889 23891 13923
rect 27445 13889 27479 13923
rect 13645 13821 13679 13855
rect 13737 13821 13771 13855
rect 13921 13821 13955 13855
rect 14177 13821 14211 13855
rect 16129 13821 16163 13855
rect 23213 13821 23247 13855
rect 25513 13821 25547 13855
rect 25789 13821 25823 13855
rect 26065 13821 26099 13855
rect 26709 13821 26743 13855
rect 16396 13753 16430 13787
rect 23305 13753 23339 13787
rect 23505 13753 23539 13787
rect 24102 13753 24136 13787
rect 25697 13753 25731 13787
rect 26893 13753 26927 13787
rect 16037 13685 16071 13719
rect 17601 13685 17635 13719
rect 23673 13685 23707 13719
rect 25973 13685 26007 13719
rect 26617 13685 26651 13719
rect 15761 13481 15795 13515
rect 16957 13481 16991 13515
rect 18429 13481 18463 13515
rect 23857 13481 23891 13515
rect 24317 13481 24351 13515
rect 27813 13481 27847 13515
rect 15945 13413 15979 13447
rect 24041 13413 24075 13447
rect 24225 13413 24259 13447
rect 25430 13413 25464 13447
rect 14197 13345 14231 13379
rect 14464 13345 14498 13379
rect 15669 13345 15703 13379
rect 17049 13345 17083 13379
rect 17877 13345 17911 13379
rect 18521 13345 18555 13379
rect 18981 13345 19015 13379
rect 25789 13345 25823 13379
rect 25973 13345 26007 13379
rect 26433 13345 26467 13379
rect 26689 13345 26723 13379
rect 16681 13277 16715 13311
rect 17969 13277 18003 13311
rect 19533 13277 19567 13311
rect 25697 13277 25731 13311
rect 15577 13209 15611 13243
rect 15945 13209 15979 13243
rect 18245 13209 18279 13243
rect 16129 13141 16163 13175
rect 25881 13141 25915 13175
rect 15117 12937 15151 12971
rect 16681 12937 16715 12971
rect 26249 12937 26283 12971
rect 18061 12869 18095 12903
rect 16497 12801 16531 12835
rect 17969 12801 18003 12835
rect 14933 12733 14967 12767
rect 15117 12733 15151 12767
rect 16313 12733 16347 12767
rect 16773 12733 16807 12767
rect 17049 12733 17083 12767
rect 17233 12733 17267 12767
rect 17325 12733 17359 12767
rect 18337 12733 18371 12767
rect 18889 12733 18923 12767
rect 25605 12733 25639 12767
rect 25789 12733 25823 12767
rect 25881 12733 25915 12767
rect 25973 12733 26007 12767
rect 18061 12665 18095 12699
rect 16129 12597 16163 12631
rect 17141 12597 17175 12631
rect 18245 12597 18279 12631
rect 18797 12597 18831 12631
rect 17049 12393 17083 12427
rect 17217 12393 17251 12427
rect 18153 12393 18187 12427
rect 17417 12325 17451 12359
rect 18512 12325 18546 12359
rect 15761 12257 15795 12291
rect 15945 12257 15979 12291
rect 16313 12257 16347 12291
rect 16865 12257 16899 12291
rect 17601 12257 17635 12291
rect 18245 12257 18279 12291
rect 15761 12053 15795 12087
rect 17233 12053 17267 12087
rect 19625 12053 19659 12087
rect 18245 11849 18279 11883
rect 14933 11645 14967 11679
rect 15025 11645 15059 11679
rect 15209 11645 15243 11679
rect 16865 11645 16899 11679
rect 17132 11645 17166 11679
rect 15476 11577 15510 11611
rect 16589 11509 16623 11543
rect 15669 11305 15703 11339
rect 17049 11305 17083 11339
rect 15577 11169 15611 11203
rect 15761 11169 15795 11203
rect 17141 11169 17175 11203
<< metal1 >>
rect 552 44634 31648 44656
rect 552 44582 3662 44634
rect 3714 44582 3726 44634
rect 3778 44582 3790 44634
rect 3842 44582 3854 44634
rect 3906 44582 3918 44634
rect 3970 44582 11436 44634
rect 11488 44582 11500 44634
rect 11552 44582 11564 44634
rect 11616 44582 11628 44634
rect 11680 44582 11692 44634
rect 11744 44582 19210 44634
rect 19262 44582 19274 44634
rect 19326 44582 19338 44634
rect 19390 44582 19402 44634
rect 19454 44582 19466 44634
rect 19518 44582 26984 44634
rect 27036 44582 27048 44634
rect 27100 44582 27112 44634
rect 27164 44582 27176 44634
rect 27228 44582 27240 44634
rect 27292 44582 31648 44634
rect 552 44560 31648 44582
rect 7190 44480 7196 44532
rect 7248 44480 7254 44532
rect 7650 44480 7656 44532
rect 7708 44480 7714 44532
rect 7929 44523 7987 44529
rect 7929 44489 7941 44523
rect 7975 44520 7987 44523
rect 8294 44520 8300 44532
rect 7975 44492 8300 44520
rect 7975 44489 7987 44492
rect 7929 44483 7987 44489
rect 8294 44480 8300 44492
rect 8352 44480 8358 44532
rect 8754 44480 8760 44532
rect 8812 44480 8818 44532
rect 9306 44480 9312 44532
rect 9364 44480 9370 44532
rect 11701 44523 11759 44529
rect 11701 44489 11713 44523
rect 11747 44520 11759 44523
rect 11790 44520 11796 44532
rect 11747 44492 11796 44520
rect 11747 44489 11759 44492
rect 11701 44483 11759 44489
rect 11790 44480 11796 44492
rect 11848 44480 11854 44532
rect 12802 44480 12808 44532
rect 12860 44480 12866 44532
rect 13078 44480 13084 44532
rect 13136 44480 13142 44532
rect 27430 44480 27436 44532
rect 27488 44520 27494 44532
rect 27488 44492 27936 44520
rect 27488 44480 27494 44492
rect 25222 44412 25228 44464
rect 25280 44452 25286 44464
rect 26421 44455 26479 44461
rect 26421 44452 26433 44455
rect 25280 44424 26433 44452
rect 25280 44412 25286 44424
rect 26421 44421 26433 44424
rect 26467 44421 26479 44455
rect 26421 44415 26479 44421
rect 11882 44344 11888 44396
rect 11940 44384 11946 44396
rect 26510 44384 26516 44396
rect 11940 44356 14136 44384
rect 11940 44344 11946 44356
rect 8021 44319 8079 44325
rect 8021 44285 8033 44319
rect 8067 44285 8079 44319
rect 8021 44279 8079 44285
rect 8036 44248 8064 44279
rect 8202 44276 8208 44328
rect 8260 44316 8266 44328
rect 8573 44319 8631 44325
rect 8573 44316 8585 44319
rect 8260 44288 8585 44316
rect 8260 44276 8266 44288
rect 8573 44285 8585 44288
rect 8619 44316 8631 44319
rect 9125 44319 9183 44325
rect 9125 44316 9137 44319
rect 8619 44288 9137 44316
rect 8619 44285 8631 44288
rect 8573 44279 8631 44285
rect 9125 44285 9137 44288
rect 9171 44285 9183 44319
rect 12345 44319 12403 44325
rect 12345 44316 12357 44319
rect 9125 44279 9183 44285
rect 11072 44288 12357 44316
rect 11072 44260 11100 44288
rect 12345 44285 12357 44288
rect 12391 44316 12403 44319
rect 12437 44319 12495 44325
rect 12437 44316 12449 44319
rect 12391 44288 12449 44316
rect 12391 44285 12403 44288
rect 12345 44279 12403 44285
rect 12437 44285 12449 44288
rect 12483 44285 12495 44319
rect 12437 44279 12495 44285
rect 11054 44248 11060 44260
rect 8036 44220 11060 44248
rect 11054 44208 11060 44220
rect 11112 44208 11118 44260
rect 12452 44248 12480 44279
rect 13722 44276 13728 44328
rect 13780 44276 13786 44328
rect 13814 44276 13820 44328
rect 13872 44276 13878 44328
rect 13998 44276 14004 44328
rect 14056 44276 14062 44328
rect 14108 44325 14136 44356
rect 25792 44356 26516 44384
rect 14093 44319 14151 44325
rect 14093 44285 14105 44319
rect 14139 44285 14151 44319
rect 14093 44279 14151 44285
rect 14553 44319 14611 44325
rect 14553 44285 14565 44319
rect 14599 44285 14611 44319
rect 14553 44279 14611 44285
rect 15197 44319 15255 44325
rect 15197 44285 15209 44319
rect 15243 44316 15255 44319
rect 15838 44316 15844 44328
rect 15243 44288 15844 44316
rect 15243 44285 15255 44288
rect 15197 44279 15255 44285
rect 14568 44248 14596 44279
rect 15838 44276 15844 44288
rect 15896 44276 15902 44328
rect 16482 44276 16488 44328
rect 16540 44316 16546 44328
rect 17037 44319 17095 44325
rect 17037 44316 17049 44319
rect 16540 44288 17049 44316
rect 16540 44276 16546 44288
rect 17037 44285 17049 44288
rect 17083 44316 17095 44319
rect 19337 44319 19395 44325
rect 19337 44316 19349 44319
rect 17083 44288 19349 44316
rect 17083 44285 17095 44288
rect 17037 44279 17095 44285
rect 19337 44285 19349 44288
rect 19383 44285 19395 44319
rect 19337 44279 19395 44285
rect 21634 44276 21640 44328
rect 21692 44276 21698 44328
rect 24026 44276 24032 44328
rect 24084 44276 24090 44328
rect 24394 44276 24400 44328
rect 24452 44276 24458 44328
rect 24946 44276 24952 44328
rect 25004 44276 25010 44328
rect 25498 44276 25504 44328
rect 25556 44276 25562 44328
rect 25792 44325 25820 44356
rect 26510 44344 26516 44356
rect 26568 44344 26574 44396
rect 25777 44319 25835 44325
rect 25777 44285 25789 44319
rect 25823 44285 25835 44319
rect 25777 44279 25835 44285
rect 26050 44276 26056 44328
rect 26108 44276 26114 44328
rect 27908 44325 27936 44492
rect 28994 44344 29000 44396
rect 29052 44344 29058 44396
rect 27801 44319 27859 44325
rect 27801 44316 27813 44319
rect 27448 44288 27813 44316
rect 27448 44260 27476 44288
rect 27801 44285 27813 44288
rect 27847 44285 27859 44319
rect 27801 44279 27859 44285
rect 27893 44319 27951 44325
rect 27893 44285 27905 44319
rect 27939 44285 27951 44319
rect 27893 44279 27951 44285
rect 28166 44276 28172 44328
rect 28224 44276 28230 44328
rect 29270 44276 29276 44328
rect 29328 44276 29334 44328
rect 12452 44220 14596 44248
rect 25976 44220 26924 44248
rect 8113 44183 8171 44189
rect 8113 44149 8125 44183
rect 8159 44180 8171 44183
rect 8294 44180 8300 44192
rect 8159 44152 8300 44180
rect 8159 44149 8171 44152
rect 8113 44143 8171 44149
rect 8294 44140 8300 44152
rect 8352 44140 8358 44192
rect 12253 44183 12311 44189
rect 12253 44149 12265 44183
rect 12299 44180 12311 44183
rect 12434 44180 12440 44192
rect 12299 44152 12440 44180
rect 12299 44149 12311 44152
rect 12253 44143 12311 44149
rect 12434 44140 12440 44152
rect 12492 44140 12498 44192
rect 12526 44140 12532 44192
rect 12584 44140 12590 44192
rect 13538 44140 13544 44192
rect 13596 44140 13602 44192
rect 14274 44140 14280 44192
rect 14332 44180 14338 44192
rect 14461 44183 14519 44189
rect 14461 44180 14473 44183
rect 14332 44152 14473 44180
rect 14332 44140 14338 44152
rect 14461 44149 14473 44152
rect 14507 44149 14519 44183
rect 14461 44143 14519 44149
rect 15013 44183 15071 44189
rect 15013 44149 15025 44183
rect 15059 44180 15071 44183
rect 15746 44180 15752 44192
rect 15059 44152 15752 44180
rect 15059 44149 15071 44152
rect 15013 44143 15071 44149
rect 15746 44140 15752 44152
rect 15804 44140 15810 44192
rect 16758 44140 16764 44192
rect 16816 44180 16822 44192
rect 16945 44183 17003 44189
rect 16945 44180 16957 44183
rect 16816 44152 16957 44180
rect 16816 44140 16822 44152
rect 16945 44149 16957 44152
rect 16991 44149 17003 44183
rect 16945 44143 17003 44149
rect 19242 44140 19248 44192
rect 19300 44180 19306 44192
rect 19429 44183 19487 44189
rect 19429 44180 19441 44183
rect 19300 44152 19441 44180
rect 19300 44140 19306 44152
rect 19429 44149 19441 44152
rect 19475 44149 19487 44183
rect 19429 44143 19487 44149
rect 21818 44140 21824 44192
rect 21876 44140 21882 44192
rect 22002 44140 22008 44192
rect 22060 44180 22066 44192
rect 23845 44183 23903 44189
rect 23845 44180 23857 44183
rect 22060 44152 23857 44180
rect 22060 44140 22066 44152
rect 23845 44149 23857 44152
rect 23891 44149 23903 44183
rect 23845 44143 23903 44149
rect 24578 44140 24584 44192
rect 24636 44140 24642 44192
rect 25130 44140 25136 44192
rect 25188 44140 25194 44192
rect 25682 44140 25688 44192
rect 25740 44140 25746 44192
rect 25976 44189 26004 44220
rect 25961 44183 26019 44189
rect 25961 44149 25973 44183
rect 26007 44149 26019 44183
rect 25961 44143 26019 44149
rect 26234 44140 26240 44192
rect 26292 44140 26298 44192
rect 26896 44180 26924 44220
rect 27430 44208 27436 44260
rect 27488 44208 27494 44260
rect 27534 44251 27592 44257
rect 27534 44217 27546 44251
rect 27580 44217 27592 44251
rect 27534 44211 27592 44217
rect 27540 44180 27568 44211
rect 26896 44152 27568 44180
rect 28074 44140 28080 44192
rect 28132 44140 28138 44192
rect 28353 44183 28411 44189
rect 28353 44149 28365 44183
rect 28399 44180 28411 44183
rect 28994 44180 29000 44192
rect 28399 44152 29000 44180
rect 28399 44149 28411 44152
rect 28353 44143 28411 44149
rect 28994 44140 29000 44152
rect 29052 44140 29058 44192
rect 552 44090 31648 44112
rect 552 44038 4322 44090
rect 4374 44038 4386 44090
rect 4438 44038 4450 44090
rect 4502 44038 4514 44090
rect 4566 44038 4578 44090
rect 4630 44038 12096 44090
rect 12148 44038 12160 44090
rect 12212 44038 12224 44090
rect 12276 44038 12288 44090
rect 12340 44038 12352 44090
rect 12404 44038 19870 44090
rect 19922 44038 19934 44090
rect 19986 44038 19998 44090
rect 20050 44038 20062 44090
rect 20114 44038 20126 44090
rect 20178 44038 27644 44090
rect 27696 44038 27708 44090
rect 27760 44038 27772 44090
rect 27824 44038 27836 44090
rect 27888 44038 27900 44090
rect 27952 44038 31648 44090
rect 552 44016 31648 44038
rect 6546 43936 6552 43988
rect 6604 43936 6610 43988
rect 6914 43936 6920 43988
rect 6972 43936 6978 43988
rect 8202 43936 8208 43988
rect 8260 43976 8266 43988
rect 9677 43979 9735 43985
rect 9677 43976 9689 43979
rect 8260 43948 9689 43976
rect 8260 43936 8266 43948
rect 9677 43945 9689 43948
rect 9723 43945 9735 43979
rect 9677 43939 9735 43945
rect 6733 43843 6791 43849
rect 6733 43809 6745 43843
rect 6779 43840 6791 43843
rect 7101 43843 7159 43849
rect 7101 43840 7113 43843
rect 6779 43812 7113 43840
rect 6779 43809 6791 43812
rect 6733 43803 6791 43809
rect 7101 43809 7113 43812
rect 7147 43840 7159 43843
rect 8202 43840 8208 43852
rect 7147 43812 8208 43840
rect 7147 43809 7159 43812
rect 7101 43803 7159 43809
rect 8202 43800 8208 43812
rect 8260 43800 8266 43852
rect 8294 43800 8300 43852
rect 8352 43800 8358 43852
rect 8564 43843 8622 43849
rect 8564 43809 8576 43843
rect 8610 43840 8622 43843
rect 8846 43840 8852 43852
rect 8610 43812 8852 43840
rect 8610 43809 8622 43812
rect 8564 43803 8622 43809
rect 8846 43800 8852 43812
rect 8904 43800 8910 43852
rect 9692 43840 9720 43939
rect 10686 43936 10692 43988
rect 10744 43936 10750 43988
rect 13262 43936 13268 43988
rect 13320 43936 13326 43988
rect 13541 43979 13599 43985
rect 13541 43945 13553 43979
rect 13587 43976 13599 43979
rect 13814 43976 13820 43988
rect 13587 43948 13820 43976
rect 13587 43945 13599 43948
rect 13541 43939 13599 43945
rect 13814 43936 13820 43948
rect 13872 43936 13878 43988
rect 18138 43936 18144 43988
rect 18196 43936 18202 43988
rect 26421 43979 26479 43985
rect 26421 43976 26433 43979
rect 23216 43948 26433 43976
rect 15933 43911 15991 43917
rect 15933 43877 15945 43911
rect 15979 43908 15991 43911
rect 16574 43908 16580 43920
rect 15979 43880 16580 43908
rect 15979 43877 15991 43880
rect 15933 43871 15991 43877
rect 16574 43868 16580 43880
rect 16632 43868 16638 43920
rect 21818 43868 21824 43920
rect 21876 43908 21882 43920
rect 23216 43917 23244 43948
rect 26421 43945 26433 43948
rect 26467 43945 26479 43979
rect 27893 43979 27951 43985
rect 27893 43976 27905 43979
rect 26421 43939 26479 43945
rect 27632 43948 27905 43976
rect 22382 43911 22440 43917
rect 22382 43908 22394 43911
rect 21876 43880 22394 43908
rect 21876 43868 21882 43880
rect 22382 43877 22394 43880
rect 22428 43877 22440 43911
rect 22382 43871 22440 43877
rect 23201 43911 23259 43917
rect 23201 43877 23213 43911
rect 23247 43877 23259 43911
rect 23201 43871 23259 43877
rect 25130 43868 25136 43920
rect 25188 43917 25194 43920
rect 25188 43908 25200 43917
rect 25188 43880 25233 43908
rect 25188 43871 25200 43880
rect 25188 43868 25194 43871
rect 26234 43868 26240 43920
rect 26292 43908 26298 43920
rect 27534 43911 27592 43917
rect 27534 43908 27546 43911
rect 26292 43880 27546 43908
rect 26292 43868 26298 43880
rect 27534 43877 27546 43880
rect 27580 43877 27592 43911
rect 27534 43871 27592 43877
rect 10321 43843 10379 43849
rect 10321 43840 10333 43843
rect 9692 43812 10333 43840
rect 10321 43809 10333 43812
rect 10367 43840 10379 43843
rect 10505 43843 10563 43849
rect 10505 43840 10517 43843
rect 10367 43812 10517 43840
rect 10367 43809 10379 43812
rect 10321 43803 10379 43809
rect 10505 43809 10517 43812
rect 10551 43809 10563 43843
rect 10505 43803 10563 43809
rect 11238 43800 11244 43852
rect 11296 43840 11302 43852
rect 12078 43843 12136 43849
rect 12078 43840 12090 43843
rect 11296 43812 12090 43840
rect 11296 43800 11302 43812
rect 12078 43809 12090 43812
rect 12124 43809 12136 43843
rect 12078 43803 12136 43809
rect 12342 43800 12348 43852
rect 12400 43800 12406 43852
rect 12805 43843 12863 43849
rect 12805 43809 12817 43843
rect 12851 43809 12863 43843
rect 12805 43803 12863 43809
rect 13357 43843 13415 43849
rect 13357 43809 13369 43843
rect 13403 43840 13415 43843
rect 13998 43840 14004 43852
rect 13403 43812 14004 43840
rect 13403 43809 13415 43812
rect 13357 43803 13415 43809
rect 12820 43772 12848 43803
rect 13998 43800 14004 43812
rect 14056 43800 14062 43852
rect 14274 43800 14280 43852
rect 14332 43800 14338 43852
rect 16114 43800 16120 43852
rect 16172 43840 16178 43852
rect 16301 43843 16359 43849
rect 16301 43840 16313 43843
rect 16172 43812 16313 43840
rect 16172 43800 16178 43812
rect 16301 43809 16313 43812
rect 16347 43809 16359 43843
rect 16301 43803 16359 43809
rect 16758 43800 16764 43852
rect 16816 43800 16822 43852
rect 19242 43800 19248 43852
rect 19300 43800 19306 43852
rect 22922 43800 22928 43852
rect 22980 43840 22986 43852
rect 23109 43843 23167 43849
rect 23109 43840 23121 43843
rect 22980 43812 23121 43840
rect 22980 43800 22986 43812
rect 23109 43809 23121 43812
rect 23155 43809 23167 43843
rect 23109 43803 23167 43809
rect 23293 43843 23351 43849
rect 23293 43809 23305 43843
rect 23339 43840 23351 43843
rect 23382 43840 23388 43852
rect 23339 43812 23388 43840
rect 23339 43809 23351 43812
rect 23293 43803 23351 43809
rect 23382 43800 23388 43812
rect 23440 43800 23446 43852
rect 23477 43843 23535 43849
rect 23477 43809 23489 43843
rect 23523 43840 23535 43843
rect 27632 43840 27660 43948
rect 27893 43945 27905 43948
rect 27939 43945 27951 43979
rect 27893 43939 27951 43945
rect 23523 43812 27660 43840
rect 23523 43809 23535 43812
rect 23477 43803 23535 43809
rect 28994 43800 29000 43852
rect 29052 43849 29058 43852
rect 29052 43840 29064 43849
rect 29273 43843 29331 43849
rect 29052 43812 29097 43840
rect 29052 43803 29064 43812
rect 29273 43809 29285 43843
rect 29319 43809 29331 43843
rect 29273 43803 29331 43809
rect 29052 43800 29058 43803
rect 14182 43772 14188 43784
rect 12820 43744 14188 43772
rect 14182 43732 14188 43744
rect 14240 43732 14246 43784
rect 14553 43775 14611 43781
rect 14553 43741 14565 43775
rect 14599 43772 14611 43775
rect 15286 43772 15292 43784
rect 14599 43744 15292 43772
rect 14599 43741 14611 43744
rect 14553 43735 14611 43741
rect 15286 43732 15292 43744
rect 15344 43732 15350 43784
rect 17034 43732 17040 43784
rect 17092 43732 17098 43784
rect 19521 43775 19579 43781
rect 19521 43741 19533 43775
rect 19567 43772 19579 43775
rect 19702 43772 19708 43784
rect 19567 43744 19708 43772
rect 19567 43741 19579 43744
rect 19521 43735 19579 43741
rect 19702 43732 19708 43744
rect 19760 43732 19766 43784
rect 22649 43775 22707 43781
rect 22649 43741 22661 43775
rect 22695 43741 22707 43775
rect 22649 43735 22707 43741
rect 15838 43664 15844 43716
rect 15896 43704 15902 43716
rect 16117 43707 16175 43713
rect 16117 43704 16129 43707
rect 15896 43676 16129 43704
rect 15896 43664 15902 43676
rect 16117 43673 16129 43676
rect 16163 43673 16175 43707
rect 16117 43667 16175 43673
rect 9766 43596 9772 43648
rect 9824 43596 9830 43648
rect 10962 43596 10968 43648
rect 11020 43596 11026 43648
rect 12713 43639 12771 43645
rect 12713 43605 12725 43639
rect 12759 43636 12771 43639
rect 13814 43636 13820 43648
rect 12759 43608 13820 43636
rect 12759 43605 12771 43608
rect 12713 43599 12771 43605
rect 13814 43596 13820 43608
rect 13872 43596 13878 43648
rect 19610 43596 19616 43648
rect 19668 43636 19674 43648
rect 20625 43639 20683 43645
rect 20625 43636 20637 43639
rect 19668 43608 20637 43636
rect 19668 43596 19674 43608
rect 20625 43605 20637 43608
rect 20671 43605 20683 43639
rect 20625 43599 20683 43605
rect 21269 43639 21327 43645
rect 21269 43605 21281 43639
rect 21315 43636 21327 43639
rect 21450 43636 21456 43648
rect 21315 43608 21456 43636
rect 21315 43605 21327 43608
rect 21269 43599 21327 43605
rect 21450 43596 21456 43608
rect 21508 43596 21514 43648
rect 22370 43596 22376 43648
rect 22428 43636 22434 43648
rect 22664 43636 22692 43735
rect 25406 43732 25412 43784
rect 25464 43732 25470 43784
rect 27801 43775 27859 43781
rect 27801 43741 27813 43775
rect 27847 43741 27859 43775
rect 27801 43735 27859 43741
rect 22428 43608 22692 43636
rect 22925 43639 22983 43645
rect 22428 43596 22434 43608
rect 22925 43605 22937 43639
rect 22971 43636 22983 43639
rect 23198 43636 23204 43648
rect 22971 43608 23204 43636
rect 22971 43605 22983 43608
rect 22925 43599 22983 43605
rect 23198 43596 23204 43608
rect 23256 43596 23262 43648
rect 24029 43639 24087 43645
rect 24029 43605 24041 43639
rect 24075 43636 24087 43639
rect 24394 43636 24400 43648
rect 24075 43608 24400 43636
rect 24075 43605 24087 43608
rect 24029 43599 24087 43605
rect 24394 43596 24400 43608
rect 24452 43596 24458 43648
rect 27522 43596 27528 43648
rect 27580 43636 27586 43648
rect 27816 43636 27844 43735
rect 29288 43636 29316 43803
rect 27580 43608 29316 43636
rect 27580 43596 27586 43608
rect 552 43546 31648 43568
rect 552 43494 3662 43546
rect 3714 43494 3726 43546
rect 3778 43494 3790 43546
rect 3842 43494 3854 43546
rect 3906 43494 3918 43546
rect 3970 43494 11436 43546
rect 11488 43494 11500 43546
rect 11552 43494 11564 43546
rect 11616 43494 11628 43546
rect 11680 43494 11692 43546
rect 11744 43494 19210 43546
rect 19262 43494 19274 43546
rect 19326 43494 19338 43546
rect 19390 43494 19402 43546
rect 19454 43494 19466 43546
rect 19518 43494 26984 43546
rect 27036 43494 27048 43546
rect 27100 43494 27112 43546
rect 27164 43494 27176 43546
rect 27228 43494 27240 43546
rect 27292 43494 31648 43546
rect 552 43472 31648 43494
rect 8846 43392 8852 43444
rect 8904 43392 8910 43444
rect 11330 43392 11336 43444
rect 11388 43432 11394 43444
rect 11609 43435 11667 43441
rect 11609 43432 11621 43435
rect 11388 43404 11621 43432
rect 11388 43392 11394 43404
rect 11609 43401 11621 43404
rect 11655 43401 11667 43435
rect 11609 43395 11667 43401
rect 13633 43435 13691 43441
rect 13633 43401 13645 43435
rect 13679 43432 13691 43435
rect 14366 43432 14372 43444
rect 13679 43404 14372 43432
rect 13679 43401 13691 43404
rect 13633 43395 13691 43401
rect 14366 43392 14372 43404
rect 14424 43392 14430 43444
rect 15286 43392 15292 43444
rect 15344 43392 15350 43444
rect 23474 43432 23480 43444
rect 20088 43404 23480 43432
rect 9766 43324 9772 43376
rect 9824 43324 9830 43376
rect 13357 43367 13415 43373
rect 13357 43333 13369 43367
rect 13403 43364 13415 43367
rect 14182 43364 14188 43376
rect 13403 43336 14188 43364
rect 13403 43333 13415 43336
rect 13357 43327 13415 43333
rect 14182 43324 14188 43336
rect 14240 43324 14246 43376
rect 17126 43324 17132 43376
rect 17184 43364 17190 43376
rect 20088 43364 20116 43404
rect 23474 43392 23480 43404
rect 23532 43392 23538 43444
rect 17184 43336 20116 43364
rect 17184 43324 17190 43336
rect 9784 43296 9812 43324
rect 15105 43299 15163 43305
rect 15105 43296 15117 43299
rect 9232 43268 9812 43296
rect 13832 43268 15117 43296
rect 9232 43237 9260 43268
rect 9217 43231 9275 43237
rect 9217 43197 9229 43231
rect 9263 43197 9275 43231
rect 9217 43191 9275 43197
rect 9398 43188 9404 43240
rect 9456 43228 9462 43240
rect 9585 43231 9643 43237
rect 9585 43228 9597 43231
rect 9456 43200 9597 43228
rect 9456 43188 9462 43200
rect 9585 43197 9597 43200
rect 9631 43197 9643 43231
rect 9585 43191 9643 43197
rect 9677 43231 9735 43237
rect 9677 43197 9689 43231
rect 9723 43197 9735 43231
rect 9677 43191 9735 43197
rect 9769 43231 9827 43237
rect 9769 43197 9781 43231
rect 9815 43228 9827 43231
rect 10318 43228 10324 43240
rect 9815 43200 10324 43228
rect 9815 43197 9827 43200
rect 9769 43191 9827 43197
rect 9033 43163 9091 43169
rect 9033 43129 9045 43163
rect 9079 43129 9091 43163
rect 9692 43160 9720 43191
rect 10318 43188 10324 43200
rect 10376 43188 10382 43240
rect 10962 43188 10968 43240
rect 11020 43228 11026 43240
rect 11425 43231 11483 43237
rect 11425 43228 11437 43231
rect 11020 43200 11437 43228
rect 11020 43188 11026 43200
rect 11425 43197 11437 43200
rect 11471 43197 11483 43231
rect 11425 43191 11483 43197
rect 11974 43188 11980 43240
rect 12032 43188 12038 43240
rect 12244 43231 12302 43237
rect 12244 43197 12256 43231
rect 12290 43228 12302 43231
rect 13538 43228 13544 43240
rect 12290 43200 13544 43228
rect 12290 43197 12302 43200
rect 12244 43191 12302 43197
rect 13538 43188 13544 43200
rect 13596 43188 13602 43240
rect 13832 43237 13860 43268
rect 15105 43265 15117 43268
rect 15151 43265 15163 43299
rect 15105 43259 15163 43265
rect 15580 43268 16436 43296
rect 13817 43231 13875 43237
rect 13817 43197 13829 43231
rect 13863 43197 13875 43231
rect 13817 43191 13875 43197
rect 13998 43188 14004 43240
rect 14056 43228 14062 43240
rect 14093 43231 14151 43237
rect 14093 43228 14105 43231
rect 14056 43200 14105 43228
rect 14056 43188 14062 43200
rect 14093 43197 14105 43200
rect 14139 43197 14151 43231
rect 14093 43191 14151 43197
rect 14182 43188 14188 43240
rect 14240 43228 14246 43240
rect 14829 43231 14887 43237
rect 14829 43228 14841 43231
rect 14240 43200 14841 43228
rect 14240 43188 14246 43200
rect 14829 43197 14841 43200
rect 14875 43197 14887 43231
rect 14829 43191 14887 43197
rect 15010 43188 15016 43240
rect 15068 43188 15074 43240
rect 15580 43237 15608 43268
rect 15565 43231 15623 43237
rect 15565 43197 15577 43231
rect 15611 43197 15623 43231
rect 15565 43191 15623 43197
rect 15654 43188 15660 43240
rect 15712 43188 15718 43240
rect 15749 43231 15807 43237
rect 15749 43197 15761 43231
rect 15795 43197 15807 43231
rect 15749 43191 15807 43197
rect 11054 43160 11060 43172
rect 9692 43132 11060 43160
rect 9033 43123 9091 43129
rect 9048 43092 9076 43123
rect 11054 43120 11060 43132
rect 11112 43120 11118 43172
rect 9861 43095 9919 43101
rect 9861 43092 9873 43095
rect 9048 43064 9873 43092
rect 9861 43061 9873 43064
rect 9907 43092 9919 43095
rect 11882 43092 11888 43104
rect 9907 43064 11888 43092
rect 9907 43061 9919 43064
rect 9861 43055 9919 43061
rect 11882 43052 11888 43064
rect 11940 43052 11946 43104
rect 14182 43052 14188 43104
rect 14240 43092 14246 43104
rect 14737 43095 14795 43101
rect 14737 43092 14749 43095
rect 14240 43064 14749 43092
rect 14240 43052 14246 43064
rect 14737 43061 14749 43064
rect 14783 43061 14795 43095
rect 14737 43055 14795 43061
rect 15562 43052 15568 43104
rect 15620 43092 15626 43104
rect 15764 43092 15792 43191
rect 15838 43188 15844 43240
rect 15896 43228 15902 43240
rect 15933 43231 15991 43237
rect 15933 43228 15945 43231
rect 15896 43200 15945 43228
rect 15896 43188 15902 43200
rect 15933 43197 15945 43200
rect 15979 43197 15991 43231
rect 15933 43191 15991 43197
rect 16022 43188 16028 43240
rect 16080 43188 16086 43240
rect 16298 43188 16304 43240
rect 16356 43188 16362 43240
rect 16408 43228 16436 43268
rect 16482 43256 16488 43308
rect 16540 43296 16546 43308
rect 18785 43299 18843 43305
rect 16540 43268 18736 43296
rect 16540 43256 16546 43268
rect 16574 43228 16580 43240
rect 16408 43200 16580 43228
rect 16574 43188 16580 43200
rect 16632 43228 16638 43240
rect 16761 43231 16819 43237
rect 16761 43228 16773 43231
rect 16632 43200 16773 43228
rect 16632 43188 16638 43200
rect 16761 43197 16773 43200
rect 16807 43197 16819 43231
rect 16761 43191 16819 43197
rect 17037 43231 17095 43237
rect 17037 43197 17049 43231
rect 17083 43228 17095 43231
rect 17126 43228 17132 43240
rect 17083 43200 17132 43228
rect 17083 43197 17095 43200
rect 17037 43191 17095 43197
rect 17126 43188 17132 43200
rect 17184 43188 17190 43240
rect 17402 43188 17408 43240
rect 17460 43188 17466 43240
rect 17494 43188 17500 43240
rect 17552 43228 17558 43240
rect 17681 43231 17739 43237
rect 17681 43228 17693 43231
rect 17552 43200 17693 43228
rect 17552 43188 17558 43200
rect 17681 43197 17693 43200
rect 17727 43197 17739 43231
rect 17681 43191 17739 43197
rect 17770 43188 17776 43240
rect 17828 43228 17834 43240
rect 18708 43237 18736 43268
rect 18785 43265 18797 43299
rect 18831 43296 18843 43299
rect 19518 43296 19524 43308
rect 18831 43268 19524 43296
rect 18831 43265 18843 43268
rect 18785 43259 18843 43265
rect 19518 43256 19524 43268
rect 19576 43256 19582 43308
rect 17911 43231 17969 43237
rect 17911 43228 17923 43231
rect 17828 43200 17923 43228
rect 17828 43188 17834 43200
rect 17911 43197 17923 43200
rect 17957 43197 17969 43231
rect 18269 43231 18327 43237
rect 18269 43228 18281 43231
rect 17911 43191 17969 43197
rect 18248 43197 18281 43228
rect 18315 43197 18327 43231
rect 18248 43191 18327 43197
rect 18417 43231 18475 43237
rect 18417 43197 18429 43231
rect 18463 43197 18475 43231
rect 18417 43191 18475 43197
rect 18693 43231 18751 43237
rect 18693 43197 18705 43231
rect 18739 43197 18751 43231
rect 18693 43191 18751 43197
rect 16117 43163 16175 43169
rect 16117 43129 16129 43163
rect 16163 43160 16175 43163
rect 16945 43163 17003 43169
rect 16945 43160 16957 43163
rect 16163 43132 16957 43160
rect 16163 43129 16175 43132
rect 16117 43123 16175 43129
rect 16776 43104 16804 43132
rect 16945 43129 16957 43132
rect 16991 43129 17003 43163
rect 17420 43160 17448 43188
rect 18049 43163 18107 43169
rect 18049 43160 18061 43163
rect 17420 43132 18061 43160
rect 16945 43123 17003 43129
rect 18049 43129 18061 43132
rect 18095 43129 18107 43163
rect 18049 43123 18107 43129
rect 18138 43120 18144 43172
rect 18196 43120 18202 43172
rect 15620 43064 15792 43092
rect 15620 43052 15626 43064
rect 16390 43052 16396 43104
rect 16448 43092 16454 43104
rect 16485 43095 16543 43101
rect 16485 43092 16497 43095
rect 16448 43064 16497 43092
rect 16448 43052 16454 43064
rect 16485 43061 16497 43064
rect 16531 43061 16543 43095
rect 16485 43055 16543 43061
rect 16574 43052 16580 43104
rect 16632 43052 16638 43104
rect 16758 43052 16764 43104
rect 16816 43052 16822 43104
rect 17218 43052 17224 43104
rect 17276 43052 17282 43104
rect 17586 43052 17592 43104
rect 17644 43052 17650 43104
rect 17770 43052 17776 43104
rect 17828 43052 17834 43104
rect 17954 43052 17960 43104
rect 18012 43092 18018 43104
rect 18248 43092 18276 43191
rect 18432 43160 18460 43191
rect 18874 43188 18880 43240
rect 18932 43228 18938 43240
rect 19245 43231 19303 43237
rect 19245 43228 19257 43231
rect 18932 43200 19257 43228
rect 18932 43188 18938 43200
rect 19245 43197 19257 43200
rect 19291 43197 19303 43231
rect 19245 43191 19303 43197
rect 19610 43188 19616 43240
rect 19668 43188 19674 43240
rect 19705 43231 19763 43237
rect 19705 43197 19717 43231
rect 19751 43228 19763 43231
rect 19794 43228 19800 43240
rect 19751 43200 19800 43228
rect 19751 43197 19763 43200
rect 19705 43191 19763 43197
rect 19794 43188 19800 43200
rect 19852 43188 19858 43240
rect 19981 43231 20039 43237
rect 19981 43197 19993 43231
rect 20027 43197 20039 43231
rect 19981 43191 20039 43197
rect 18432 43132 19104 43160
rect 19076 43101 19104 43132
rect 19150 43120 19156 43172
rect 19208 43160 19214 43172
rect 19337 43163 19395 43169
rect 19337 43160 19349 43163
rect 19208 43132 19349 43160
rect 19208 43120 19214 43132
rect 19337 43129 19349 43132
rect 19383 43129 19395 43163
rect 19337 43123 19395 43129
rect 19429 43163 19487 43169
rect 19429 43129 19441 43163
rect 19475 43129 19487 43163
rect 19628 43160 19656 43188
rect 19996 43160 20024 43191
rect 19628 43132 20024 43160
rect 19429 43123 19487 43129
rect 18012 43064 18276 43092
rect 19061 43095 19119 43101
rect 18012 43052 18018 43064
rect 19061 43061 19073 43095
rect 19107 43061 19119 43095
rect 19444 43092 19472 43123
rect 19610 43092 19616 43104
rect 19444 43064 19616 43092
rect 19061 43055 19119 43061
rect 19610 43052 19616 43064
rect 19668 43092 19674 43104
rect 19797 43095 19855 43101
rect 19797 43092 19809 43095
rect 19668 43064 19809 43092
rect 19668 43052 19674 43064
rect 19797 43061 19809 43064
rect 19843 43092 19855 43095
rect 20088 43092 20116 43336
rect 20533 43231 20591 43237
rect 20533 43197 20545 43231
rect 20579 43228 20591 43231
rect 21269 43231 21327 43237
rect 21269 43228 21281 43231
rect 20579 43200 21281 43228
rect 20579 43197 20591 43200
rect 20533 43191 20591 43197
rect 21269 43197 21281 43200
rect 21315 43197 21327 43231
rect 21269 43191 21327 43197
rect 21545 43231 21603 43237
rect 21545 43197 21557 43231
rect 21591 43228 21603 43231
rect 21729 43231 21787 43237
rect 21729 43228 21741 43231
rect 21591 43200 21741 43228
rect 21591 43197 21603 43200
rect 21545 43191 21603 43197
rect 21729 43197 21741 43200
rect 21775 43228 21787 43231
rect 22370 43228 22376 43240
rect 21775 43200 22376 43228
rect 21775 43197 21787 43200
rect 21729 43191 21787 43197
rect 21284 43160 21312 43191
rect 22370 43188 22376 43200
rect 22428 43188 22434 43240
rect 24578 43188 24584 43240
rect 24636 43228 24642 43240
rect 24958 43231 25016 43237
rect 24958 43228 24970 43231
rect 24636 43200 24970 43228
rect 24636 43188 24642 43200
rect 24958 43197 24970 43200
rect 25004 43197 25016 43231
rect 24958 43191 25016 43197
rect 25225 43231 25283 43237
rect 25225 43197 25237 43231
rect 25271 43228 25283 43231
rect 25406 43228 25412 43240
rect 25271 43200 25412 43228
rect 25271 43197 25283 43200
rect 25225 43191 25283 43197
rect 25406 43188 25412 43200
rect 25464 43228 25470 43240
rect 26697 43231 26755 43237
rect 26697 43228 26709 43231
rect 25464 43200 26709 43228
rect 25464 43188 25470 43200
rect 26697 43197 26709 43200
rect 26743 43228 26755 43231
rect 27522 43228 27528 43240
rect 26743 43200 27528 43228
rect 26743 43197 26755 43200
rect 26697 43191 26755 43197
rect 27522 43188 27528 43200
rect 27580 43228 27586 43240
rect 28169 43231 28227 43237
rect 28169 43228 28181 43231
rect 27580 43200 28181 43228
rect 27580 43188 27586 43200
rect 28169 43197 28181 43200
rect 28215 43197 28227 43231
rect 28169 43191 28227 43197
rect 21634 43160 21640 43172
rect 21284 43132 21640 43160
rect 21634 43120 21640 43132
rect 21692 43120 21698 43172
rect 22002 43169 22008 43172
rect 21996 43123 22008 43169
rect 22002 43120 22008 43123
rect 22060 43120 22066 43172
rect 23290 43120 23296 43172
rect 23348 43120 23354 43172
rect 25682 43120 25688 43172
rect 25740 43160 25746 43172
rect 26430 43163 26488 43169
rect 26430 43160 26442 43163
rect 25740 43132 26442 43160
rect 25740 43120 25746 43132
rect 26430 43129 26442 43132
rect 26476 43129 26488 43163
rect 26430 43123 26488 43129
rect 27924 43163 27982 43169
rect 27924 43129 27936 43163
rect 27970 43160 27982 43163
rect 28074 43160 28080 43172
rect 27970 43132 28080 43160
rect 27970 43129 27982 43132
rect 27924 43123 27982 43129
rect 28074 43120 28080 43132
rect 28132 43120 28138 43172
rect 19843 43064 20116 43092
rect 20165 43095 20223 43101
rect 19843 43061 19855 43064
rect 19797 43055 19855 43061
rect 20165 43061 20177 43095
rect 20211 43092 20223 43095
rect 20254 43092 20260 43104
rect 20211 43064 20260 43092
rect 20211 43061 20223 43064
rect 20165 43055 20223 43061
rect 20254 43052 20260 43064
rect 20312 43052 20318 43104
rect 20346 43052 20352 43104
rect 20404 43052 20410 43104
rect 21082 43052 21088 43104
rect 21140 43052 21146 43104
rect 21266 43052 21272 43104
rect 21324 43092 21330 43104
rect 21453 43095 21511 43101
rect 21453 43092 21465 43095
rect 21324 43064 21465 43092
rect 21324 43052 21330 43064
rect 21453 43061 21465 43064
rect 21499 43061 21511 43095
rect 21453 43055 21511 43061
rect 23014 43052 23020 43104
rect 23072 43092 23078 43104
rect 23109 43095 23167 43101
rect 23109 43092 23121 43095
rect 23072 43064 23121 43092
rect 23072 43052 23078 43064
rect 23109 43061 23121 43064
rect 23155 43061 23167 43095
rect 23109 43055 23167 43061
rect 23566 43052 23572 43104
rect 23624 43052 23630 43104
rect 23845 43095 23903 43101
rect 23845 43061 23857 43095
rect 23891 43092 23903 43095
rect 24118 43092 24124 43104
rect 23891 43064 24124 43092
rect 23891 43061 23903 43064
rect 23845 43055 23903 43061
rect 24118 43052 24124 43064
rect 24176 43052 24182 43104
rect 25314 43052 25320 43104
rect 25372 43052 25378 43104
rect 26786 43052 26792 43104
rect 26844 43052 26850 43104
rect 552 43002 31648 43024
rect 552 42950 4322 43002
rect 4374 42950 4386 43002
rect 4438 42950 4450 43002
rect 4502 42950 4514 43002
rect 4566 42950 4578 43002
rect 4630 42950 12096 43002
rect 12148 42950 12160 43002
rect 12212 42950 12224 43002
rect 12276 42950 12288 43002
rect 12340 42950 12352 43002
rect 12404 42950 19870 43002
rect 19922 42950 19934 43002
rect 19986 42950 19998 43002
rect 20050 42950 20062 43002
rect 20114 42950 20126 43002
rect 20178 42950 27644 43002
rect 27696 42950 27708 43002
rect 27760 42950 27772 43002
rect 27824 42950 27836 43002
rect 27888 42950 27900 43002
rect 27952 42950 31648 43002
rect 552 42928 31648 42950
rect 11974 42848 11980 42900
rect 12032 42888 12038 42900
rect 12161 42891 12219 42897
rect 12161 42888 12173 42891
rect 12032 42860 12173 42888
rect 12032 42848 12038 42860
rect 12161 42857 12173 42860
rect 12207 42857 12219 42891
rect 12161 42851 12219 42857
rect 13909 42891 13967 42897
rect 13909 42857 13921 42891
rect 13955 42888 13967 42891
rect 13998 42888 14004 42900
rect 13955 42860 14004 42888
rect 13955 42857 13967 42860
rect 13909 42851 13967 42857
rect 13998 42848 14004 42860
rect 14056 42848 14062 42900
rect 14093 42891 14151 42897
rect 14093 42857 14105 42891
rect 14139 42888 14151 42891
rect 15010 42888 15016 42900
rect 14139 42860 15016 42888
rect 14139 42857 14151 42860
rect 14093 42851 14151 42857
rect 15010 42848 15016 42860
rect 15068 42848 15074 42900
rect 15470 42848 15476 42900
rect 15528 42888 15534 42900
rect 15657 42891 15715 42897
rect 15657 42888 15669 42891
rect 15528 42860 15669 42888
rect 15528 42848 15534 42860
rect 15657 42857 15669 42860
rect 15703 42888 15715 42891
rect 16298 42888 16304 42900
rect 15703 42860 16304 42888
rect 15703 42857 15715 42860
rect 15657 42851 15715 42857
rect 16298 42848 16304 42860
rect 16356 42848 16362 42900
rect 16666 42888 16672 42900
rect 16500 42860 16672 42888
rect 12268 42792 14044 42820
rect 9398 42712 9404 42764
rect 9456 42712 9462 42764
rect 9674 42761 9680 42764
rect 9668 42715 9680 42761
rect 9674 42712 9680 42715
rect 9732 42712 9738 42764
rect 11054 42712 11060 42764
rect 11112 42752 11118 42764
rect 12268 42761 12296 42792
rect 12253 42755 12311 42761
rect 12253 42752 12265 42755
rect 11112 42724 12265 42752
rect 11112 42712 11118 42724
rect 12253 42721 12265 42724
rect 12299 42721 12311 42755
rect 12253 42715 12311 42721
rect 12526 42712 12532 42764
rect 12584 42712 12590 42764
rect 12796 42755 12854 42761
rect 12796 42721 12808 42755
rect 12842 42752 12854 42755
rect 13538 42752 13544 42764
rect 12842 42724 13544 42752
rect 12842 42721 12854 42724
rect 12796 42715 12854 42721
rect 13538 42712 13544 42724
rect 13596 42712 13602 42764
rect 14016 42761 14044 42792
rect 14001 42755 14059 42761
rect 14001 42721 14013 42755
rect 14047 42752 14059 42755
rect 14642 42752 14648 42764
rect 14047 42724 14648 42752
rect 14047 42721 14059 42724
rect 14001 42715 14059 42721
rect 14642 42712 14648 42724
rect 14700 42712 14706 42764
rect 16206 42712 16212 42764
rect 16264 42752 16270 42764
rect 16500 42761 16528 42860
rect 16666 42848 16672 42860
rect 16724 42848 16730 42900
rect 19702 42848 19708 42900
rect 19760 42848 19766 42900
rect 22649 42891 22707 42897
rect 22649 42857 22661 42891
rect 22695 42888 22707 42891
rect 23290 42888 23296 42900
rect 22695 42860 23296 42888
rect 22695 42857 22707 42860
rect 22649 42851 22707 42857
rect 23290 42848 23296 42860
rect 23348 42848 23354 42900
rect 24486 42888 24492 42900
rect 23860 42860 24492 42888
rect 17126 42820 17132 42832
rect 16684 42792 17132 42820
rect 16684 42761 16712 42792
rect 17126 42780 17132 42792
rect 17184 42780 17190 42832
rect 17497 42823 17555 42829
rect 17497 42820 17509 42823
rect 17236 42792 17509 42820
rect 16942 42761 16948 42764
rect 16393 42755 16451 42761
rect 16393 42752 16405 42755
rect 16264 42724 16405 42752
rect 16264 42712 16270 42724
rect 16393 42721 16405 42724
rect 16439 42721 16451 42755
rect 16393 42715 16451 42721
rect 16486 42755 16544 42761
rect 16486 42721 16498 42755
rect 16532 42721 16544 42755
rect 16486 42715 16544 42721
rect 16669 42755 16727 42761
rect 16669 42721 16681 42755
rect 16715 42721 16727 42755
rect 16669 42715 16727 42721
rect 16761 42755 16819 42761
rect 16761 42721 16773 42755
rect 16807 42721 16819 42755
rect 16761 42715 16819 42721
rect 16897 42755 16948 42761
rect 16897 42721 16909 42755
rect 16943 42721 16948 42755
rect 16897 42715 16948 42721
rect 11330 42684 11336 42696
rect 10796 42656 11336 42684
rect 10796 42625 10824 42656
rect 11330 42644 11336 42656
rect 11388 42684 11394 42696
rect 11517 42687 11575 42693
rect 11517 42684 11529 42687
rect 11388 42656 11529 42684
rect 11388 42644 11394 42656
rect 11517 42653 11529 42656
rect 11563 42653 11575 42687
rect 11517 42647 11575 42653
rect 14274 42644 14280 42696
rect 14332 42644 14338 42696
rect 14553 42687 14611 42693
rect 14553 42653 14565 42687
rect 14599 42684 14611 42687
rect 15010 42684 15016 42696
rect 14599 42656 15016 42684
rect 14599 42653 14611 42656
rect 14553 42647 14611 42653
rect 15010 42644 15016 42656
rect 15068 42644 15074 42696
rect 16298 42644 16304 42696
rect 16356 42684 16362 42696
rect 16776 42684 16804 42715
rect 16356 42656 16804 42684
rect 16914 42712 16948 42715
rect 17000 42752 17006 42764
rect 17236 42752 17264 42792
rect 17497 42789 17509 42792
rect 17543 42820 17555 42823
rect 18138 42820 18144 42832
rect 17543 42792 18144 42820
rect 17543 42789 17555 42792
rect 17497 42783 17555 42789
rect 18138 42780 18144 42792
rect 18196 42780 18202 42832
rect 20530 42780 20536 42832
rect 20588 42820 20594 42832
rect 20588 42792 22968 42820
rect 20588 42780 20594 42792
rect 22940 42764 22968 42792
rect 17000 42724 17264 42752
rect 17000 42712 17006 42724
rect 17402 42712 17408 42764
rect 17460 42712 17466 42764
rect 17681 42755 17739 42761
rect 17681 42721 17693 42755
rect 17727 42752 17739 42755
rect 17954 42752 17960 42764
rect 17727 42724 17960 42752
rect 17727 42721 17739 42724
rect 17681 42715 17739 42721
rect 17954 42712 17960 42724
rect 18012 42712 18018 42764
rect 19518 42712 19524 42764
rect 19576 42752 19582 42764
rect 19613 42755 19671 42761
rect 19613 42752 19625 42755
rect 19576 42724 19625 42752
rect 19576 42712 19582 42724
rect 19613 42721 19625 42724
rect 19659 42721 19671 42755
rect 19613 42715 19671 42721
rect 19981 42755 20039 42761
rect 19981 42721 19993 42755
rect 20027 42721 20039 42755
rect 19981 42715 20039 42721
rect 16356 42644 16362 42656
rect 10781 42619 10839 42625
rect 10781 42585 10793 42619
rect 10827 42585 10839 42619
rect 10781 42579 10839 42585
rect 16022 42576 16028 42628
rect 16080 42616 16086 42628
rect 16914 42616 16942 42712
rect 19337 42687 19395 42693
rect 19337 42653 19349 42687
rect 19383 42684 19395 42687
rect 19383 42656 19656 42684
rect 19383 42653 19395 42656
rect 19337 42647 19395 42653
rect 19628 42628 19656 42656
rect 16080 42588 16942 42616
rect 16080 42576 16086 42588
rect 19610 42576 19616 42628
rect 19668 42576 19674 42628
rect 10962 42508 10968 42560
rect 11020 42508 11026 42560
rect 17037 42551 17095 42557
rect 17037 42517 17049 42551
rect 17083 42548 17095 42551
rect 17494 42548 17500 42560
rect 17083 42520 17500 42548
rect 17083 42517 17095 42520
rect 17037 42511 17095 42517
rect 17494 42508 17500 42520
rect 17552 42508 17558 42560
rect 17865 42551 17923 42557
rect 17865 42517 17877 42551
rect 17911 42548 17923 42551
rect 18966 42548 18972 42560
rect 17911 42520 18972 42548
rect 17911 42517 17923 42520
rect 17865 42511 17923 42517
rect 18966 42508 18972 42520
rect 19024 42508 19030 42560
rect 19150 42508 19156 42560
rect 19208 42548 19214 42560
rect 19996 42548 20024 42715
rect 20070 42712 20076 42764
rect 20128 42712 20134 42764
rect 20165 42755 20223 42761
rect 20165 42721 20177 42755
rect 20211 42752 20223 42755
rect 20254 42752 20260 42764
rect 20211 42724 20260 42752
rect 20211 42721 20223 42724
rect 20165 42715 20223 42721
rect 20254 42712 20260 42724
rect 20312 42712 20318 42764
rect 20346 42712 20352 42764
rect 20404 42712 20410 42764
rect 21266 42712 21272 42764
rect 21324 42712 21330 42764
rect 21358 42712 21364 42764
rect 21416 42752 21422 42764
rect 21525 42755 21583 42761
rect 21525 42752 21537 42755
rect 21416 42724 21537 42752
rect 21416 42712 21422 42724
rect 21525 42721 21537 42724
rect 21571 42721 21583 42755
rect 21525 42715 21583 42721
rect 22922 42712 22928 42764
rect 22980 42712 22986 42764
rect 23014 42712 23020 42764
rect 23072 42712 23078 42764
rect 23201 42755 23259 42761
rect 23201 42721 23213 42755
rect 23247 42721 23259 42755
rect 23201 42715 23259 42721
rect 23216 42684 23244 42715
rect 23290 42712 23296 42764
rect 23348 42712 23354 42764
rect 23474 42712 23480 42764
rect 23532 42752 23538 42764
rect 23569 42755 23627 42761
rect 23569 42752 23581 42755
rect 23532 42724 23581 42752
rect 23532 42712 23538 42724
rect 23569 42721 23581 42724
rect 23615 42721 23627 42755
rect 23569 42715 23627 42721
rect 23661 42755 23719 42761
rect 23661 42721 23673 42755
rect 23707 42721 23719 42755
rect 23661 42715 23719 42721
rect 23385 42687 23443 42693
rect 23385 42684 23397 42687
rect 23216 42656 23397 42684
rect 23385 42653 23397 42656
rect 23431 42653 23443 42687
rect 23676 42684 23704 42715
rect 23750 42712 23756 42764
rect 23808 42752 23814 42764
rect 23860 42761 23888 42860
rect 24486 42848 24492 42860
rect 24544 42848 24550 42900
rect 25222 42820 25228 42832
rect 24412 42792 25228 42820
rect 23845 42755 23903 42761
rect 23845 42752 23857 42755
rect 23808 42724 23857 42752
rect 23808 42712 23814 42724
rect 23845 42721 23857 42724
rect 23891 42721 23903 42755
rect 23845 42715 23903 42721
rect 23934 42712 23940 42764
rect 23992 42712 23998 42764
rect 24026 42712 24032 42764
rect 24084 42752 24090 42764
rect 24213 42755 24271 42761
rect 24213 42752 24225 42755
rect 24084 42724 24225 42752
rect 24084 42712 24090 42724
rect 24213 42721 24225 42724
rect 24259 42721 24271 42755
rect 24213 42715 24271 42721
rect 24305 42755 24363 42761
rect 24305 42721 24317 42755
rect 24351 42752 24363 42755
rect 24412 42752 24440 42792
rect 25222 42780 25228 42792
rect 25280 42780 25286 42832
rect 24351 42724 24440 42752
rect 24351 42721 24363 42724
rect 24305 42715 24363 42721
rect 24486 42712 24492 42764
rect 24544 42712 24550 42764
rect 24578 42712 24584 42764
rect 24636 42712 24642 42764
rect 27522 42712 27528 42764
rect 27580 42752 27586 42764
rect 29641 42755 29699 42761
rect 29641 42752 29653 42755
rect 27580 42724 29653 42752
rect 27580 42712 27586 42724
rect 29641 42721 29653 42724
rect 29687 42721 29699 42755
rect 29641 42715 29699 42721
rect 25314 42684 25320 42696
rect 23676 42656 25320 42684
rect 23385 42647 23443 42653
rect 25314 42644 25320 42656
rect 25372 42644 25378 42696
rect 22646 42576 22652 42628
rect 22704 42616 22710 42628
rect 23934 42616 23940 42628
rect 22704 42588 23940 42616
rect 22704 42576 22710 42588
rect 23934 42576 23940 42588
rect 23992 42576 23998 42628
rect 24210 42576 24216 42628
rect 24268 42616 24274 42628
rect 29270 42616 29276 42628
rect 24268 42588 29276 42616
rect 24268 42576 24274 42588
rect 29270 42576 29276 42588
rect 29328 42576 29334 42628
rect 19208 42520 20024 42548
rect 19208 42508 19214 42520
rect 22278 42508 22284 42560
rect 22336 42548 22342 42560
rect 22741 42551 22799 42557
rect 22741 42548 22753 42551
rect 22336 42520 22753 42548
rect 22336 42508 22342 42520
rect 22741 42517 22753 42520
rect 22787 42517 22799 42551
rect 22741 42511 22799 42517
rect 23382 42508 23388 42560
rect 23440 42548 23446 42560
rect 24029 42551 24087 42557
rect 24029 42548 24041 42551
rect 23440 42520 24041 42548
rect 23440 42508 23446 42520
rect 24029 42517 24041 42520
rect 24075 42517 24087 42551
rect 24029 42511 24087 42517
rect 29362 42508 29368 42560
rect 29420 42548 29426 42560
rect 29549 42551 29607 42557
rect 29549 42548 29561 42551
rect 29420 42520 29561 42548
rect 29420 42508 29426 42520
rect 29549 42517 29561 42520
rect 29595 42517 29607 42551
rect 29549 42511 29607 42517
rect 552 42458 31648 42480
rect 552 42406 3662 42458
rect 3714 42406 3726 42458
rect 3778 42406 3790 42458
rect 3842 42406 3854 42458
rect 3906 42406 3918 42458
rect 3970 42406 11436 42458
rect 11488 42406 11500 42458
rect 11552 42406 11564 42458
rect 11616 42406 11628 42458
rect 11680 42406 11692 42458
rect 11744 42406 19210 42458
rect 19262 42406 19274 42458
rect 19326 42406 19338 42458
rect 19390 42406 19402 42458
rect 19454 42406 19466 42458
rect 19518 42406 26984 42458
rect 27036 42406 27048 42458
rect 27100 42406 27112 42458
rect 27164 42406 27176 42458
rect 27228 42406 27240 42458
rect 27292 42406 31648 42458
rect 552 42384 31648 42406
rect 13538 42304 13544 42356
rect 13596 42304 13602 42356
rect 14274 42304 14280 42356
rect 14332 42344 14338 42356
rect 14737 42347 14795 42353
rect 14737 42344 14749 42347
rect 14332 42316 14749 42344
rect 14332 42304 14338 42316
rect 14737 42313 14749 42316
rect 14783 42313 14795 42347
rect 14737 42307 14795 42313
rect 15010 42304 15016 42356
rect 15068 42304 15074 42356
rect 17034 42304 17040 42356
rect 17092 42344 17098 42356
rect 17129 42347 17187 42353
rect 17129 42344 17141 42347
rect 17092 42316 17141 42344
rect 17092 42304 17098 42316
rect 17129 42313 17141 42316
rect 17175 42313 17187 42347
rect 17129 42307 17187 42313
rect 17310 42304 17316 42356
rect 17368 42304 17374 42356
rect 18690 42344 18696 42356
rect 17512 42316 18696 42344
rect 15470 42276 15476 42288
rect 15212 42248 15476 42276
rect 13722 42100 13728 42152
rect 13780 42100 13786 42152
rect 13998 42100 14004 42152
rect 14056 42100 14062 42152
rect 14182 42100 14188 42152
rect 14240 42100 14246 42152
rect 14642 42100 14648 42152
rect 14700 42100 14706 42152
rect 15212 42149 15240 42248
rect 15470 42236 15476 42248
rect 15528 42236 15534 42288
rect 16390 42236 16396 42288
rect 16448 42236 16454 42288
rect 15381 42211 15439 42217
rect 15381 42177 15393 42211
rect 15427 42208 15439 42211
rect 15654 42208 15660 42220
rect 15427 42180 15660 42208
rect 15427 42177 15439 42180
rect 15381 42171 15439 42177
rect 15654 42168 15660 42180
rect 15712 42168 15718 42220
rect 16408 42208 16436 42236
rect 16850 42208 16856 42220
rect 16408 42180 16528 42208
rect 15197 42143 15255 42149
rect 15197 42109 15209 42143
rect 15243 42109 15255 42143
rect 15197 42103 15255 42109
rect 15470 42100 15476 42152
rect 15528 42100 15534 42152
rect 15565 42143 15623 42149
rect 15565 42109 15577 42143
rect 15611 42109 15623 42143
rect 15565 42103 15623 42109
rect 15580 42072 15608 42103
rect 15746 42100 15752 42152
rect 15804 42100 15810 42152
rect 16500 42149 16528 42180
rect 16684 42180 16856 42208
rect 16684 42149 16712 42180
rect 16850 42168 16856 42180
rect 16908 42168 16914 42220
rect 16301 42143 16359 42149
rect 16301 42109 16313 42143
rect 16347 42109 16359 42143
rect 16301 42103 16359 42109
rect 16393 42143 16451 42149
rect 16393 42109 16405 42143
rect 16439 42109 16451 42143
rect 16393 42103 16451 42109
rect 16485 42143 16543 42149
rect 16485 42109 16497 42143
rect 16531 42109 16543 42143
rect 16485 42103 16543 42109
rect 16669 42143 16727 42149
rect 16669 42109 16681 42143
rect 16715 42109 16727 42143
rect 16669 42103 16727 42109
rect 16025 42075 16083 42081
rect 16025 42072 16037 42075
rect 15580 42044 16037 42072
rect 16025 42041 16037 42044
rect 16071 42041 16083 42075
rect 16025 42035 16083 42041
rect 15194 41964 15200 42016
rect 15252 42004 15258 42016
rect 15746 42004 15752 42016
rect 15252 41976 15752 42004
rect 15252 41964 15258 41976
rect 15746 41964 15752 41976
rect 15804 41964 15810 42016
rect 16316 42004 16344 42103
rect 16408 42072 16436 42103
rect 16758 42100 16764 42152
rect 16816 42100 16822 42152
rect 16942 42100 16948 42152
rect 17000 42100 17006 42152
rect 16853 42075 16911 42081
rect 16853 42072 16865 42075
rect 16408 42044 16865 42072
rect 16853 42041 16865 42044
rect 16899 42041 16911 42075
rect 16853 42035 16911 42041
rect 17218 42032 17224 42084
rect 17276 42081 17282 42084
rect 17512 42081 17540 42316
rect 18690 42304 18696 42316
rect 18748 42304 18754 42356
rect 19426 42304 19432 42356
rect 19484 42344 19490 42356
rect 19610 42344 19616 42356
rect 19484 42316 19616 42344
rect 19484 42304 19490 42316
rect 19610 42304 19616 42316
rect 19668 42304 19674 42356
rect 20993 42347 21051 42353
rect 20993 42313 21005 42347
rect 21039 42344 21051 42347
rect 21358 42344 21364 42356
rect 21039 42316 21364 42344
rect 21039 42313 21051 42316
rect 20993 42307 21051 42313
rect 21358 42304 21364 42316
rect 21416 42304 21422 42356
rect 23290 42304 23296 42356
rect 23348 42344 23354 42356
rect 23845 42347 23903 42353
rect 23845 42344 23857 42347
rect 23348 42316 23857 42344
rect 23348 42304 23354 42316
rect 23845 42313 23857 42316
rect 23891 42313 23903 42347
rect 23845 42307 23903 42313
rect 18417 42279 18475 42285
rect 18417 42245 18429 42279
rect 18463 42245 18475 42279
rect 18417 42239 18475 42245
rect 18432 42208 18460 42239
rect 18966 42236 18972 42288
rect 19024 42236 19030 42288
rect 19521 42279 19579 42285
rect 19521 42245 19533 42279
rect 19567 42276 19579 42279
rect 20070 42276 20076 42288
rect 19567 42248 20076 42276
rect 19567 42245 19579 42248
rect 19521 42239 19579 42245
rect 20070 42236 20076 42248
rect 20128 42236 20134 42288
rect 23658 42276 23664 42288
rect 22066 42248 23664 42276
rect 18984 42208 19012 42236
rect 21082 42208 21088 42220
rect 18432 42180 18828 42208
rect 18506 42149 18512 42152
rect 18484 42143 18512 42149
rect 18325 42133 18383 42139
rect 18325 42099 18337 42133
rect 18371 42099 18383 42133
rect 18484 42109 18496 42143
rect 18484 42103 18512 42109
rect 18506 42100 18512 42103
rect 18564 42100 18570 42152
rect 18690 42100 18696 42152
rect 18748 42100 18754 42152
rect 18325 42093 18383 42099
rect 17276 42075 17339 42081
rect 17276 42041 17293 42075
rect 17327 42041 17339 42075
rect 17276 42035 17339 42041
rect 17497 42075 17555 42081
rect 17497 42041 17509 42075
rect 17543 42041 17555 42075
rect 17497 42035 17555 42041
rect 17276 42032 17282 42035
rect 18340 42016 18368 42093
rect 18138 42004 18144 42016
rect 16316 41976 18144 42004
rect 18138 41964 18144 41976
rect 18196 41964 18202 42016
rect 18322 41964 18328 42016
rect 18380 41964 18386 42016
rect 18708 42004 18736 42100
rect 18800 42072 18828 42180
rect 18892 42180 19012 42208
rect 20364 42180 21088 42208
rect 18892 42149 18920 42180
rect 18877 42143 18935 42149
rect 18877 42109 18889 42143
rect 18923 42109 18935 42143
rect 18877 42103 18935 42109
rect 18969 42143 19027 42149
rect 18969 42109 18981 42143
rect 19015 42109 19027 42143
rect 18969 42103 19027 42109
rect 18984 42072 19012 42103
rect 19058 42100 19064 42152
rect 19116 42100 19122 42152
rect 19150 42100 19156 42152
rect 19208 42140 19214 42152
rect 19429 42143 19487 42149
rect 19429 42140 19441 42143
rect 19208 42112 19441 42140
rect 19208 42100 19214 42112
rect 19429 42109 19441 42112
rect 19475 42109 19487 42143
rect 19429 42103 19487 42109
rect 18800 42044 19012 42072
rect 19334 42032 19340 42084
rect 19392 42032 19398 42084
rect 19444 42072 19472 42103
rect 19518 42100 19524 42152
rect 19576 42140 19582 42152
rect 19613 42143 19671 42149
rect 19613 42140 19625 42143
rect 19576 42112 19625 42140
rect 19576 42100 19582 42112
rect 19613 42109 19625 42112
rect 19659 42109 19671 42143
rect 19613 42103 19671 42109
rect 19702 42100 19708 42152
rect 19760 42140 19766 42152
rect 20073 42143 20131 42149
rect 20073 42140 20085 42143
rect 19760 42112 20085 42140
rect 19760 42100 19766 42112
rect 20073 42109 20085 42112
rect 20119 42109 20131 42143
rect 20073 42103 20131 42109
rect 20254 42100 20260 42152
rect 20312 42100 20318 42152
rect 20364 42149 20392 42180
rect 21082 42168 21088 42180
rect 21140 42168 21146 42220
rect 21269 42211 21327 42217
rect 21269 42177 21281 42211
rect 21315 42208 21327 42211
rect 22066 42208 22094 42248
rect 23658 42236 23664 42248
rect 23716 42276 23722 42288
rect 24210 42276 24216 42288
rect 23716 42248 24216 42276
rect 23716 42236 23722 42248
rect 24210 42236 24216 42248
rect 24268 42236 24274 42288
rect 26786 42208 26792 42220
rect 21315 42180 22094 42208
rect 23124 42180 26792 42208
rect 21315 42177 21327 42180
rect 21269 42171 21327 42177
rect 20349 42143 20407 42149
rect 20349 42109 20361 42143
rect 20395 42109 20407 42143
rect 20349 42103 20407 42109
rect 20533 42143 20591 42149
rect 20533 42109 20545 42143
rect 20579 42109 20591 42143
rect 20533 42103 20591 42109
rect 20625 42143 20683 42149
rect 20625 42109 20637 42143
rect 20671 42109 20683 42143
rect 20625 42103 20683 42109
rect 20717 42143 20775 42149
rect 20717 42109 20729 42143
rect 20763 42140 20775 42143
rect 20806 42140 20812 42152
rect 20763 42112 20812 42140
rect 20763 42109 20775 42112
rect 20717 42103 20775 42109
rect 19794 42072 19800 42084
rect 19444 42044 19800 42072
rect 19794 42032 19800 42044
rect 19852 42032 19858 42084
rect 20165 42075 20223 42081
rect 20165 42041 20177 42075
rect 20211 42072 20223 42075
rect 20548 42072 20576 42103
rect 20211 42044 20576 42072
rect 20211 42041 20223 42044
rect 20165 42035 20223 42041
rect 20346 42004 20352 42016
rect 18708 41976 20352 42004
rect 20346 41964 20352 41976
rect 20404 41964 20410 42016
rect 20438 41964 20444 42016
rect 20496 42004 20502 42016
rect 20640 42004 20668 42103
rect 20806 42100 20812 42112
rect 20864 42100 20870 42152
rect 20990 42100 20996 42152
rect 21048 42140 21054 42152
rect 21284 42140 21312 42171
rect 21048 42112 21312 42140
rect 21545 42143 21603 42149
rect 21048 42100 21054 42112
rect 21545 42109 21557 42143
rect 21591 42140 21603 42143
rect 21634 42140 21640 42152
rect 21591 42112 21640 42140
rect 21591 42109 21603 42112
rect 21545 42103 21603 42109
rect 21634 42100 21640 42112
rect 21692 42140 21698 42152
rect 22002 42140 22008 42152
rect 21692 42112 22008 42140
rect 21692 42100 21698 42112
rect 22002 42100 22008 42112
rect 22060 42100 22066 42152
rect 22370 42100 22376 42152
rect 22428 42100 22434 42152
rect 22922 42100 22928 42152
rect 22980 42140 22986 42152
rect 23124 42149 23152 42180
rect 26786 42168 26792 42180
rect 26844 42168 26850 42220
rect 23017 42143 23075 42149
rect 23017 42140 23029 42143
rect 22980 42112 23029 42140
rect 22980 42100 22986 42112
rect 23017 42109 23029 42112
rect 23063 42109 23075 42143
rect 23017 42103 23075 42109
rect 23109 42143 23167 42149
rect 23109 42109 23121 42143
rect 23155 42109 23167 42143
rect 23109 42103 23167 42109
rect 23198 42100 23204 42152
rect 23256 42140 23262 42152
rect 23293 42143 23351 42149
rect 23293 42140 23305 42143
rect 23256 42112 23305 42140
rect 23256 42100 23262 42112
rect 23293 42109 23305 42112
rect 23339 42109 23351 42143
rect 23293 42103 23351 42109
rect 23382 42100 23388 42152
rect 23440 42100 23446 42152
rect 24026 42100 24032 42152
rect 24084 42100 24090 42152
rect 24118 42100 24124 42152
rect 24176 42100 24182 42152
rect 24394 42100 24400 42152
rect 24452 42100 24458 42152
rect 26234 42100 26240 42152
rect 26292 42140 26298 42152
rect 26697 42143 26755 42149
rect 26697 42140 26709 42143
rect 26292 42112 26709 42140
rect 26292 42100 26298 42112
rect 26697 42109 26709 42112
rect 26743 42140 26755 42143
rect 27522 42140 27528 42152
rect 26743 42112 27528 42140
rect 26743 42109 26755 42112
rect 26697 42103 26755 42109
rect 27522 42100 27528 42112
rect 27580 42140 27586 42152
rect 28169 42143 28227 42149
rect 28169 42140 28181 42143
rect 27580 42112 28181 42140
rect 27580 42100 27586 42112
rect 28169 42109 28181 42112
rect 28215 42109 28227 42143
rect 28169 42103 28227 42109
rect 29546 42100 29552 42152
rect 29604 42100 29610 42152
rect 30377 42143 30435 42149
rect 30377 42109 30389 42143
rect 30423 42140 30435 42143
rect 30742 42140 30748 42152
rect 30423 42112 30748 42140
rect 30423 42109 30435 42112
rect 30377 42103 30435 42109
rect 20824 42072 20852 42100
rect 23566 42072 23572 42084
rect 20824 42044 23572 42072
rect 23566 42032 23572 42044
rect 23624 42032 23630 42084
rect 24213 42075 24271 42081
rect 24213 42041 24225 42075
rect 24259 42041 24271 42075
rect 24213 42035 24271 42041
rect 20496 41976 20668 42004
rect 20496 41964 20502 41976
rect 20990 41964 20996 42016
rect 21048 42004 21054 42016
rect 21085 42007 21143 42013
rect 21085 42004 21097 42007
rect 21048 41976 21097 42004
rect 21048 41964 21054 41976
rect 21085 41973 21097 41976
rect 21131 41973 21143 42007
rect 21085 41967 21143 41973
rect 21266 41964 21272 42016
rect 21324 42004 21330 42016
rect 22281 42007 22339 42013
rect 22281 42004 22293 42007
rect 21324 41976 22293 42004
rect 21324 41964 21330 41976
rect 22281 41973 22293 41976
rect 22327 41973 22339 42007
rect 22281 41967 22339 41973
rect 22830 41964 22836 42016
rect 22888 41964 22894 42016
rect 22922 41964 22928 42016
rect 22980 42004 22986 42016
rect 24228 42004 24256 42035
rect 28718 42032 28724 42084
rect 28776 42072 28782 42084
rect 30392 42072 30420 42103
rect 30742 42100 30748 42112
rect 30800 42100 30806 42152
rect 28776 42044 30420 42072
rect 28776 42032 28782 42044
rect 22980 41976 24256 42004
rect 22980 41964 22986 41976
rect 26418 41964 26424 42016
rect 26476 42004 26482 42016
rect 26605 42007 26663 42013
rect 26605 42004 26617 42007
rect 26476 41976 26617 42004
rect 26476 41964 26482 41976
rect 26605 41973 26617 41976
rect 26651 41973 26663 42007
rect 26605 41967 26663 41973
rect 27982 41964 27988 42016
rect 28040 42004 28046 42016
rect 28077 42007 28135 42013
rect 28077 42004 28089 42007
rect 28040 41976 28089 42004
rect 28040 41964 28046 41976
rect 28077 41973 28089 41976
rect 28123 41973 28135 42007
rect 28077 41967 28135 41973
rect 28994 41964 29000 42016
rect 29052 41964 29058 42016
rect 29270 41964 29276 42016
rect 29328 42004 29334 42016
rect 29733 42007 29791 42013
rect 29733 42004 29745 42007
rect 29328 41976 29745 42004
rect 29328 41964 29334 41976
rect 29733 41973 29745 41976
rect 29779 41973 29791 42007
rect 29733 41967 29791 41973
rect 552 41914 31648 41936
rect 552 41862 4322 41914
rect 4374 41862 4386 41914
rect 4438 41862 4450 41914
rect 4502 41862 4514 41914
rect 4566 41862 4578 41914
rect 4630 41862 12096 41914
rect 12148 41862 12160 41914
rect 12212 41862 12224 41914
rect 12276 41862 12288 41914
rect 12340 41862 12352 41914
rect 12404 41862 19870 41914
rect 19922 41862 19934 41914
rect 19986 41862 19998 41914
rect 20050 41862 20062 41914
rect 20114 41862 20126 41914
rect 20178 41862 27644 41914
rect 27696 41862 27708 41914
rect 27760 41862 27772 41914
rect 27824 41862 27836 41914
rect 27888 41862 27900 41914
rect 27952 41862 31648 41914
rect 552 41840 31648 41862
rect 9674 41760 9680 41812
rect 9732 41760 9738 41812
rect 13814 41760 13820 41812
rect 13872 41800 13878 41812
rect 14274 41800 14280 41812
rect 13872 41772 14280 41800
rect 13872 41760 13878 41772
rect 14274 41760 14280 41772
rect 14332 41760 14338 41812
rect 16758 41760 16764 41812
rect 16816 41800 16822 41812
rect 17126 41800 17132 41812
rect 16816 41772 17132 41800
rect 16816 41760 16822 41772
rect 17126 41760 17132 41772
rect 17184 41800 17190 41812
rect 18049 41803 18107 41809
rect 18049 41800 18061 41803
rect 17184 41772 18061 41800
rect 17184 41760 17190 41772
rect 18049 41769 18061 41772
rect 18095 41769 18107 41803
rect 18049 41763 18107 41769
rect 18506 41760 18512 41812
rect 18564 41800 18570 41812
rect 20070 41800 20076 41812
rect 18564 41772 20076 41800
rect 18564 41760 18570 41772
rect 20070 41760 20076 41772
rect 20128 41800 20134 41812
rect 24026 41800 24032 41812
rect 20128 41772 24032 41800
rect 20128 41760 20134 41772
rect 24026 41760 24032 41772
rect 24084 41760 24090 41812
rect 28810 41760 28816 41812
rect 28868 41800 28874 41812
rect 29273 41803 29331 41809
rect 29273 41800 29285 41803
rect 28868 41772 29285 41800
rect 28868 41760 28874 41772
rect 29273 41769 29285 41772
rect 29319 41800 29331 41803
rect 29546 41800 29552 41812
rect 29319 41772 29552 41800
rect 29319 41769 29331 41772
rect 29273 41763 29331 41769
rect 29546 41760 29552 41772
rect 29604 41760 29610 41812
rect 30742 41760 30748 41812
rect 30800 41760 30806 41812
rect 10962 41732 10968 41744
rect 9968 41704 10968 41732
rect 9968 41673 9996 41704
rect 10962 41692 10968 41704
rect 11020 41692 11026 41744
rect 16206 41692 16212 41744
rect 16264 41732 16270 41744
rect 20254 41732 20260 41744
rect 16264 41704 20260 41732
rect 16264 41692 16270 41704
rect 20254 41692 20260 41704
rect 20312 41732 20318 41744
rect 22646 41732 22652 41744
rect 20312 41704 22652 41732
rect 20312 41692 20318 41704
rect 22646 41692 22652 41704
rect 22704 41692 22710 41744
rect 9953 41667 10011 41673
rect 9953 41633 9965 41667
rect 9999 41633 10011 41667
rect 9953 41627 10011 41633
rect 10045 41667 10103 41673
rect 10045 41633 10057 41667
rect 10091 41633 10103 41667
rect 10045 41627 10103 41633
rect 10060 41596 10088 41627
rect 10134 41624 10140 41676
rect 10192 41624 10198 41676
rect 10318 41624 10324 41676
rect 10376 41664 10382 41676
rect 10778 41664 10784 41676
rect 10376 41636 10784 41664
rect 10376 41624 10382 41636
rect 10778 41624 10784 41636
rect 10836 41624 10842 41676
rect 13725 41667 13783 41673
rect 13725 41633 13737 41667
rect 13771 41633 13783 41667
rect 13725 41627 13783 41633
rect 13909 41667 13967 41673
rect 13909 41633 13921 41667
rect 13955 41664 13967 41667
rect 13998 41664 14004 41676
rect 13955 41636 14004 41664
rect 13955 41633 13967 41636
rect 13909 41627 13967 41633
rect 10410 41596 10416 41608
rect 10060 41568 10416 41596
rect 10410 41556 10416 41568
rect 10468 41556 10474 41608
rect 12710 41556 12716 41608
rect 12768 41596 12774 41608
rect 12989 41599 13047 41605
rect 12989 41596 13001 41599
rect 12768 41568 13001 41596
rect 12768 41556 12774 41568
rect 12989 41565 13001 41568
rect 13035 41565 13047 41599
rect 13740 41596 13768 41627
rect 13998 41624 14004 41636
rect 14056 41664 14062 41676
rect 14826 41664 14832 41676
rect 14056 41636 14832 41664
rect 14056 41624 14062 41636
rect 14826 41624 14832 41636
rect 14884 41624 14890 41676
rect 17862 41624 17868 41676
rect 17920 41624 17926 41676
rect 21266 41624 21272 41676
rect 21324 41624 21330 41676
rect 21358 41624 21364 41676
rect 21416 41664 21422 41676
rect 21525 41667 21583 41673
rect 21525 41664 21537 41667
rect 21416 41636 21537 41664
rect 21416 41624 21422 41636
rect 21525 41633 21537 41636
rect 21571 41633 21583 41667
rect 22741 41667 22799 41673
rect 22741 41664 22753 41667
rect 21525 41627 21583 41633
rect 22664 41636 22753 41664
rect 19610 41596 19616 41608
rect 13740 41568 19616 41596
rect 12989 41559 13047 41565
rect 19610 41556 19616 41568
rect 19668 41596 19674 41608
rect 20438 41596 20444 41608
rect 19668 41568 20444 41596
rect 19668 41556 19674 41568
rect 20438 41556 20444 41568
rect 20496 41556 20502 41608
rect 15010 41488 15016 41540
rect 15068 41528 15074 41540
rect 15838 41528 15844 41540
rect 15068 41500 15844 41528
rect 15068 41488 15074 41500
rect 15838 41488 15844 41500
rect 15896 41488 15902 41540
rect 16114 41488 16120 41540
rect 16172 41528 16178 41540
rect 20990 41528 20996 41540
rect 16172 41500 20996 41528
rect 16172 41488 16178 41500
rect 20990 41488 20996 41500
rect 21048 41488 21054 41540
rect 22664 41537 22692 41636
rect 22741 41633 22753 41636
rect 22787 41633 22799 41667
rect 22741 41627 22799 41633
rect 23198 41624 23204 41676
rect 23256 41624 23262 41676
rect 23934 41624 23940 41676
rect 23992 41624 23998 41676
rect 26418 41624 26424 41676
rect 26476 41624 26482 41676
rect 26694 41673 26700 41676
rect 26688 41627 26700 41673
rect 26694 41624 26700 41627
rect 26752 41624 26758 41676
rect 27893 41667 27951 41673
rect 27893 41633 27905 41667
rect 27939 41664 27951 41667
rect 27982 41664 27988 41676
rect 27939 41636 27988 41664
rect 27939 41633 27951 41636
rect 27893 41627 27951 41633
rect 27982 41624 27988 41636
rect 28040 41624 28046 41676
rect 28166 41673 28172 41676
rect 28160 41664 28172 41673
rect 28127 41636 28172 41664
rect 28160 41627 28172 41636
rect 28166 41624 28172 41627
rect 28224 41624 28230 41676
rect 29362 41624 29368 41676
rect 29420 41624 29426 41676
rect 29454 41624 29460 41676
rect 29512 41664 29518 41676
rect 29621 41667 29679 41673
rect 29621 41664 29633 41667
rect 29512 41636 29633 41664
rect 29512 41624 29518 41636
rect 29621 41633 29633 41636
rect 29667 41633 29679 41667
rect 29621 41627 29679 41633
rect 22649 41531 22707 41537
rect 22649 41497 22661 41531
rect 22695 41497 22707 41531
rect 22649 41491 22707 41497
rect 22925 41531 22983 41537
rect 22925 41497 22937 41531
rect 22971 41528 22983 41531
rect 23934 41528 23940 41540
rect 22971 41500 23940 41528
rect 22971 41497 22983 41500
rect 22925 41491 22983 41497
rect 23934 41488 23940 41500
rect 23992 41488 23998 41540
rect 12434 41420 12440 41472
rect 12492 41420 12498 41472
rect 15378 41420 15384 41472
rect 15436 41460 15442 41472
rect 15654 41460 15660 41472
rect 15436 41432 15660 41460
rect 15436 41420 15442 41432
rect 15654 41420 15660 41432
rect 15712 41420 15718 41472
rect 17586 41420 17592 41472
rect 17644 41460 17650 41472
rect 20530 41460 20536 41472
rect 17644 41432 20536 41460
rect 17644 41420 17650 41432
rect 20530 41420 20536 41432
rect 20588 41420 20594 41472
rect 23474 41420 23480 41472
rect 23532 41420 23538 41472
rect 23750 41420 23756 41472
rect 23808 41460 23814 41472
rect 24578 41460 24584 41472
rect 23808 41432 24584 41460
rect 23808 41420 23814 41432
rect 24578 41420 24584 41432
rect 24636 41420 24642 41472
rect 27798 41420 27804 41472
rect 27856 41420 27862 41472
rect 552 41370 31648 41392
rect 552 41318 3662 41370
rect 3714 41318 3726 41370
rect 3778 41318 3790 41370
rect 3842 41318 3854 41370
rect 3906 41318 3918 41370
rect 3970 41318 11436 41370
rect 11488 41318 11500 41370
rect 11552 41318 11564 41370
rect 11616 41318 11628 41370
rect 11680 41318 11692 41370
rect 11744 41318 19210 41370
rect 19262 41318 19274 41370
rect 19326 41318 19338 41370
rect 19390 41318 19402 41370
rect 19454 41318 19466 41370
rect 19518 41318 26984 41370
rect 27036 41318 27048 41370
rect 27100 41318 27112 41370
rect 27164 41318 27176 41370
rect 27228 41318 27240 41370
rect 27292 41318 31648 41370
rect 552 41296 31648 41318
rect 9674 41256 9680 41268
rect 8864 41228 9680 41256
rect 8294 41012 8300 41064
rect 8352 41052 8358 41064
rect 8864 41061 8892 41228
rect 9674 41216 9680 41228
rect 9732 41216 9738 41268
rect 10134 41216 10140 41268
rect 10192 41256 10198 41268
rect 10597 41259 10655 41265
rect 10597 41256 10609 41259
rect 10192 41228 10609 41256
rect 10192 41216 10198 41228
rect 10597 41225 10609 41228
rect 10643 41225 10655 41259
rect 12618 41256 12624 41268
rect 10597 41219 10655 41225
rect 10796 41228 12624 41256
rect 9214 41148 9220 41200
rect 9272 41188 9278 41200
rect 10796 41188 10824 41228
rect 12618 41216 12624 41228
rect 12676 41216 12682 41268
rect 15028 41228 15516 41256
rect 9272 41160 10824 41188
rect 9272 41148 9278 41160
rect 9140 41092 9444 41120
rect 8573 41055 8631 41061
rect 8573 41052 8585 41055
rect 8352 41024 8585 41052
rect 8352 41012 8358 41024
rect 8573 41021 8585 41024
rect 8619 41021 8631 41055
rect 8573 41015 8631 41021
rect 8849 41055 8907 41061
rect 8849 41021 8861 41055
rect 8895 41021 8907 41055
rect 8849 41015 8907 41021
rect 8588 40984 8616 41015
rect 8938 41012 8944 41064
rect 8996 41012 9002 41064
rect 9140 41061 9168 41092
rect 9125 41055 9183 41061
rect 9125 41021 9137 41055
rect 9171 41021 9183 41055
rect 9125 41015 9183 41021
rect 9214 41012 9220 41064
rect 9272 41012 9278 41064
rect 9416 41052 9444 41092
rect 9490 41080 9496 41132
rect 9548 41120 9554 41132
rect 9861 41123 9919 41129
rect 9861 41120 9873 41123
rect 9548 41092 9873 41120
rect 9548 41080 9554 41092
rect 9861 41089 9873 41092
rect 9907 41089 9919 41123
rect 10594 41120 10600 41132
rect 9861 41083 9919 41089
rect 10060 41092 10600 41120
rect 9766 41052 9772 41064
rect 9416 41024 9772 41052
rect 9766 41012 9772 41024
rect 9824 41012 9830 41064
rect 10060 41061 10088 41092
rect 10594 41080 10600 41092
rect 10652 41080 10658 41132
rect 10778 41080 10784 41132
rect 10836 41120 10842 41132
rect 10836 41092 11468 41120
rect 10836 41080 10842 41092
rect 10045 41055 10103 41061
rect 10045 41021 10057 41055
rect 10091 41021 10103 41055
rect 10045 41015 10103 41021
rect 10134 41012 10140 41064
rect 10192 41012 10198 41064
rect 10318 41012 10324 41064
rect 10376 41012 10382 41064
rect 10413 41055 10471 41061
rect 10413 41021 10425 41055
rect 10459 41052 10471 41055
rect 10962 41052 10968 41064
rect 10459 41024 10968 41052
rect 10459 41021 10471 41024
rect 10413 41015 10471 41021
rect 10962 41012 10968 41024
rect 11020 41012 11026 41064
rect 11054 41012 11060 41064
rect 11112 41012 11118 41064
rect 11149 41055 11207 41061
rect 11149 41021 11161 41055
rect 11195 41052 11207 41055
rect 11333 41055 11391 41061
rect 11333 41052 11345 41055
rect 11195 41024 11345 41052
rect 11195 41021 11207 41024
rect 11149 41015 11207 41021
rect 11333 41021 11345 41024
rect 11379 41021 11391 41055
rect 11440 41052 11468 41092
rect 14369 41055 14427 41061
rect 11440 41024 13216 41052
rect 11333 41015 11391 41021
rect 11072 40984 11100 41012
rect 8588 40956 11100 40984
rect 11600 40987 11658 40993
rect 11600 40953 11612 40987
rect 11646 40984 11658 40987
rect 11790 40984 11796 40996
rect 11646 40956 11796 40984
rect 11646 40953 11658 40956
rect 11600 40947 11658 40953
rect 11790 40944 11796 40956
rect 11848 40944 11854 40996
rect 8110 40876 8116 40928
rect 8168 40916 8174 40928
rect 8481 40919 8539 40925
rect 8481 40916 8493 40919
rect 8168 40888 8493 40916
rect 8168 40876 8174 40888
rect 8481 40885 8493 40888
rect 8527 40885 8539 40919
rect 8481 40879 8539 40885
rect 8662 40876 8668 40928
rect 8720 40876 8726 40928
rect 9122 40876 9128 40928
rect 9180 40916 9186 40928
rect 9309 40919 9367 40925
rect 9309 40916 9321 40919
rect 9180 40888 9321 40916
rect 9180 40876 9186 40888
rect 9309 40885 9321 40888
rect 9355 40885 9367 40919
rect 12406 40916 12434 41024
rect 12802 40944 12808 40996
rect 12860 40944 12866 40996
rect 12989 40987 13047 40993
rect 12989 40953 13001 40987
rect 13035 40984 13047 40987
rect 13078 40984 13084 40996
rect 13035 40956 13084 40984
rect 13035 40953 13047 40956
rect 12989 40947 13047 40953
rect 12526 40916 12532 40928
rect 12406 40888 12532 40916
rect 9309 40879 9367 40885
rect 12526 40876 12532 40888
rect 12584 40876 12590 40928
rect 12710 40876 12716 40928
rect 12768 40916 12774 40928
rect 13004 40916 13032 40947
rect 13078 40944 13084 40956
rect 13136 40944 13142 40996
rect 13188 40984 13216 41024
rect 14369 41021 14381 41055
rect 14415 41052 14427 41055
rect 15028 41052 15056 41228
rect 15194 41148 15200 41200
rect 15252 41148 15258 41200
rect 15488 41188 15516 41228
rect 15562 41216 15568 41268
rect 15620 41216 15626 41268
rect 16482 41256 16488 41268
rect 15764 41228 16488 41256
rect 15764 41188 15792 41228
rect 16482 41216 16488 41228
rect 16540 41216 16546 41268
rect 17310 41216 17316 41268
rect 17368 41256 17374 41268
rect 17957 41259 18015 41265
rect 17957 41256 17969 41259
rect 17368 41228 17969 41256
rect 17368 41216 17374 41228
rect 17957 41225 17969 41228
rect 18003 41225 18015 41259
rect 17957 41219 18015 41225
rect 18138 41216 18144 41268
rect 18196 41256 18202 41268
rect 19058 41256 19064 41268
rect 18196 41228 19064 41256
rect 18196 41216 18202 41228
rect 19058 41216 19064 41228
rect 19116 41216 19122 41268
rect 19521 41259 19579 41265
rect 19521 41225 19533 41259
rect 19567 41256 19579 41259
rect 20346 41256 20352 41268
rect 19567 41228 20352 41256
rect 19567 41225 19579 41228
rect 19521 41219 19579 41225
rect 20346 41216 20352 41228
rect 20404 41216 20410 41268
rect 20809 41259 20867 41265
rect 20809 41225 20821 41259
rect 20855 41256 20867 41259
rect 21358 41256 21364 41268
rect 20855 41228 21364 41256
rect 20855 41225 20867 41228
rect 20809 41219 20867 41225
rect 21358 41216 21364 41228
rect 21416 41216 21422 41268
rect 22646 41216 22652 41268
rect 22704 41256 22710 41268
rect 22833 41259 22891 41265
rect 22833 41256 22845 41259
rect 22704 41228 22845 41256
rect 22704 41216 22710 41228
rect 22833 41225 22845 41228
rect 22879 41225 22891 41259
rect 22833 41219 22891 41225
rect 26602 41216 26608 41268
rect 26660 41256 26666 41268
rect 26789 41259 26847 41265
rect 26789 41256 26801 41259
rect 26660 41228 26801 41256
rect 26660 41216 26666 41228
rect 26789 41225 26801 41228
rect 26835 41225 26847 41259
rect 26789 41219 26847 41225
rect 28166 41216 28172 41268
rect 28224 41216 28230 41268
rect 28813 41259 28871 41265
rect 28813 41225 28825 41259
rect 28859 41256 28871 41259
rect 29454 41256 29460 41268
rect 28859 41228 29460 41256
rect 28859 41225 28871 41228
rect 28813 41219 28871 41225
rect 29454 41216 29460 41228
rect 29512 41216 29518 41268
rect 26237 41191 26295 41197
rect 15488 41160 15792 41188
rect 15856 41160 20300 41188
rect 15212 41120 15240 41148
rect 15212 41092 15516 41120
rect 14415 41024 15056 41052
rect 14415 41021 14427 41024
rect 14369 41015 14427 41021
rect 15102 41012 15108 41064
rect 15160 41012 15166 41064
rect 15194 41012 15200 41064
rect 15252 41012 15258 41064
rect 15289 41055 15347 41061
rect 15289 41021 15301 41055
rect 15335 41052 15347 41055
rect 15378 41052 15384 41064
rect 15335 41024 15384 41052
rect 15335 41021 15347 41024
rect 15289 41015 15347 41021
rect 15378 41012 15384 41024
rect 15436 41012 15442 41064
rect 15488 41061 15516 41092
rect 15473 41055 15531 41061
rect 15473 41021 15485 41055
rect 15519 41021 15531 41055
rect 15473 41015 15531 41021
rect 15488 40984 15516 41015
rect 15562 41012 15568 41064
rect 15620 41052 15626 41064
rect 15856 41061 15884 41160
rect 17126 41120 17132 41132
rect 16592 41092 17132 41120
rect 15749 41055 15807 41061
rect 15749 41052 15761 41055
rect 15620 41024 15761 41052
rect 15620 41012 15626 41024
rect 15749 41021 15761 41024
rect 15795 41021 15807 41055
rect 15749 41015 15807 41021
rect 15841 41055 15899 41061
rect 15841 41021 15853 41055
rect 15887 41021 15899 41055
rect 15841 41015 15899 41021
rect 13188 40956 15516 40984
rect 15764 40984 15792 41015
rect 15930 41012 15936 41064
rect 15988 41052 15994 41064
rect 16025 41055 16083 41061
rect 16025 41052 16037 41055
rect 15988 41024 16037 41052
rect 15988 41012 15994 41024
rect 16025 41021 16037 41024
rect 16071 41021 16083 41055
rect 16025 41015 16083 41021
rect 16114 41012 16120 41064
rect 16172 41012 16178 41064
rect 16298 41012 16304 41064
rect 16356 41052 16362 41064
rect 16592 41061 16620 41092
rect 17126 41080 17132 41092
rect 17184 41080 17190 41132
rect 17586 41080 17592 41132
rect 17644 41120 17650 41132
rect 20272 41120 20300 41160
rect 26237 41157 26249 41191
rect 26283 41157 26295 41191
rect 26237 41151 26295 41157
rect 23474 41120 23480 41132
rect 17644 41092 17724 41120
rect 17644 41080 17650 41092
rect 16577 41055 16635 41061
rect 16356 41024 16528 41052
rect 16356 41012 16362 41024
rect 16209 40987 16267 40993
rect 16209 40984 16221 40987
rect 15764 40956 16221 40984
rect 15212 40928 15240 40956
rect 16209 40953 16221 40956
rect 16255 40953 16267 40987
rect 16209 40947 16267 40953
rect 16393 40987 16451 40993
rect 16393 40953 16405 40987
rect 16439 40953 16451 40987
rect 16500 40984 16528 41024
rect 16577 41021 16589 41055
rect 16623 41021 16635 41055
rect 16577 41015 16635 41021
rect 16761 41055 16819 41061
rect 16761 41021 16773 41055
rect 16807 41052 16819 41055
rect 17034 41052 17040 41064
rect 16807 41024 17040 41052
rect 16807 41021 16819 41024
rect 16761 41015 16819 41021
rect 17034 41012 17040 41024
rect 17092 41012 17098 41064
rect 17696 41061 17724 41092
rect 17788 41092 19840 41120
rect 20272 41092 23480 41120
rect 17313 41055 17371 41061
rect 17313 41021 17325 41055
rect 17359 41021 17371 41055
rect 17313 41015 17371 41021
rect 17681 41055 17739 41061
rect 17681 41021 17693 41055
rect 17727 41021 17739 41055
rect 17681 41015 17739 41021
rect 17328 40984 17356 41015
rect 16500 40956 17356 40984
rect 16393 40947 16451 40953
rect 12768 40888 13032 40916
rect 13173 40919 13231 40925
rect 12768 40876 12774 40888
rect 13173 40885 13185 40919
rect 13219 40916 13231 40919
rect 13262 40916 13268 40928
rect 13219 40888 13268 40916
rect 13219 40885 13231 40888
rect 13173 40879 13231 40885
rect 13262 40876 13268 40888
rect 13320 40876 13326 40928
rect 14090 40876 14096 40928
rect 14148 40916 14154 40928
rect 14277 40919 14335 40925
rect 14277 40916 14289 40919
rect 14148 40888 14289 40916
rect 14148 40876 14154 40888
rect 14277 40885 14289 40888
rect 14323 40885 14335 40919
rect 14277 40879 14335 40885
rect 14366 40876 14372 40928
rect 14424 40916 14430 40928
rect 14829 40919 14887 40925
rect 14829 40916 14841 40919
rect 14424 40888 14841 40916
rect 14424 40876 14430 40888
rect 14829 40885 14841 40888
rect 14875 40885 14887 40919
rect 14829 40879 14887 40885
rect 15194 40876 15200 40928
rect 15252 40876 15258 40928
rect 15286 40876 15292 40928
rect 15344 40916 15350 40928
rect 16408 40916 16436 40947
rect 17402 40944 17408 40996
rect 17460 40984 17466 40996
rect 17497 40987 17555 40993
rect 17497 40984 17509 40987
rect 17460 40956 17509 40984
rect 17460 40944 17466 40956
rect 17497 40953 17509 40956
rect 17543 40953 17555 40987
rect 17497 40947 17555 40953
rect 17586 40944 17592 40996
rect 17644 40944 17650 40996
rect 15344 40888 16436 40916
rect 15344 40876 15350 40888
rect 16666 40876 16672 40928
rect 16724 40876 16730 40928
rect 17310 40876 17316 40928
rect 17368 40916 17374 40928
rect 17788 40916 17816 41092
rect 17862 41012 17868 41064
rect 17920 41012 17926 41064
rect 17954 41012 17960 41064
rect 18012 41052 18018 41064
rect 18141 41055 18199 41061
rect 18141 41052 18153 41055
rect 18012 41024 18153 41052
rect 18012 41012 18018 41024
rect 18141 41021 18153 41024
rect 18187 41021 18199 41055
rect 18141 41015 18199 41021
rect 18509 41055 18567 41061
rect 18509 41021 18521 41055
rect 18555 41052 18567 41055
rect 19334 41052 19340 41064
rect 18555 41024 19340 41052
rect 18555 41021 18567 41024
rect 18509 41015 18567 41021
rect 19334 41012 19340 41024
rect 19392 41012 19398 41064
rect 19429 41055 19487 41061
rect 19429 41021 19441 41055
rect 19475 41052 19487 41055
rect 19518 41052 19524 41064
rect 19475 41024 19524 41052
rect 19475 41021 19487 41024
rect 19429 41015 19487 41021
rect 19518 41012 19524 41024
rect 19576 41012 19582 41064
rect 19613 41055 19671 41061
rect 19613 41021 19625 41055
rect 19659 41052 19671 41055
rect 19702 41052 19708 41064
rect 19659 41024 19708 41052
rect 19659 41021 19671 41024
rect 19613 41015 19671 41021
rect 19702 41012 19708 41024
rect 19760 41012 19766 41064
rect 19812 41061 19840 41092
rect 23474 41080 23480 41092
rect 23532 41080 23538 41132
rect 26252 41120 26280 41151
rect 26326 41148 26332 41200
rect 26384 41188 26390 41200
rect 26384 41160 28304 41188
rect 26384 41148 26390 41160
rect 25240 41092 26280 41120
rect 26605 41123 26663 41129
rect 19797 41055 19855 41061
rect 19797 41021 19809 41055
rect 19843 41021 19855 41055
rect 19797 41015 19855 41021
rect 19981 41055 20039 41061
rect 19981 41021 19993 41055
rect 20027 41021 20039 41055
rect 19981 41015 20039 41021
rect 20165 41055 20223 41061
rect 20165 41021 20177 41055
rect 20211 41052 20223 41055
rect 20254 41052 20260 41064
rect 20211 41024 20260 41052
rect 20211 41021 20223 41024
rect 20165 41015 20223 41021
rect 17880 40984 17908 41012
rect 19242 40984 19248 40996
rect 17880 40956 19248 40984
rect 19242 40944 19248 40956
rect 19300 40944 19306 40996
rect 19720 40984 19748 41012
rect 19996 40984 20024 41015
rect 20254 41012 20260 41024
rect 20312 41012 20318 41064
rect 20346 41012 20352 41064
rect 20404 41012 20410 41064
rect 20438 41012 20444 41064
rect 20496 41012 20502 41064
rect 20533 41055 20591 41061
rect 20533 41021 20545 41055
rect 20579 41021 20591 41055
rect 22094 41052 22100 41064
rect 20533 41015 20591 41021
rect 19720 40956 20024 40984
rect 20070 40944 20076 40996
rect 20128 40944 20134 40996
rect 20548 40984 20576 41015
rect 22066 41012 22100 41052
rect 22152 41012 22158 41064
rect 22189 41055 22247 41061
rect 22189 41021 22201 41055
rect 22235 41052 22247 41055
rect 22370 41052 22376 41064
rect 22235 41024 22376 41052
rect 22235 41021 22247 41024
rect 22189 41015 22247 41021
rect 22370 41012 22376 41024
rect 22428 41012 22434 41064
rect 22741 41055 22799 41061
rect 22741 41021 22753 41055
rect 22787 41052 22799 41055
rect 23750 41052 23756 41064
rect 22787 41024 23756 41052
rect 22787 41021 22799 41024
rect 22741 41015 22799 41021
rect 22066 40984 22094 41012
rect 22756 40984 22784 41015
rect 23750 41012 23756 41024
rect 23808 41012 23814 41064
rect 23934 41012 23940 41064
rect 23992 41012 23998 41064
rect 24204 41055 24262 41061
rect 24204 41021 24216 41055
rect 24250 41052 24262 41055
rect 25240 41052 25268 41092
rect 26605 41089 26617 41123
rect 26651 41120 26663 41123
rect 26651 41092 26740 41120
rect 26651 41089 26663 41092
rect 26605 41083 26663 41089
rect 24250 41024 25268 41052
rect 24250 41021 24262 41024
rect 24204 41015 24262 41021
rect 25314 41012 25320 41064
rect 25372 41052 25378 41064
rect 26053 41055 26111 41061
rect 26053 41052 26065 41055
rect 25372 41024 26065 41052
rect 25372 41012 25378 41024
rect 26053 41021 26065 41024
rect 26099 41021 26111 41055
rect 26053 41015 26111 41021
rect 26142 41012 26148 41064
rect 26200 41052 26206 41064
rect 26513 41055 26571 41061
rect 26513 41052 26525 41055
rect 26200 41024 26525 41052
rect 26200 41012 26206 41024
rect 26513 41021 26525 41024
rect 26559 41021 26571 41055
rect 26513 41015 26571 41021
rect 20364 40956 22784 40984
rect 23385 40987 23443 40993
rect 17368 40888 17816 40916
rect 17865 40919 17923 40925
rect 17368 40876 17374 40888
rect 17865 40885 17877 40919
rect 17911 40916 17923 40919
rect 18046 40916 18052 40928
rect 17911 40888 18052 40916
rect 17911 40885 17923 40888
rect 17865 40879 17923 40885
rect 18046 40876 18052 40888
rect 18104 40876 18110 40928
rect 19981 40919 20039 40925
rect 19981 40885 19993 40919
rect 20027 40916 20039 40919
rect 20088 40916 20116 40944
rect 20364 40928 20392 40956
rect 23385 40953 23397 40987
rect 23431 40984 23443 40987
rect 23474 40984 23480 40996
rect 23431 40956 23480 40984
rect 23431 40953 23443 40956
rect 23385 40947 23443 40953
rect 23474 40944 23480 40956
rect 23532 40984 23538 40996
rect 24670 40984 24676 40996
rect 23532 40956 24676 40984
rect 23532 40944 23538 40956
rect 24670 40944 24676 40956
rect 24728 40944 24734 40996
rect 24854 40944 24860 40996
rect 24912 40984 24918 40996
rect 26237 40987 26295 40993
rect 26237 40984 26249 40987
rect 24912 40956 26249 40984
rect 24912 40944 24918 40956
rect 26237 40953 26249 40956
rect 26283 40953 26295 40987
rect 26712 40984 26740 41092
rect 26786 41080 26792 41132
rect 26844 41120 26850 41132
rect 27709 41123 27767 41129
rect 27709 41120 27721 41123
rect 26844 41092 27721 41120
rect 26844 41080 26850 41092
rect 27709 41089 27721 41092
rect 27755 41120 27767 41123
rect 27798 41120 27804 41132
rect 27755 41092 27804 41120
rect 27755 41089 27767 41092
rect 27709 41083 27767 41089
rect 27798 41080 27804 41092
rect 27856 41080 27862 41132
rect 28276 41129 28304 41160
rect 28261 41123 28319 41129
rect 28261 41089 28273 41123
rect 28307 41089 28319 41123
rect 28902 41120 28908 41132
rect 28261 41083 28319 41089
rect 28368 41092 28908 41120
rect 26881 41055 26939 41061
rect 26881 41021 26893 41055
rect 26927 41052 26939 41055
rect 27157 41055 27215 41061
rect 27157 41052 27169 41055
rect 26927 41024 27169 41052
rect 26927 41021 26939 41024
rect 26881 41015 26939 41021
rect 27157 41021 27169 41024
rect 27203 41021 27215 41055
rect 27157 41015 27215 41021
rect 27893 41055 27951 41061
rect 27893 41021 27905 41055
rect 27939 41021 27951 41055
rect 27893 41015 27951 41021
rect 27985 41055 28043 41061
rect 27985 41021 27997 41055
rect 28031 41052 28043 41055
rect 28368 41052 28396 41092
rect 28552 41061 28580 41092
rect 28902 41080 28908 41092
rect 28960 41080 28966 41132
rect 28997 41123 29055 41129
rect 28997 41089 29009 41123
rect 29043 41120 29055 41123
rect 29546 41120 29552 41132
rect 29043 41092 29552 41120
rect 29043 41089 29055 41092
rect 28997 41083 29055 41089
rect 29546 41080 29552 41092
rect 29604 41080 29610 41132
rect 28031 41024 28396 41052
rect 28445 41055 28503 41061
rect 28031 41021 28043 41024
rect 27985 41015 28043 41021
rect 28445 41021 28457 41055
rect 28491 41021 28503 41055
rect 28445 41015 28503 41021
rect 28537 41055 28595 41061
rect 28537 41021 28549 41055
rect 28583 41021 28595 41055
rect 28537 41015 28595 41021
rect 27430 40984 27436 40996
rect 26712 40956 27436 40984
rect 26237 40947 26295 40953
rect 27430 40944 27436 40956
rect 27488 40944 27494 40996
rect 27908 40984 27936 41015
rect 28169 40987 28227 40993
rect 27908 40956 28028 40984
rect 20027 40888 20116 40916
rect 20027 40885 20039 40888
rect 19981 40879 20039 40885
rect 20346 40876 20352 40928
rect 20404 40876 20410 40928
rect 21910 40876 21916 40928
rect 21968 40916 21974 40928
rect 22097 40919 22155 40925
rect 22097 40916 22109 40919
rect 21968 40888 22109 40916
rect 21968 40876 21974 40888
rect 22097 40885 22109 40888
rect 22143 40885 22155 40919
rect 22097 40879 22155 40885
rect 23290 40876 23296 40928
rect 23348 40876 23354 40928
rect 25222 40876 25228 40928
rect 25280 40916 25286 40928
rect 25317 40919 25375 40925
rect 25317 40916 25329 40919
rect 25280 40888 25329 40916
rect 25280 40876 25286 40888
rect 25317 40885 25329 40888
rect 25363 40885 25375 40919
rect 25317 40879 25375 40885
rect 25498 40876 25504 40928
rect 25556 40916 25562 40928
rect 26421 40919 26479 40925
rect 26421 40916 26433 40919
rect 25556 40888 26433 40916
rect 25556 40876 25562 40888
rect 26421 40885 26433 40888
rect 26467 40885 26479 40919
rect 26421 40879 26479 40885
rect 26510 40876 26516 40928
rect 26568 40916 26574 40928
rect 26605 40919 26663 40925
rect 26605 40916 26617 40919
rect 26568 40888 26617 40916
rect 26568 40876 26574 40888
rect 26605 40885 26617 40888
rect 26651 40885 26663 40919
rect 28000 40916 28028 40956
rect 28169 40953 28181 40987
rect 28215 40984 28227 40987
rect 28261 40987 28319 40993
rect 28261 40984 28273 40987
rect 28215 40956 28273 40984
rect 28215 40953 28227 40956
rect 28169 40947 28227 40953
rect 28261 40953 28273 40956
rect 28307 40953 28319 40987
rect 28261 40947 28319 40953
rect 28460 40984 28488 41015
rect 28626 41012 28632 41064
rect 28684 41012 28690 41064
rect 28813 41055 28871 41061
rect 28813 41021 28825 41055
rect 28859 41021 28871 41055
rect 28813 41015 28871 41021
rect 29181 41055 29239 41061
rect 29181 41021 29193 41055
rect 29227 41021 29239 41055
rect 29181 41015 29239 41021
rect 28644 40984 28672 41012
rect 28460 40956 28672 40984
rect 28828 40984 28856 41015
rect 28997 40987 29055 40993
rect 28997 40984 29009 40987
rect 28828 40956 29009 40984
rect 28460 40916 28488 40956
rect 28997 40953 29009 40956
rect 29043 40953 29055 40987
rect 28997 40947 29055 40953
rect 29196 40984 29224 41015
rect 29270 41012 29276 41064
rect 29328 41012 29334 41064
rect 30837 41055 30895 41061
rect 30837 41021 30849 41055
rect 30883 41052 30895 41055
rect 31110 41052 31116 41064
rect 30883 41024 31116 41052
rect 30883 41021 30895 41024
rect 30837 41015 30895 41021
rect 31110 41012 31116 41024
rect 31168 41012 31174 41064
rect 30592 40987 30650 40993
rect 29196 40956 29592 40984
rect 28000 40888 28488 40916
rect 26605 40879 26663 40885
rect 28534 40876 28540 40928
rect 28592 40916 28598 40928
rect 29196 40916 29224 40956
rect 28592 40888 29224 40916
rect 28592 40876 28598 40888
rect 29454 40876 29460 40928
rect 29512 40876 29518 40928
rect 29564 40916 29592 40956
rect 30592 40953 30604 40987
rect 30638 40984 30650 40987
rect 30742 40984 30748 40996
rect 30638 40956 30748 40984
rect 30638 40953 30650 40956
rect 30592 40947 30650 40953
rect 30742 40944 30748 40956
rect 30800 40944 30806 40996
rect 30926 40916 30932 40928
rect 29564 40888 30932 40916
rect 30926 40876 30932 40888
rect 30984 40876 30990 40928
rect 552 40826 31648 40848
rect 552 40774 4322 40826
rect 4374 40774 4386 40826
rect 4438 40774 4450 40826
rect 4502 40774 4514 40826
rect 4566 40774 4578 40826
rect 4630 40774 12096 40826
rect 12148 40774 12160 40826
rect 12212 40774 12224 40826
rect 12276 40774 12288 40826
rect 12340 40774 12352 40826
rect 12404 40774 19870 40826
rect 19922 40774 19934 40826
rect 19986 40774 19998 40826
rect 20050 40774 20062 40826
rect 20114 40774 20126 40826
rect 20178 40774 27644 40826
rect 27696 40774 27708 40826
rect 27760 40774 27772 40826
rect 27824 40774 27836 40826
rect 27888 40774 27900 40826
rect 27952 40774 31648 40826
rect 552 40752 31648 40774
rect 10134 40672 10140 40724
rect 10192 40712 10198 40724
rect 10781 40715 10839 40721
rect 10781 40712 10793 40715
rect 10192 40684 10793 40712
rect 10192 40672 10198 40684
rect 10781 40681 10793 40684
rect 10827 40681 10839 40715
rect 10781 40675 10839 40681
rect 10962 40672 10968 40724
rect 11020 40672 11026 40724
rect 11790 40672 11796 40724
rect 11848 40672 11854 40724
rect 12434 40712 12440 40724
rect 12084 40684 12440 40712
rect 8938 40604 8944 40656
rect 8996 40644 9002 40656
rect 10226 40644 10232 40656
rect 8996 40616 10232 40644
rect 8996 40604 9002 40616
rect 10226 40604 10232 40616
rect 10284 40604 10290 40656
rect 11974 40644 11980 40656
rect 10428 40616 11980 40644
rect 8110 40536 8116 40588
rect 8168 40536 8174 40588
rect 8380 40579 8438 40585
rect 8380 40545 8392 40579
rect 8426 40576 8438 40579
rect 8846 40576 8852 40588
rect 8426 40548 8852 40576
rect 8426 40545 8438 40548
rect 8380 40539 8438 40545
rect 8846 40536 8852 40548
rect 8904 40536 8910 40588
rect 9582 40536 9588 40588
rect 9640 40576 9646 40588
rect 10428 40585 10456 40616
rect 11974 40604 11980 40616
rect 12032 40604 12038 40656
rect 12084 40585 12112 40684
rect 12434 40672 12440 40684
rect 12492 40672 12498 40724
rect 15102 40672 15108 40724
rect 15160 40712 15166 40724
rect 15473 40715 15531 40721
rect 15473 40712 15485 40715
rect 15160 40684 15485 40712
rect 15160 40672 15166 40684
rect 15473 40681 15485 40684
rect 15519 40681 15531 40715
rect 15473 40675 15531 40681
rect 12710 40644 12716 40656
rect 12360 40616 12716 40644
rect 9677 40579 9735 40585
rect 9677 40576 9689 40579
rect 9640 40548 9689 40576
rect 9640 40536 9646 40548
rect 9677 40545 9689 40548
rect 9723 40545 9735 40579
rect 9677 40539 9735 40545
rect 9861 40579 9919 40585
rect 9861 40545 9873 40579
rect 9907 40545 9919 40579
rect 9861 40539 9919 40545
rect 10045 40579 10103 40585
rect 10045 40545 10057 40579
rect 10091 40576 10103 40579
rect 10137 40579 10195 40585
rect 10137 40576 10149 40579
rect 10091 40548 10149 40576
rect 10091 40545 10103 40548
rect 10045 40539 10103 40545
rect 10137 40545 10149 40548
rect 10183 40545 10195 40579
rect 10137 40539 10195 40545
rect 10321 40579 10379 40585
rect 10321 40545 10333 40579
rect 10367 40545 10379 40579
rect 10321 40539 10379 40545
rect 10413 40579 10471 40585
rect 10413 40545 10425 40579
rect 10459 40545 10471 40579
rect 10413 40539 10471 40545
rect 10505 40579 10563 40585
rect 10505 40545 10517 40579
rect 10551 40576 10563 40579
rect 11333 40579 11391 40585
rect 11333 40576 11345 40579
rect 10551 40548 11345 40576
rect 10551 40545 10563 40548
rect 10505 40539 10563 40545
rect 11333 40545 11345 40548
rect 11379 40576 11391 40579
rect 12069 40579 12127 40585
rect 11379 40548 11652 40576
rect 11379 40545 11391 40548
rect 11333 40539 11391 40545
rect 9876 40508 9904 40539
rect 9508 40480 9904 40508
rect 9508 40384 9536 40480
rect 9858 40400 9864 40452
rect 9916 40440 9922 40452
rect 10336 40440 10364 40539
rect 10686 40468 10692 40520
rect 10744 40508 10750 40520
rect 11425 40511 11483 40517
rect 11425 40508 11437 40511
rect 10744 40480 11437 40508
rect 10744 40468 10750 40480
rect 11425 40477 11437 40480
rect 11471 40477 11483 40511
rect 11425 40471 11483 40477
rect 11517 40511 11575 40517
rect 11517 40477 11529 40511
rect 11563 40477 11575 40511
rect 11624 40508 11652 40548
rect 12069 40545 12081 40579
rect 12115 40545 12127 40579
rect 12069 40539 12127 40545
rect 12158 40536 12164 40588
rect 12216 40536 12222 40588
rect 12250 40536 12256 40588
rect 12308 40536 12314 40588
rect 12360 40508 12388 40616
rect 12710 40604 12716 40616
rect 12768 40604 12774 40656
rect 15488 40644 15516 40675
rect 16758 40672 16764 40724
rect 16816 40712 16822 40724
rect 17218 40712 17224 40724
rect 16816 40684 17224 40712
rect 16816 40672 16822 40684
rect 17218 40672 17224 40684
rect 17276 40672 17282 40724
rect 17402 40672 17408 40724
rect 17460 40712 17466 40724
rect 17460 40684 18460 40712
rect 17460 40672 17466 40684
rect 18432 40656 18460 40684
rect 19242 40672 19248 40724
rect 19300 40712 19306 40724
rect 20346 40712 20352 40724
rect 19300 40684 20352 40712
rect 19300 40672 19306 40684
rect 20346 40672 20352 40684
rect 20404 40672 20410 40724
rect 23198 40672 23204 40724
rect 23256 40712 23262 40724
rect 23293 40715 23351 40721
rect 23293 40712 23305 40715
rect 23256 40684 23305 40712
rect 23256 40672 23262 40684
rect 23293 40681 23305 40684
rect 23339 40681 23351 40715
rect 23293 40675 23351 40681
rect 23934 40672 23940 40724
rect 23992 40712 23998 40724
rect 24121 40715 24179 40721
rect 24121 40712 24133 40715
rect 23992 40684 24133 40712
rect 23992 40672 23998 40684
rect 24121 40681 24133 40684
rect 24167 40681 24179 40715
rect 24121 40675 24179 40681
rect 24854 40672 24860 40724
rect 24912 40672 24918 40724
rect 25961 40715 26019 40721
rect 25961 40681 25973 40715
rect 26007 40712 26019 40715
rect 26694 40712 26700 40724
rect 26007 40684 26700 40712
rect 26007 40681 26019 40684
rect 25961 40675 26019 40681
rect 26694 40672 26700 40684
rect 26752 40672 26758 40724
rect 30742 40672 30748 40724
rect 30800 40712 30806 40724
rect 30837 40715 30895 40721
rect 30837 40712 30849 40715
rect 30800 40684 30849 40712
rect 30800 40672 30806 40684
rect 30837 40681 30849 40684
rect 30883 40681 30895 40715
rect 30837 40675 30895 40681
rect 31110 40672 31116 40724
rect 31168 40672 31174 40724
rect 17586 40644 17592 40656
rect 15488 40616 17592 40644
rect 12431 40579 12489 40585
rect 12431 40545 12443 40579
rect 12477 40576 12489 40579
rect 12526 40576 12532 40588
rect 12477 40548 12532 40576
rect 12477 40545 12489 40548
rect 12431 40539 12489 40545
rect 12526 40536 12532 40548
rect 12584 40536 12590 40588
rect 12894 40536 12900 40588
rect 12952 40536 12958 40588
rect 12986 40536 12992 40588
rect 13044 40536 13050 40588
rect 13081 40579 13139 40585
rect 13081 40545 13093 40579
rect 13127 40545 13139 40579
rect 13081 40539 13139 40545
rect 11624 40480 12388 40508
rect 11517 40471 11575 40477
rect 9916 40412 10364 40440
rect 9916 40400 9922 40412
rect 10962 40400 10968 40452
rect 11020 40440 11026 40452
rect 11532 40440 11560 40471
rect 11020 40412 11560 40440
rect 11020 40400 11026 40412
rect 11790 40400 11796 40452
rect 11848 40440 11854 40452
rect 13096 40440 13124 40539
rect 13262 40536 13268 40588
rect 13320 40536 13326 40588
rect 14090 40536 14096 40588
rect 14148 40536 14154 40588
rect 14366 40536 14372 40588
rect 14424 40536 14430 40588
rect 16206 40536 16212 40588
rect 16264 40576 16270 40588
rect 16485 40579 16543 40585
rect 16485 40576 16497 40579
rect 16264 40548 16497 40576
rect 16264 40536 16270 40548
rect 16485 40545 16497 40548
rect 16531 40545 16543 40579
rect 16485 40539 16543 40545
rect 16758 40536 16764 40588
rect 16816 40536 16822 40588
rect 16945 40579 17003 40585
rect 16945 40545 16957 40579
rect 16991 40576 17003 40579
rect 16991 40548 17080 40576
rect 16991 40545 17003 40548
rect 16945 40539 17003 40545
rect 16577 40511 16635 40517
rect 16577 40477 16589 40511
rect 16623 40508 16635 40511
rect 16850 40508 16856 40520
rect 16623 40480 16856 40508
rect 16623 40477 16635 40480
rect 16577 40471 16635 40477
rect 16850 40468 16856 40480
rect 16908 40468 16914 40520
rect 17052 40517 17080 40548
rect 17126 40536 17132 40588
rect 17184 40576 17190 40588
rect 17512 40585 17540 40616
rect 17586 40604 17592 40616
rect 17644 40604 17650 40656
rect 17770 40604 17776 40656
rect 17828 40644 17834 40656
rect 18049 40647 18107 40653
rect 18049 40644 18061 40647
rect 17828 40616 18061 40644
rect 17828 40604 17834 40616
rect 18049 40613 18061 40616
rect 18095 40613 18107 40647
rect 18049 40607 18107 40613
rect 18414 40604 18420 40656
rect 18472 40644 18478 40656
rect 18598 40644 18604 40656
rect 18472 40616 18604 40644
rect 18472 40604 18478 40616
rect 18598 40604 18604 40616
rect 18656 40644 18662 40656
rect 19061 40647 19119 40653
rect 19061 40644 19073 40647
rect 18656 40616 19073 40644
rect 18656 40604 18662 40616
rect 19061 40613 19073 40616
rect 19107 40613 19119 40647
rect 19061 40607 19119 40613
rect 21450 40604 21456 40656
rect 21508 40604 21514 40656
rect 26234 40644 26240 40656
rect 24964 40616 26240 40644
rect 24964 40588 24992 40616
rect 26234 40604 26240 40616
rect 26292 40644 26298 40656
rect 27338 40644 27344 40656
rect 26292 40616 27344 40644
rect 26292 40604 26298 40616
rect 27338 40604 27344 40616
rect 27396 40604 27402 40656
rect 30653 40647 30711 40653
rect 30653 40613 30665 40647
rect 30699 40644 30711 40647
rect 30699 40616 30788 40644
rect 30699 40613 30711 40616
rect 30653 40607 30711 40613
rect 17497 40579 17555 40585
rect 17184 40548 17448 40576
rect 17184 40536 17190 40548
rect 17037 40511 17095 40517
rect 17037 40477 17049 40511
rect 17083 40477 17095 40511
rect 17037 40471 17095 40477
rect 17221 40511 17279 40517
rect 17221 40477 17233 40511
rect 17267 40477 17279 40511
rect 17221 40471 17279 40477
rect 14090 40440 14096 40452
rect 11848 40412 14096 40440
rect 11848 40400 11854 40412
rect 14090 40400 14096 40412
rect 14148 40400 14154 40452
rect 16669 40443 16727 40449
rect 16669 40409 16681 40443
rect 16715 40440 16727 40443
rect 16758 40440 16764 40452
rect 16715 40412 16764 40440
rect 16715 40409 16727 40412
rect 16669 40403 16727 40409
rect 16758 40400 16764 40412
rect 16816 40400 16822 40452
rect 17236 40440 17264 40471
rect 17310 40468 17316 40520
rect 17368 40468 17374 40520
rect 17420 40517 17448 40548
rect 17497 40545 17509 40579
rect 17543 40545 17555 40579
rect 17497 40539 17555 40545
rect 17681 40579 17739 40585
rect 17681 40545 17693 40579
rect 17727 40576 17739 40579
rect 17954 40576 17960 40588
rect 17727 40548 17960 40576
rect 17727 40545 17739 40548
rect 17681 40539 17739 40545
rect 17954 40536 17960 40548
rect 18012 40536 18018 40588
rect 18874 40536 18880 40588
rect 18932 40536 18938 40588
rect 19153 40579 19211 40585
rect 19153 40545 19165 40579
rect 19199 40576 19211 40579
rect 19334 40576 19340 40588
rect 19199 40548 19340 40576
rect 19199 40545 19211 40548
rect 19153 40539 19211 40545
rect 19334 40536 19340 40548
rect 19392 40576 19398 40588
rect 19610 40576 19616 40588
rect 19392 40548 19616 40576
rect 19392 40536 19398 40548
rect 19610 40536 19616 40548
rect 19668 40576 19674 40588
rect 19794 40576 19800 40588
rect 19668 40548 19800 40576
rect 19668 40536 19674 40548
rect 19794 40536 19800 40548
rect 19852 40536 19858 40588
rect 20714 40536 20720 40588
rect 20772 40576 20778 40588
rect 21269 40579 21327 40585
rect 21269 40576 21281 40579
rect 20772 40548 21281 40576
rect 20772 40536 20778 40548
rect 21269 40545 21281 40548
rect 21315 40545 21327 40579
rect 21269 40539 21327 40545
rect 21910 40536 21916 40588
rect 21968 40536 21974 40588
rect 22186 40585 22192 40588
rect 22180 40539 22192 40585
rect 22186 40536 22192 40539
rect 22244 40536 22250 40588
rect 23477 40579 23535 40585
rect 23477 40545 23489 40579
rect 23523 40576 23535 40579
rect 23566 40576 23572 40588
rect 23523 40548 23572 40576
rect 23523 40545 23535 40548
rect 23477 40539 23535 40545
rect 23566 40536 23572 40548
rect 23624 40536 23630 40588
rect 24213 40579 24271 40585
rect 24213 40545 24225 40579
rect 24259 40576 24271 40579
rect 24946 40576 24952 40588
rect 24259 40548 24952 40576
rect 24259 40545 24271 40548
rect 24213 40539 24271 40545
rect 24946 40536 24952 40548
rect 25004 40536 25010 40588
rect 25133 40579 25191 40585
rect 25133 40545 25145 40579
rect 25179 40576 25191 40579
rect 25498 40576 25504 40588
rect 25179 40548 25504 40576
rect 25179 40545 25191 40548
rect 25133 40539 25191 40545
rect 25498 40536 25504 40548
rect 25556 40536 25562 40588
rect 25869 40579 25927 40585
rect 25869 40545 25881 40579
rect 25915 40545 25927 40579
rect 25869 40539 25927 40545
rect 26053 40579 26111 40585
rect 26053 40545 26065 40579
rect 26099 40576 26111 40579
rect 26510 40576 26516 40588
rect 26099 40548 26516 40576
rect 26099 40545 26111 40548
rect 26053 40539 26111 40545
rect 17405 40511 17463 40517
rect 17405 40477 17417 40511
rect 17451 40508 17463 40511
rect 17865 40511 17923 40517
rect 17865 40508 17877 40511
rect 17451 40480 17877 40508
rect 17451 40477 17463 40480
rect 17405 40471 17463 40477
rect 17865 40477 17877 40480
rect 17911 40477 17923 40511
rect 17865 40471 17923 40477
rect 24857 40511 24915 40517
rect 24857 40477 24869 40511
rect 24903 40477 24915 40511
rect 24857 40471 24915 40477
rect 17236 40412 17448 40440
rect 17420 40384 17448 40412
rect 17678 40400 17684 40452
rect 17736 40440 17742 40452
rect 17880 40440 17908 40471
rect 17736 40412 17908 40440
rect 17979 40443 18037 40449
rect 17736 40400 17742 40412
rect 17979 40409 17991 40443
rect 18025 40440 18037 40443
rect 19058 40440 19064 40452
rect 18025 40412 19064 40440
rect 18025 40409 18037 40412
rect 17979 40403 18037 40409
rect 19058 40400 19064 40412
rect 19116 40400 19122 40452
rect 24872 40440 24900 40471
rect 25038 40468 25044 40520
rect 25096 40508 25102 40520
rect 25884 40508 25912 40539
rect 26510 40536 26516 40548
rect 26568 40536 26574 40588
rect 26602 40536 26608 40588
rect 26660 40536 26666 40588
rect 28350 40536 28356 40588
rect 28408 40536 28414 40588
rect 28445 40579 28503 40585
rect 28445 40545 28457 40579
rect 28491 40576 28503 40579
rect 28534 40576 28540 40588
rect 28491 40548 28540 40576
rect 28491 40545 28503 40548
rect 28445 40539 28503 40545
rect 28534 40536 28540 40548
rect 28592 40536 28598 40588
rect 29454 40536 29460 40588
rect 29512 40576 29518 40588
rect 30760 40585 30788 40616
rect 29641 40579 29699 40585
rect 29641 40576 29653 40579
rect 29512 40548 29653 40576
rect 29512 40536 29518 40548
rect 29641 40545 29653 40548
rect 29687 40545 29699 40579
rect 29641 40539 29699 40545
rect 30285 40579 30343 40585
rect 30285 40545 30297 40579
rect 30331 40576 30343 40579
rect 30377 40579 30435 40585
rect 30377 40576 30389 40579
rect 30331 40548 30389 40576
rect 30331 40545 30343 40548
rect 30285 40539 30343 40545
rect 30377 40545 30389 40548
rect 30423 40545 30435 40579
rect 30377 40539 30435 40545
rect 30745 40579 30803 40585
rect 30745 40545 30757 40579
rect 30791 40545 30803 40579
rect 30745 40539 30803 40545
rect 30926 40536 30932 40588
rect 30984 40536 30990 40588
rect 31018 40536 31024 40588
rect 31076 40536 31082 40588
rect 26142 40508 26148 40520
rect 25096 40480 26148 40508
rect 25096 40468 25102 40480
rect 26142 40468 26148 40480
rect 26200 40508 26206 40520
rect 26421 40511 26479 40517
rect 26421 40508 26433 40511
rect 26200 40480 26433 40508
rect 26200 40468 26206 40480
rect 26421 40477 26433 40480
rect 26467 40477 26479 40511
rect 26421 40471 26479 40477
rect 26786 40468 26792 40520
rect 26844 40468 26850 40520
rect 27430 40468 27436 40520
rect 27488 40508 27494 40520
rect 29546 40508 29552 40520
rect 27488 40480 29552 40508
rect 27488 40468 27494 40480
rect 29546 40468 29552 40480
rect 29604 40508 29610 40520
rect 30653 40511 30711 40517
rect 30653 40508 30665 40511
rect 29604 40480 30665 40508
rect 29604 40468 29610 40480
rect 30653 40477 30665 40480
rect 30699 40477 30711 40511
rect 30653 40471 30711 40477
rect 25130 40440 25136 40452
rect 24872 40412 25136 40440
rect 25130 40400 25136 40412
rect 25188 40400 25194 40452
rect 9490 40332 9496 40384
rect 9548 40372 9554 40384
rect 10686 40372 10692 40384
rect 9548 40344 10692 40372
rect 9548 40332 9554 40344
rect 10686 40332 10692 40344
rect 10744 40332 10750 40384
rect 12618 40332 12624 40384
rect 12676 40332 12682 40384
rect 15838 40332 15844 40384
rect 15896 40372 15902 40384
rect 16301 40375 16359 40381
rect 16301 40372 16313 40375
rect 15896 40344 16313 40372
rect 15896 40332 15902 40344
rect 16301 40341 16313 40344
rect 16347 40341 16359 40375
rect 16301 40335 16359 40341
rect 17402 40332 17408 40384
rect 17460 40332 17466 40384
rect 17494 40332 17500 40384
rect 17552 40372 17558 40384
rect 17773 40375 17831 40381
rect 17773 40372 17785 40375
rect 17552 40344 17785 40372
rect 17552 40332 17558 40344
rect 17773 40341 17785 40344
rect 17819 40341 17831 40375
rect 17773 40335 17831 40341
rect 18690 40332 18696 40384
rect 18748 40332 18754 40384
rect 21450 40332 21456 40384
rect 21508 40372 21514 40384
rect 21637 40375 21695 40381
rect 21637 40372 21649 40375
rect 21508 40344 21649 40372
rect 21508 40332 21514 40344
rect 21637 40341 21649 40344
rect 21683 40341 21695 40375
rect 21637 40335 21695 40341
rect 23474 40332 23480 40384
rect 23532 40372 23538 40384
rect 23569 40375 23627 40381
rect 23569 40372 23581 40375
rect 23532 40344 23581 40372
rect 23532 40332 23538 40344
rect 23569 40341 23581 40344
rect 23615 40341 23627 40375
rect 23569 40335 23627 40341
rect 28626 40332 28632 40384
rect 28684 40332 28690 40384
rect 30374 40332 30380 40384
rect 30432 40372 30438 40384
rect 30469 40375 30527 40381
rect 30469 40372 30481 40375
rect 30432 40344 30481 40372
rect 30432 40332 30438 40344
rect 30469 40341 30481 40344
rect 30515 40341 30527 40375
rect 30469 40335 30527 40341
rect 552 40282 31648 40304
rect 552 40230 3662 40282
rect 3714 40230 3726 40282
rect 3778 40230 3790 40282
rect 3842 40230 3854 40282
rect 3906 40230 3918 40282
rect 3970 40230 11436 40282
rect 11488 40230 11500 40282
rect 11552 40230 11564 40282
rect 11616 40230 11628 40282
rect 11680 40230 11692 40282
rect 11744 40230 19210 40282
rect 19262 40230 19274 40282
rect 19326 40230 19338 40282
rect 19390 40230 19402 40282
rect 19454 40230 19466 40282
rect 19518 40230 26984 40282
rect 27036 40230 27048 40282
rect 27100 40230 27112 40282
rect 27164 40230 27176 40282
rect 27228 40230 27240 40282
rect 27292 40230 31648 40282
rect 552 40208 31648 40230
rect 8846 40128 8852 40180
rect 8904 40128 8910 40180
rect 9674 40128 9680 40180
rect 9732 40128 9738 40180
rect 11149 40171 11207 40177
rect 11149 40137 11161 40171
rect 11195 40168 11207 40171
rect 12250 40168 12256 40180
rect 11195 40140 12256 40168
rect 11195 40137 11207 40140
rect 11149 40131 11207 40137
rect 12250 40128 12256 40140
rect 12308 40128 12314 40180
rect 15378 40128 15384 40180
rect 15436 40128 15442 40180
rect 16114 40128 16120 40180
rect 16172 40128 16178 40180
rect 16850 40128 16856 40180
rect 16908 40168 16914 40180
rect 17221 40171 17279 40177
rect 17221 40168 17233 40171
rect 16908 40140 17233 40168
rect 16908 40128 16914 40140
rect 17221 40137 17233 40140
rect 17267 40168 17279 40171
rect 17862 40168 17868 40180
rect 17267 40140 17868 40168
rect 17267 40137 17279 40140
rect 17221 40131 17279 40137
rect 17862 40128 17868 40140
rect 17920 40128 17926 40180
rect 25133 40171 25191 40177
rect 18248 40140 22968 40168
rect 10134 40060 10140 40112
rect 10192 40100 10198 40112
rect 10962 40100 10968 40112
rect 10192 40072 10968 40100
rect 10192 40060 10198 40072
rect 8662 39992 8668 40044
rect 8720 40032 8726 40044
rect 9582 40032 9588 40044
rect 8720 40004 9352 40032
rect 8720 39992 8726 40004
rect 9122 39924 9128 39976
rect 9180 39924 9186 39976
rect 9214 39924 9220 39976
rect 9272 39924 9278 39976
rect 9324 39973 9352 40004
rect 9416 40004 9588 40032
rect 9309 39967 9367 39973
rect 9309 39933 9321 39967
rect 9355 39933 9367 39967
rect 9309 39927 9367 39933
rect 8573 39899 8631 39905
rect 8573 39865 8585 39899
rect 8619 39865 8631 39899
rect 8573 39859 8631 39865
rect 8757 39899 8815 39905
rect 8757 39865 8769 39899
rect 8803 39896 8815 39899
rect 9416 39896 9444 40004
rect 9582 39992 9588 40004
rect 9640 39992 9646 40044
rect 10244 40041 10272 40072
rect 10962 40060 10968 40072
rect 11020 40100 11026 40112
rect 13262 40100 13268 40112
rect 11020 40072 11836 40100
rect 11020 40060 11026 40072
rect 10229 40035 10287 40041
rect 10229 40001 10241 40035
rect 10275 40001 10287 40035
rect 11330 40032 11336 40044
rect 10229 39995 10287 40001
rect 10520 40004 11336 40032
rect 9493 39967 9551 39973
rect 9493 39933 9505 39967
rect 9539 39933 9551 39967
rect 9493 39927 9551 39933
rect 8803 39868 9444 39896
rect 9508 39896 9536 39927
rect 9950 39924 9956 39976
rect 10008 39964 10014 39976
rect 10045 39967 10103 39973
rect 10045 39964 10057 39967
rect 10008 39936 10057 39964
rect 10008 39924 10014 39936
rect 10045 39933 10057 39936
rect 10091 39964 10103 39967
rect 10520 39964 10548 40004
rect 11330 39992 11336 40004
rect 11388 40032 11394 40044
rect 11808 40041 11836 40072
rect 13188 40072 13268 40100
rect 11701 40035 11759 40041
rect 11701 40032 11713 40035
rect 11388 40004 11713 40032
rect 11388 39992 11394 40004
rect 11701 40001 11713 40004
rect 11747 40001 11759 40035
rect 11701 39995 11759 40001
rect 11793 40035 11851 40041
rect 11793 40001 11805 40035
rect 11839 40001 11851 40035
rect 11793 39995 11851 40001
rect 10091 39936 10548 39964
rect 10091 39933 10103 39936
rect 10045 39927 10103 39933
rect 10594 39924 10600 39976
rect 10652 39924 10658 39976
rect 10686 39924 10692 39976
rect 10744 39924 10750 39976
rect 10870 39924 10876 39976
rect 10928 39924 10934 39976
rect 10965 39967 11023 39973
rect 10965 39933 10977 39967
rect 11011 39964 11023 39967
rect 11716 39964 11744 39995
rect 13078 39992 13084 40044
rect 13136 39992 13142 40044
rect 13188 40041 13216 40072
rect 13262 40060 13268 40072
rect 13320 40060 13326 40112
rect 16758 40100 16764 40112
rect 16408 40072 16764 40100
rect 13173 40035 13231 40041
rect 13173 40001 13185 40035
rect 13219 40001 13231 40035
rect 13173 39995 13231 40001
rect 15010 39992 15016 40044
rect 15068 40032 15074 40044
rect 15378 40032 15384 40044
rect 15068 40004 15384 40032
rect 15068 39992 15074 40004
rect 15378 39992 15384 40004
rect 15436 39992 15442 40044
rect 12253 39967 12311 39973
rect 12253 39964 12265 39967
rect 11011 39936 11284 39964
rect 11716 39936 12265 39964
rect 11011 39933 11023 39936
rect 10965 39927 11023 39933
rect 10226 39896 10232 39908
rect 9508 39868 10232 39896
rect 8803 39865 8815 39868
rect 8757 39859 8815 39865
rect 8386 39788 8392 39840
rect 8444 39788 8450 39840
rect 8588 39828 8616 39859
rect 10226 39856 10232 39868
rect 10284 39856 10290 39908
rect 10318 39856 10324 39908
rect 10376 39896 10382 39908
rect 10888 39896 10916 39924
rect 10376 39868 10916 39896
rect 10376 39856 10382 39868
rect 9582 39828 9588 39840
rect 8588 39800 9588 39828
rect 9582 39788 9588 39800
rect 9640 39828 9646 39840
rect 11256 39837 11284 39936
rect 12253 39933 12265 39936
rect 12299 39933 12311 39967
rect 12253 39927 12311 39933
rect 13538 39924 13544 39976
rect 13596 39924 13602 39976
rect 14090 39924 14096 39976
rect 14148 39964 14154 39976
rect 15562 39964 15568 39976
rect 14148 39936 15568 39964
rect 14148 39924 14154 39936
rect 15562 39924 15568 39936
rect 15620 39924 15626 39976
rect 15657 39967 15715 39973
rect 15657 39933 15669 39967
rect 15703 39933 15715 39967
rect 15657 39927 15715 39933
rect 11330 39856 11336 39908
rect 11388 39896 11394 39908
rect 12158 39896 12164 39908
rect 11388 39868 12164 39896
rect 11388 39856 11394 39868
rect 12158 39856 12164 39868
rect 12216 39856 12222 39908
rect 12437 39899 12495 39905
rect 12437 39865 12449 39899
rect 12483 39896 12495 39899
rect 12710 39896 12716 39908
rect 12483 39868 12716 39896
rect 12483 39865 12495 39868
rect 12437 39859 12495 39865
rect 12710 39856 12716 39868
rect 12768 39856 12774 39908
rect 13446 39856 13452 39908
rect 13504 39896 13510 39908
rect 13786 39899 13844 39905
rect 13786 39896 13798 39899
rect 13504 39868 13798 39896
rect 13504 39856 13510 39868
rect 13786 39865 13798 39868
rect 13832 39865 13844 39899
rect 13786 39859 13844 39865
rect 10137 39831 10195 39837
rect 10137 39828 10149 39831
rect 9640 39800 10149 39828
rect 9640 39788 9646 39800
rect 10137 39797 10149 39800
rect 10183 39797 10195 39831
rect 10137 39791 10195 39797
rect 11241 39831 11299 39837
rect 11241 39797 11253 39831
rect 11287 39797 11299 39831
rect 11241 39791 11299 39797
rect 11606 39788 11612 39840
rect 11664 39788 11670 39840
rect 11882 39788 11888 39840
rect 11940 39828 11946 39840
rect 12069 39831 12127 39837
rect 12069 39828 12081 39831
rect 11940 39800 12081 39828
rect 11940 39788 11946 39800
rect 12069 39797 12081 39800
rect 12115 39797 12127 39831
rect 12069 39791 12127 39797
rect 12526 39788 12532 39840
rect 12584 39828 12590 39840
rect 12621 39831 12679 39837
rect 12621 39828 12633 39831
rect 12584 39800 12633 39828
rect 12584 39788 12590 39800
rect 12621 39797 12633 39800
rect 12667 39797 12679 39831
rect 12621 39791 12679 39797
rect 12894 39788 12900 39840
rect 12952 39828 12958 39840
rect 12989 39831 13047 39837
rect 12989 39828 13001 39831
rect 12952 39800 13001 39828
rect 12952 39788 12958 39800
rect 12989 39797 13001 39800
rect 13035 39828 13047 39831
rect 13630 39828 13636 39840
rect 13035 39800 13636 39828
rect 13035 39797 13047 39800
rect 12989 39791 13047 39797
rect 13630 39788 13636 39800
rect 13688 39788 13694 39840
rect 14918 39788 14924 39840
rect 14976 39788 14982 39840
rect 15672 39828 15700 39927
rect 15838 39924 15844 39976
rect 15896 39924 15902 39976
rect 15930 39924 15936 39976
rect 15988 39924 15994 39976
rect 16408 39973 16436 40072
rect 16758 40060 16764 40072
rect 16816 40100 16822 40112
rect 17770 40100 17776 40112
rect 16816 40072 17776 40100
rect 16816 40060 16822 40072
rect 17770 40060 17776 40072
rect 17828 40100 17834 40112
rect 18138 40100 18144 40112
rect 17828 40072 18144 40100
rect 17828 40060 17834 40072
rect 18138 40060 18144 40072
rect 18196 40060 18202 40112
rect 16666 40032 16672 40044
rect 16500 40004 16672 40032
rect 16500 39973 16528 40004
rect 16666 39992 16672 40004
rect 16724 39992 16730 40044
rect 18248 40032 18276 40140
rect 17420 40004 18276 40032
rect 17420 39976 17448 40004
rect 18874 39992 18880 40044
rect 18932 40032 18938 40044
rect 20073 40035 20131 40041
rect 20073 40032 20085 40035
rect 18932 40004 20085 40032
rect 18932 39992 18938 40004
rect 20073 40001 20085 40004
rect 20119 40001 20131 40035
rect 21560 40032 21588 40140
rect 22186 40100 22192 40112
rect 22066 40072 22192 40100
rect 21913 40035 21971 40041
rect 21560 40004 21680 40032
rect 20073 39995 20131 40001
rect 16393 39967 16451 39973
rect 16393 39933 16405 39967
rect 16439 39933 16451 39967
rect 16393 39927 16451 39933
rect 16485 39967 16543 39973
rect 16485 39933 16497 39967
rect 16531 39933 16543 39967
rect 16485 39927 16543 39933
rect 16574 39924 16580 39976
rect 16632 39924 16638 39976
rect 16761 39967 16819 39973
rect 16761 39933 16773 39967
rect 16807 39964 16819 39967
rect 16942 39964 16948 39976
rect 16807 39936 16948 39964
rect 16807 39933 16819 39936
rect 16761 39927 16819 39933
rect 16942 39924 16948 39936
rect 17000 39924 17006 39976
rect 17126 39924 17132 39976
rect 17184 39924 17190 39976
rect 17313 39967 17371 39973
rect 17313 39933 17325 39967
rect 17359 39964 17371 39967
rect 17402 39964 17408 39976
rect 17359 39936 17408 39964
rect 17359 39933 17371 39936
rect 17313 39927 17371 39933
rect 17402 39924 17408 39936
rect 17460 39924 17466 39976
rect 18325 39967 18383 39973
rect 18325 39933 18337 39967
rect 18371 39933 18383 39967
rect 18325 39927 18383 39933
rect 18417 39967 18475 39973
rect 18417 39933 18429 39967
rect 18463 39964 18475 39967
rect 18693 39967 18751 39973
rect 18693 39964 18705 39967
rect 18463 39936 18705 39964
rect 18463 39933 18475 39936
rect 18417 39927 18475 39933
rect 18693 39933 18705 39936
rect 18739 39933 18751 39967
rect 18693 39927 18751 39933
rect 18340 39896 18368 39927
rect 18966 39924 18972 39976
rect 19024 39924 19030 39976
rect 19794 39924 19800 39976
rect 19852 39964 19858 39976
rect 20441 39967 20499 39973
rect 20441 39964 20453 39967
rect 19852 39936 20453 39964
rect 19852 39924 19858 39936
rect 20441 39933 20453 39936
rect 20487 39933 20499 39967
rect 20441 39927 20499 39933
rect 20625 39967 20683 39973
rect 20625 39933 20637 39967
rect 20671 39933 20683 39967
rect 20625 39927 20683 39933
rect 16500 39868 18368 39896
rect 16500 39840 16528 39868
rect 20346 39856 20352 39908
rect 20404 39896 20410 39908
rect 20640 39896 20668 39927
rect 21082 39924 21088 39976
rect 21140 39964 21146 39976
rect 21269 39967 21327 39973
rect 21269 39964 21281 39967
rect 21140 39936 21281 39964
rect 21140 39924 21146 39936
rect 21269 39933 21281 39936
rect 21315 39933 21327 39967
rect 21269 39927 21327 39933
rect 21450 39924 21456 39976
rect 21508 39924 21514 39976
rect 21652 39973 21680 40004
rect 21913 40001 21925 40035
rect 21959 40032 21971 40035
rect 22066 40032 22094 40072
rect 22186 40060 22192 40072
rect 22244 40060 22250 40112
rect 22940 40109 22968 40140
rect 25133 40137 25145 40171
rect 25179 40168 25191 40171
rect 26878 40168 26884 40180
rect 25179 40140 26884 40168
rect 25179 40137 25191 40140
rect 25133 40131 25191 40137
rect 26878 40128 26884 40140
rect 26936 40128 26942 40180
rect 27430 40128 27436 40180
rect 27488 40128 27494 40180
rect 28534 40128 28540 40180
rect 28592 40168 28598 40180
rect 28629 40171 28687 40177
rect 28629 40168 28641 40171
rect 28592 40140 28641 40168
rect 28592 40128 28598 40140
rect 28629 40137 28641 40140
rect 28675 40137 28687 40171
rect 28629 40131 28687 40137
rect 22925 40103 22983 40109
rect 22925 40069 22937 40103
rect 22971 40100 22983 40103
rect 23014 40100 23020 40112
rect 22971 40072 23020 40100
rect 22971 40069 22983 40072
rect 22925 40063 22983 40069
rect 23014 40060 23020 40072
rect 23072 40100 23078 40112
rect 23382 40100 23388 40112
rect 23072 40072 23388 40100
rect 23072 40060 23078 40072
rect 23382 40060 23388 40072
rect 23440 40060 23446 40112
rect 26050 40060 26056 40112
rect 26108 40100 26114 40112
rect 26145 40103 26203 40109
rect 26145 40100 26157 40103
rect 26108 40072 26157 40100
rect 26108 40060 26114 40072
rect 26145 40069 26157 40072
rect 26191 40100 26203 40103
rect 27448 40100 27476 40128
rect 28442 40100 28448 40112
rect 26191 40072 27476 40100
rect 28000 40072 28448 40100
rect 26191 40069 26203 40072
rect 26145 40063 26203 40069
rect 28000 40041 28028 40072
rect 28442 40060 28448 40072
rect 28500 40100 28506 40112
rect 28902 40100 28908 40112
rect 28500 40072 28908 40100
rect 28500 40060 28506 40072
rect 28902 40060 28908 40072
rect 28960 40060 28966 40112
rect 27985 40035 28043 40041
rect 21959 40004 22094 40032
rect 22388 40004 24348 40032
rect 21959 40001 21971 40004
rect 21913 39995 21971 40001
rect 22388 39976 22416 40004
rect 21545 39967 21603 39973
rect 21545 39933 21557 39967
rect 21591 39933 21603 39967
rect 21545 39927 21603 39933
rect 21637 39967 21695 39973
rect 21637 39933 21649 39967
rect 21683 39933 21695 39967
rect 21637 39927 21695 39933
rect 22189 39967 22247 39973
rect 22189 39933 22201 39967
rect 22235 39964 22247 39967
rect 22370 39964 22376 39976
rect 22235 39936 22376 39964
rect 22235 39933 22247 39936
rect 22189 39927 22247 39933
rect 20404 39868 20668 39896
rect 20404 39856 20410 39868
rect 16390 39828 16396 39840
rect 15672 39800 16396 39828
rect 16390 39788 16396 39800
rect 16448 39788 16454 39840
rect 16482 39788 16488 39840
rect 16540 39788 16546 39840
rect 16666 39788 16672 39840
rect 16724 39828 16730 39840
rect 17310 39828 17316 39840
rect 16724 39800 17316 39828
rect 16724 39788 16730 39800
rect 17310 39788 17316 39800
rect 17368 39788 17374 39840
rect 20530 39788 20536 39840
rect 20588 39788 20594 39840
rect 20622 39788 20628 39840
rect 20680 39828 20686 39840
rect 21560 39828 21588 39927
rect 22370 39924 22376 39936
rect 22428 39924 22434 39976
rect 23198 39924 23204 39976
rect 23256 39964 23262 39976
rect 23293 39967 23351 39973
rect 23293 39964 23305 39967
rect 23256 39936 23305 39964
rect 23256 39924 23262 39936
rect 23293 39933 23305 39936
rect 23339 39933 23351 39967
rect 23293 39927 23351 39933
rect 23382 39924 23388 39976
rect 23440 39964 23446 39976
rect 23477 39967 23535 39973
rect 23477 39964 23489 39967
rect 23440 39936 23489 39964
rect 23440 39924 23446 39936
rect 23477 39933 23489 39936
rect 23523 39933 23535 39967
rect 23477 39927 23535 39933
rect 23658 39924 23664 39976
rect 23716 39924 23722 39976
rect 24320 39973 24348 40004
rect 27985 40001 27997 40035
rect 28031 40001 28043 40035
rect 27985 39995 28043 40001
rect 28169 40035 28227 40041
rect 28169 40001 28181 40035
rect 28215 40032 28227 40035
rect 28350 40032 28356 40044
rect 28215 40004 28356 40032
rect 28215 40001 28227 40004
rect 28169 39995 28227 40001
rect 28350 39992 28356 40004
rect 28408 40032 28414 40044
rect 28718 40032 28724 40044
rect 28408 40004 28724 40032
rect 28408 39992 28414 40004
rect 28718 39992 28724 40004
rect 28776 39992 28782 40044
rect 30929 40035 30987 40041
rect 30929 40032 30941 40035
rect 30392 40004 30941 40032
rect 24305 39967 24363 39973
rect 24305 39933 24317 39967
rect 24351 39933 24363 39967
rect 24305 39927 24363 39933
rect 25590 39924 25596 39976
rect 25648 39964 25654 39976
rect 25961 39967 26019 39973
rect 25961 39964 25973 39967
rect 25648 39936 25973 39964
rect 25648 39924 25654 39936
rect 25961 39933 25973 39936
rect 26007 39933 26019 39967
rect 25961 39927 26019 39933
rect 26326 39924 26332 39976
rect 26384 39924 26390 39976
rect 26510 39924 26516 39976
rect 26568 39964 26574 39976
rect 27065 39967 27123 39973
rect 27065 39964 27077 39967
rect 26568 39936 27077 39964
rect 26568 39924 26574 39936
rect 27065 39933 27077 39936
rect 27111 39964 27123 39967
rect 28077 39967 28135 39973
rect 27111 39936 27936 39964
rect 27111 39933 27123 39936
rect 27065 39927 27123 39933
rect 22649 39899 22707 39905
rect 22649 39865 22661 39899
rect 22695 39896 22707 39899
rect 23566 39896 23572 39908
rect 22695 39868 23572 39896
rect 22695 39865 22707 39868
rect 22649 39859 22707 39865
rect 23566 39856 23572 39868
rect 23624 39856 23630 39908
rect 25038 39856 25044 39908
rect 25096 39905 25102 39908
rect 25096 39899 25159 39905
rect 25096 39865 25113 39899
rect 25147 39865 25159 39899
rect 25096 39859 25159 39865
rect 25096 39856 25102 39859
rect 25222 39856 25228 39908
rect 25280 39896 25286 39908
rect 25317 39899 25375 39905
rect 25317 39896 25329 39899
rect 25280 39868 25329 39896
rect 25280 39856 25286 39868
rect 25317 39865 25329 39868
rect 25363 39865 25375 39899
rect 25317 39859 25375 39865
rect 27433 39899 27491 39905
rect 27433 39865 27445 39899
rect 27479 39896 27491 39899
rect 27479 39868 27844 39896
rect 27479 39865 27491 39868
rect 27433 39859 27491 39865
rect 20680 39800 21588 39828
rect 20680 39788 20686 39800
rect 22094 39788 22100 39840
rect 22152 39788 22158 39840
rect 22465 39831 22523 39837
rect 22465 39797 22477 39831
rect 22511 39828 22523 39831
rect 22738 39828 22744 39840
rect 22511 39800 22744 39828
rect 22511 39797 22523 39800
rect 22465 39791 22523 39797
rect 22738 39788 22744 39800
rect 22796 39788 22802 39840
rect 22922 39788 22928 39840
rect 22980 39828 22986 39840
rect 23109 39831 23167 39837
rect 23109 39828 23121 39831
rect 22980 39800 23121 39828
rect 22980 39788 22986 39800
rect 23109 39797 23121 39800
rect 23155 39797 23167 39831
rect 23109 39791 23167 39797
rect 24210 39788 24216 39840
rect 24268 39828 24274 39840
rect 24397 39831 24455 39837
rect 24397 39828 24409 39831
rect 24268 39800 24409 39828
rect 24268 39788 24274 39800
rect 24397 39797 24409 39800
rect 24443 39797 24455 39831
rect 24397 39791 24455 39797
rect 24854 39788 24860 39840
rect 24912 39828 24918 39840
rect 24949 39831 25007 39837
rect 24949 39828 24961 39831
rect 24912 39800 24961 39828
rect 24912 39788 24918 39800
rect 24949 39797 24961 39800
rect 24995 39797 25007 39831
rect 24949 39791 25007 39797
rect 25406 39788 25412 39840
rect 25464 39788 25470 39840
rect 27617 39831 27675 39837
rect 27617 39797 27629 39831
rect 27663 39828 27675 39831
rect 27706 39828 27712 39840
rect 27663 39800 27712 39828
rect 27663 39797 27675 39800
rect 27617 39791 27675 39797
rect 27706 39788 27712 39800
rect 27764 39788 27770 39840
rect 27816 39837 27844 39868
rect 27801 39831 27859 39837
rect 27801 39797 27813 39831
rect 27847 39797 27859 39831
rect 27908 39828 27936 39936
rect 28077 39933 28089 39967
rect 28123 39933 28135 39967
rect 28077 39927 28135 39933
rect 28261 39967 28319 39973
rect 28261 39933 28273 39967
rect 28307 39964 28319 39967
rect 28534 39964 28540 39976
rect 28307 39936 28540 39964
rect 28307 39933 28319 39936
rect 28261 39927 28319 39933
rect 28092 39896 28120 39927
rect 28534 39924 28540 39936
rect 28592 39924 28598 39976
rect 29914 39924 29920 39976
rect 29972 39964 29978 39976
rect 30392 39973 30420 40004
rect 30929 40001 30941 40004
rect 30975 40001 30987 40035
rect 30929 39995 30987 40001
rect 30377 39967 30435 39973
rect 30377 39964 30389 39967
rect 29972 39936 30389 39964
rect 29972 39924 29978 39936
rect 30377 39933 30389 39936
rect 30423 39933 30435 39967
rect 30377 39927 30435 39933
rect 30558 39924 30564 39976
rect 30616 39964 30622 39976
rect 30745 39967 30803 39973
rect 30745 39964 30757 39967
rect 30616 39936 30757 39964
rect 30616 39924 30622 39936
rect 30745 39933 30757 39936
rect 30791 39933 30803 39967
rect 30745 39927 30803 39933
rect 31018 39924 31024 39976
rect 31076 39924 31082 39976
rect 28350 39896 28356 39908
rect 28092 39868 28356 39896
rect 28350 39856 28356 39868
rect 28408 39896 28414 39908
rect 28810 39896 28816 39908
rect 28408 39868 28816 39896
rect 28408 39856 28414 39868
rect 28810 39856 28816 39868
rect 28868 39856 28874 39908
rect 29270 39856 29276 39908
rect 29328 39896 29334 39908
rect 31036 39896 31064 39924
rect 29328 39868 31064 39896
rect 29328 39856 29334 39868
rect 28626 39837 28632 39840
rect 28445 39831 28503 39837
rect 28445 39828 28457 39831
rect 27908 39800 28457 39828
rect 27801 39791 27859 39797
rect 28445 39797 28457 39800
rect 28491 39797 28503 39831
rect 28445 39791 28503 39797
rect 28613 39831 28632 39837
rect 28613 39797 28625 39831
rect 28613 39791 28632 39797
rect 28626 39788 28632 39791
rect 28684 39788 28690 39840
rect 29822 39788 29828 39840
rect 29880 39788 29886 39840
rect 30374 39788 30380 39840
rect 30432 39828 30438 39840
rect 30561 39831 30619 39837
rect 30561 39828 30573 39831
rect 30432 39800 30573 39828
rect 30432 39788 30438 39800
rect 30561 39797 30573 39800
rect 30607 39797 30619 39831
rect 30561 39791 30619 39797
rect 31113 39831 31171 39837
rect 31113 39797 31125 39831
rect 31159 39828 31171 39831
rect 31159 39800 31708 39828
rect 31159 39797 31171 39800
rect 31113 39791 31171 39797
rect 552 39738 31648 39760
rect 552 39686 4322 39738
rect 4374 39686 4386 39738
rect 4438 39686 4450 39738
rect 4502 39686 4514 39738
rect 4566 39686 4578 39738
rect 4630 39686 12096 39738
rect 12148 39686 12160 39738
rect 12212 39686 12224 39738
rect 12276 39686 12288 39738
rect 12340 39686 12352 39738
rect 12404 39686 19870 39738
rect 19922 39686 19934 39738
rect 19986 39686 19998 39738
rect 20050 39686 20062 39738
rect 20114 39686 20126 39738
rect 20178 39686 27644 39738
rect 27696 39686 27708 39738
rect 27760 39686 27772 39738
rect 27824 39686 27836 39738
rect 27888 39686 27900 39738
rect 27952 39686 31648 39738
rect 552 39664 31648 39686
rect 9766 39584 9772 39636
rect 9824 39624 9830 39636
rect 10229 39627 10287 39633
rect 10229 39624 10241 39627
rect 9824 39596 10241 39624
rect 9824 39584 9830 39596
rect 10229 39593 10241 39596
rect 10275 39593 10287 39627
rect 10229 39587 10287 39593
rect 10686 39584 10692 39636
rect 10744 39624 10750 39636
rect 11241 39627 11299 39633
rect 11241 39624 11253 39627
rect 10744 39596 11253 39624
rect 10744 39584 10750 39596
rect 11241 39593 11253 39596
rect 11287 39593 11299 39627
rect 11606 39624 11612 39636
rect 11241 39587 11299 39593
rect 11532 39596 11612 39624
rect 10042 39556 10048 39568
rect 9876 39528 10048 39556
rect 8386 39448 8392 39500
rect 8444 39488 8450 39500
rect 9585 39491 9643 39497
rect 9585 39488 9597 39491
rect 8444 39460 9597 39488
rect 8444 39448 8450 39460
rect 9585 39457 9597 39460
rect 9631 39457 9643 39491
rect 9585 39451 9643 39457
rect 9766 39448 9772 39500
rect 9824 39448 9830 39500
rect 9876 39497 9904 39528
rect 10042 39516 10048 39528
rect 10100 39556 10106 39568
rect 10962 39556 10968 39568
rect 10100 39528 10968 39556
rect 10100 39516 10106 39528
rect 10962 39516 10968 39528
rect 11020 39516 11026 39568
rect 9861 39491 9919 39497
rect 9861 39457 9873 39491
rect 9907 39457 9919 39491
rect 9861 39451 9919 39457
rect 9950 39448 9956 39500
rect 10008 39448 10014 39500
rect 11532 39497 11560 39596
rect 11606 39584 11612 39596
rect 11664 39624 11670 39636
rect 11664 39596 12112 39624
rect 11664 39584 11670 39596
rect 11974 39556 11980 39568
rect 11624 39528 11980 39556
rect 11624 39497 11652 39528
rect 11974 39516 11980 39528
rect 12032 39516 12038 39568
rect 11517 39491 11575 39497
rect 11517 39457 11529 39491
rect 11563 39457 11575 39491
rect 11517 39451 11575 39457
rect 11609 39491 11667 39497
rect 11609 39457 11621 39491
rect 11655 39457 11667 39491
rect 11609 39451 11667 39457
rect 11698 39448 11704 39500
rect 11756 39448 11762 39500
rect 11882 39448 11888 39500
rect 11940 39448 11946 39500
rect 9214 39380 9220 39432
rect 9272 39420 9278 39432
rect 11330 39420 11336 39432
rect 9272 39392 11336 39420
rect 9272 39380 9278 39392
rect 11330 39380 11336 39392
rect 11388 39380 11394 39432
rect 9766 39312 9772 39364
rect 9824 39352 9830 39364
rect 11716 39352 11744 39448
rect 12084 39420 12112 39596
rect 12434 39584 12440 39636
rect 12492 39624 12498 39636
rect 12492 39596 12756 39624
rect 12492 39584 12498 39596
rect 12526 39556 12532 39568
rect 12360 39528 12532 39556
rect 12360 39497 12388 39528
rect 12526 39516 12532 39528
rect 12584 39516 12590 39568
rect 12345 39491 12403 39497
rect 12345 39457 12357 39491
rect 12391 39457 12403 39491
rect 12345 39451 12403 39457
rect 12437 39491 12495 39497
rect 12437 39457 12449 39491
rect 12483 39488 12495 39491
rect 12483 39460 12572 39488
rect 12483 39457 12495 39460
rect 12437 39451 12495 39457
rect 12544 39432 12572 39460
rect 12618 39448 12624 39500
rect 12676 39448 12682 39500
rect 12728 39497 12756 39596
rect 13446 39584 13452 39636
rect 13504 39584 13510 39636
rect 13538 39584 13544 39636
rect 13596 39624 13602 39636
rect 13725 39627 13783 39633
rect 13725 39624 13737 39627
rect 13596 39596 13737 39624
rect 13596 39584 13602 39596
rect 13725 39593 13737 39596
rect 13771 39593 13783 39627
rect 13725 39587 13783 39593
rect 15289 39627 15347 39633
rect 15289 39593 15301 39627
rect 15335 39624 15347 39627
rect 15470 39624 15476 39636
rect 15335 39596 15476 39624
rect 15335 39593 15347 39596
rect 15289 39587 15347 39593
rect 15470 39584 15476 39596
rect 15528 39584 15534 39636
rect 15657 39627 15715 39633
rect 15657 39593 15669 39627
rect 15703 39624 15715 39627
rect 17678 39624 17684 39636
rect 15703 39596 17684 39624
rect 15703 39593 15715 39596
rect 15657 39587 15715 39593
rect 17678 39584 17684 39596
rect 17736 39584 17742 39636
rect 18966 39584 18972 39636
rect 19024 39624 19030 39636
rect 19153 39627 19211 39633
rect 19153 39624 19165 39627
rect 19024 39596 19165 39624
rect 19024 39584 19030 39596
rect 19153 39593 19165 39596
rect 19199 39593 19211 39627
rect 22649 39627 22707 39633
rect 19153 39587 19211 39593
rect 20824 39596 22600 39624
rect 16482 39556 16488 39568
rect 13832 39528 16488 39556
rect 12713 39491 12771 39497
rect 12713 39457 12725 39491
rect 12759 39457 12771 39491
rect 12713 39451 12771 39457
rect 12805 39491 12863 39497
rect 12805 39457 12817 39491
rect 12851 39488 12863 39491
rect 12851 39460 12940 39488
rect 12851 39457 12863 39460
rect 12805 39451 12863 39457
rect 12084 39392 12434 39420
rect 9824 39324 11744 39352
rect 9824 39312 9830 39324
rect 12406 39296 12434 39392
rect 12526 39380 12532 39432
rect 12584 39380 12590 39432
rect 12618 39312 12624 39364
rect 12676 39352 12682 39364
rect 12728 39352 12756 39451
rect 12676 39324 12756 39352
rect 12676 39312 12682 39324
rect 9674 39244 9680 39296
rect 9732 39284 9738 39296
rect 10410 39284 10416 39296
rect 9732 39256 10416 39284
rect 9732 39244 9738 39256
rect 10410 39244 10416 39256
rect 10468 39244 10474 39296
rect 11882 39244 11888 39296
rect 11940 39284 11946 39296
rect 12161 39287 12219 39293
rect 12161 39284 12173 39287
rect 11940 39256 12173 39284
rect 11940 39244 11946 39256
rect 12161 39253 12173 39256
rect 12207 39253 12219 39287
rect 12406 39256 12440 39296
rect 12161 39247 12219 39253
rect 12434 39244 12440 39256
rect 12492 39244 12498 39296
rect 12912 39284 12940 39460
rect 12986 39448 12992 39500
rect 13044 39448 13050 39500
rect 13832 39497 13860 39528
rect 16482 39516 16488 39528
rect 16540 39516 16546 39568
rect 17126 39516 17132 39568
rect 17184 39556 17190 39568
rect 20824 39556 20852 39596
rect 22094 39556 22100 39568
rect 17184 39528 20852 39556
rect 17184 39516 17190 39528
rect 13081 39491 13139 39497
rect 13081 39457 13093 39491
rect 13127 39457 13139 39491
rect 13081 39451 13139 39457
rect 13173 39491 13231 39497
rect 13173 39457 13185 39491
rect 13219 39457 13231 39491
rect 13173 39451 13231 39457
rect 13817 39491 13875 39497
rect 13817 39457 13829 39491
rect 13863 39457 13875 39491
rect 13817 39451 13875 39457
rect 15473 39491 15531 39497
rect 15473 39457 15485 39491
rect 15519 39457 15531 39491
rect 15473 39451 15531 39457
rect 13096 39352 13124 39451
rect 13188 39420 13216 39451
rect 14001 39423 14059 39429
rect 14001 39420 14013 39423
rect 13188 39392 14013 39420
rect 14001 39389 14013 39392
rect 14047 39389 14059 39423
rect 14001 39383 14059 39389
rect 14553 39423 14611 39429
rect 14553 39389 14565 39423
rect 14599 39420 14611 39423
rect 14918 39420 14924 39432
rect 14599 39392 14924 39420
rect 14599 39389 14611 39392
rect 14553 39383 14611 39389
rect 13630 39352 13636 39364
rect 13096 39324 13636 39352
rect 13630 39312 13636 39324
rect 13688 39312 13694 39364
rect 13722 39312 13728 39364
rect 13780 39352 13786 39364
rect 14568 39352 14596 39383
rect 14918 39380 14924 39392
rect 14976 39380 14982 39432
rect 15488 39420 15516 39451
rect 15562 39448 15568 39500
rect 15620 39488 15626 39500
rect 15749 39491 15807 39497
rect 15749 39488 15761 39491
rect 15620 39460 15761 39488
rect 15620 39448 15626 39460
rect 15749 39457 15761 39460
rect 15795 39457 15807 39491
rect 15749 39451 15807 39457
rect 18506 39448 18512 39500
rect 18564 39448 18570 39500
rect 18690 39448 18696 39500
rect 18748 39448 18754 39500
rect 18785 39491 18843 39497
rect 18785 39457 18797 39491
rect 18831 39457 18843 39491
rect 18785 39451 18843 39457
rect 15838 39420 15844 39432
rect 15488 39392 15844 39420
rect 15838 39380 15844 39392
rect 15896 39380 15902 39432
rect 18800 39420 18828 39451
rect 18874 39448 18880 39500
rect 18932 39448 18938 39500
rect 19242 39448 19248 39500
rect 19300 39448 19306 39500
rect 19429 39491 19487 39497
rect 19429 39457 19441 39491
rect 19475 39488 19487 39491
rect 19610 39488 19616 39500
rect 19475 39460 19616 39488
rect 19475 39457 19487 39460
rect 19429 39451 19487 39457
rect 19610 39448 19616 39460
rect 19668 39448 19674 39500
rect 19812 39497 19840 39528
rect 19797 39491 19855 39497
rect 19797 39457 19809 39491
rect 19843 39457 19855 39491
rect 19797 39451 19855 39457
rect 20162 39448 20168 39500
rect 20220 39448 20226 39500
rect 20346 39448 20352 39500
rect 20404 39448 20410 39500
rect 20438 39448 20444 39500
rect 20496 39448 20502 39500
rect 20824 39497 20852 39528
rect 21284 39528 22100 39556
rect 21284 39497 21312 39528
rect 22094 39516 22100 39528
rect 22152 39516 22158 39568
rect 22572 39556 22600 39596
rect 22649 39593 22661 39627
rect 22695 39624 22707 39627
rect 23566 39624 23572 39636
rect 22695 39596 23572 39624
rect 22695 39593 22707 39596
rect 22649 39587 22707 39593
rect 23566 39584 23572 39596
rect 23624 39584 23630 39636
rect 25590 39584 25596 39636
rect 25648 39584 25654 39636
rect 26053 39627 26111 39633
rect 26053 39593 26065 39627
rect 26099 39624 26111 39627
rect 26421 39627 26479 39633
rect 26421 39624 26433 39627
rect 26099 39596 26433 39624
rect 26099 39593 26111 39596
rect 26053 39587 26111 39593
rect 26421 39593 26433 39596
rect 26467 39593 26479 39627
rect 26421 39587 26479 39593
rect 23198 39556 23204 39568
rect 22572 39528 23204 39556
rect 23198 39516 23204 39528
rect 23256 39516 23262 39568
rect 26326 39516 26332 39568
rect 26384 39556 26390 39568
rect 26786 39556 26792 39568
rect 26384 39528 26792 39556
rect 26384 39516 26390 39528
rect 26786 39516 26792 39528
rect 26844 39516 26850 39568
rect 29454 39556 29460 39568
rect 29288 39528 29460 39556
rect 20625 39491 20683 39497
rect 20625 39457 20637 39491
rect 20671 39457 20683 39491
rect 20625 39451 20683 39457
rect 20717 39491 20775 39497
rect 20717 39457 20729 39491
rect 20763 39457 20775 39491
rect 20717 39451 20775 39457
rect 20809 39491 20867 39497
rect 20809 39457 20821 39491
rect 20855 39457 20867 39491
rect 20809 39451 20867 39457
rect 21269 39491 21327 39497
rect 21269 39457 21281 39491
rect 21315 39457 21327 39491
rect 21525 39491 21583 39497
rect 21525 39488 21537 39491
rect 21269 39451 21327 39457
rect 21376 39460 21537 39488
rect 19337 39423 19395 39429
rect 19337 39420 19349 39423
rect 18800 39392 19349 39420
rect 19337 39389 19349 39392
rect 19383 39389 19395 39423
rect 19337 39383 19395 39389
rect 20257 39423 20315 39429
rect 20257 39389 20269 39423
rect 20303 39420 20315 39423
rect 20640 39420 20668 39451
rect 20303 39392 20668 39420
rect 20303 39389 20315 39392
rect 20257 39383 20315 39389
rect 13780 39324 14596 39352
rect 13780 39312 13786 39324
rect 17770 39312 17776 39364
rect 17828 39352 17834 39364
rect 18874 39352 18880 39364
rect 17828 39324 18880 39352
rect 17828 39312 17834 39324
rect 18874 39312 18880 39324
rect 18932 39312 18938 39364
rect 20162 39312 20168 39364
rect 20220 39352 20226 39364
rect 20622 39352 20628 39364
rect 20220 39324 20628 39352
rect 20220 39312 20226 39324
rect 20622 39312 20628 39324
rect 20680 39352 20686 39364
rect 20732 39352 20760 39451
rect 21085 39423 21143 39429
rect 21085 39389 21097 39423
rect 21131 39420 21143 39423
rect 21376 39420 21404 39460
rect 21525 39457 21537 39460
rect 21571 39457 21583 39491
rect 21525 39451 21583 39457
rect 22738 39448 22744 39500
rect 22796 39448 22802 39500
rect 23008 39491 23066 39497
rect 23008 39457 23020 39491
rect 23054 39488 23066 39491
rect 23566 39488 23572 39500
rect 23054 39460 23572 39488
rect 23054 39457 23066 39460
rect 23008 39451 23066 39457
rect 23566 39448 23572 39460
rect 23624 39448 23630 39500
rect 24210 39448 24216 39500
rect 24268 39448 24274 39500
rect 24486 39497 24492 39500
rect 24480 39451 24492 39497
rect 24486 39448 24492 39451
rect 24544 39448 24550 39500
rect 24854 39448 24860 39500
rect 24912 39488 24918 39500
rect 25685 39491 25743 39497
rect 25685 39488 25697 39491
rect 24912 39460 25697 39488
rect 24912 39448 24918 39460
rect 25685 39457 25697 39460
rect 25731 39457 25743 39491
rect 25685 39451 25743 39457
rect 21131 39392 21404 39420
rect 21131 39389 21143 39392
rect 21085 39383 21143 39389
rect 26510 39380 26516 39432
rect 26568 39420 26574 39432
rect 26804 39429 26832 39516
rect 27338 39448 27344 39500
rect 27396 39448 27402 39500
rect 28350 39448 28356 39500
rect 28408 39497 28414 39500
rect 29288 39497 29316 39528
rect 29454 39516 29460 39528
rect 29512 39516 29518 39568
rect 28408 39491 28457 39497
rect 28408 39457 28411 39491
rect 28445 39457 28457 39491
rect 28408 39451 28457 39457
rect 29273 39491 29331 39497
rect 29273 39457 29285 39491
rect 29319 39457 29331 39491
rect 29273 39451 29331 39457
rect 28408 39448 28414 39451
rect 29822 39448 29828 39500
rect 29880 39448 29886 39500
rect 30190 39448 30196 39500
rect 30248 39488 30254 39500
rect 31030 39491 31088 39497
rect 31030 39488 31042 39491
rect 30248 39460 31042 39488
rect 30248 39448 30254 39460
rect 31030 39457 31042 39460
rect 31076 39457 31088 39491
rect 31030 39451 31088 39457
rect 31297 39491 31355 39497
rect 31297 39457 31309 39491
rect 31343 39488 31355 39491
rect 31680 39488 31708 39800
rect 31343 39460 31708 39488
rect 31343 39457 31355 39460
rect 31297 39451 31355 39457
rect 26605 39423 26663 39429
rect 26605 39420 26617 39423
rect 26568 39392 26617 39420
rect 26568 39380 26574 39392
rect 26605 39389 26617 39392
rect 26651 39389 26663 39423
rect 26605 39383 26663 39389
rect 26697 39423 26755 39429
rect 26697 39389 26709 39423
rect 26743 39389 26755 39423
rect 26697 39383 26755 39389
rect 26789 39423 26847 39429
rect 26789 39389 26801 39423
rect 26835 39389 26847 39423
rect 26789 39383 26847 39389
rect 20680 39324 20760 39352
rect 20680 39312 20686 39324
rect 25222 39312 25228 39364
rect 25280 39352 25286 39364
rect 26712 39352 26740 39383
rect 26878 39380 26884 39432
rect 26936 39380 26942 39432
rect 28074 39380 28080 39432
rect 28132 39420 28138 39432
rect 28261 39423 28319 39429
rect 28261 39420 28273 39423
rect 28132 39392 28273 39420
rect 28132 39380 28138 39392
rect 28261 39389 28273 39392
rect 28307 39389 28319 39423
rect 28261 39383 28319 39389
rect 28534 39380 28540 39432
rect 28592 39380 28598 39432
rect 28718 39380 28724 39432
rect 28776 39420 28782 39432
rect 29457 39423 29515 39429
rect 29457 39420 29469 39423
rect 28776 39392 29469 39420
rect 28776 39380 28782 39392
rect 29457 39389 29469 39392
rect 29503 39389 29515 39423
rect 29457 39383 29515 39389
rect 29546 39380 29552 39432
rect 29604 39380 29610 39432
rect 28813 39355 28871 39361
rect 28813 39352 28825 39355
rect 25280 39324 26740 39352
rect 28736 39324 28825 39352
rect 25280 39312 25286 39324
rect 28736 39296 28764 39324
rect 28813 39321 28825 39324
rect 28859 39321 28871 39355
rect 28813 39315 28871 39321
rect 29178 39312 29184 39364
rect 29236 39352 29242 39364
rect 29914 39352 29920 39364
rect 29236 39324 29920 39352
rect 29236 39312 29242 39324
rect 29914 39312 29920 39324
rect 29972 39312 29978 39364
rect 13354 39284 13360 39296
rect 12912 39256 13360 39284
rect 13354 39244 13360 39256
rect 13412 39284 13418 39296
rect 15378 39284 15384 39296
rect 13412 39256 15384 39284
rect 13412 39244 13418 39256
rect 15378 39244 15384 39256
rect 15436 39244 15442 39296
rect 18414 39244 18420 39296
rect 18472 39284 18478 39296
rect 19242 39284 19248 39296
rect 18472 39256 19248 39284
rect 18472 39244 18478 39256
rect 19242 39244 19248 39256
rect 19300 39244 19306 39296
rect 19886 39244 19892 39296
rect 19944 39244 19950 39296
rect 20438 39244 20444 39296
rect 20496 39284 20502 39296
rect 21082 39284 21088 39296
rect 20496 39256 21088 39284
rect 20496 39244 20502 39256
rect 21082 39244 21088 39256
rect 21140 39244 21146 39296
rect 23842 39244 23848 39296
rect 23900 39284 23906 39296
rect 24121 39287 24179 39293
rect 24121 39284 24133 39287
rect 23900 39256 24133 39284
rect 23900 39244 23906 39256
rect 24121 39253 24133 39256
rect 24167 39253 24179 39287
rect 24121 39247 24179 39253
rect 25130 39244 25136 39296
rect 25188 39284 25194 39296
rect 26050 39284 26056 39296
rect 25188 39256 26056 39284
rect 25188 39244 25194 39256
rect 26050 39244 26056 39256
rect 26108 39244 26114 39296
rect 26237 39287 26295 39293
rect 26237 39253 26249 39287
rect 26283 39284 26295 39287
rect 26786 39284 26792 39296
rect 26283 39256 26792 39284
rect 26283 39253 26295 39256
rect 26237 39247 26295 39253
rect 26786 39244 26792 39256
rect 26844 39244 26850 39296
rect 26878 39244 26884 39296
rect 26936 39284 26942 39296
rect 27249 39287 27307 39293
rect 27249 39284 27261 39287
rect 26936 39256 27261 39284
rect 26936 39244 26942 39256
rect 27249 39253 27261 39256
rect 27295 39253 27307 39287
rect 27249 39247 27307 39253
rect 27430 39244 27436 39296
rect 27488 39284 27494 39296
rect 27617 39287 27675 39293
rect 27617 39284 27629 39287
rect 27488 39256 27629 39284
rect 27488 39244 27494 39256
rect 27617 39253 27629 39256
rect 27663 39253 27675 39287
rect 27617 39247 27675 39253
rect 27706 39244 27712 39296
rect 27764 39284 27770 39296
rect 28718 39284 28724 39296
rect 27764 39256 28724 39284
rect 27764 39244 27770 39256
rect 28718 39244 28724 39256
rect 28776 39244 28782 39296
rect 29638 39244 29644 39296
rect 29696 39244 29702 39296
rect 29733 39287 29791 39293
rect 29733 39253 29745 39287
rect 29779 39284 29791 39287
rect 30558 39284 30564 39296
rect 29779 39256 30564 39284
rect 29779 39253 29791 39256
rect 29733 39247 29791 39253
rect 30558 39244 30564 39256
rect 30616 39244 30622 39296
rect 552 39194 31648 39216
rect 552 39142 3662 39194
rect 3714 39142 3726 39194
rect 3778 39142 3790 39194
rect 3842 39142 3854 39194
rect 3906 39142 3918 39194
rect 3970 39142 11436 39194
rect 11488 39142 11500 39194
rect 11552 39142 11564 39194
rect 11616 39142 11628 39194
rect 11680 39142 11692 39194
rect 11744 39142 19210 39194
rect 19262 39142 19274 39194
rect 19326 39142 19338 39194
rect 19390 39142 19402 39194
rect 19454 39142 19466 39194
rect 19518 39142 26984 39194
rect 27036 39142 27048 39194
rect 27100 39142 27112 39194
rect 27164 39142 27176 39194
rect 27228 39142 27240 39194
rect 27292 39142 31648 39194
rect 552 39120 31648 39142
rect 10594 39080 10600 39092
rect 9140 39052 10600 39080
rect 9140 38944 9168 39052
rect 10594 39040 10600 39052
rect 10652 39040 10658 39092
rect 10870 39040 10876 39092
rect 10928 39080 10934 39092
rect 12526 39080 12532 39092
rect 10928 39052 12532 39080
rect 10928 39040 10934 39052
rect 12526 39040 12532 39052
rect 12584 39080 12590 39092
rect 12802 39080 12808 39092
rect 12584 39052 12808 39080
rect 12584 39040 12590 39052
rect 12802 39040 12808 39052
rect 12860 39080 12866 39092
rect 16942 39080 16948 39092
rect 12860 39052 16948 39080
rect 12860 39040 12866 39052
rect 16942 39040 16948 39052
rect 17000 39040 17006 39092
rect 18506 39040 18512 39092
rect 18564 39080 18570 39092
rect 19426 39080 19432 39092
rect 18564 39052 19432 39080
rect 18564 39040 18570 39052
rect 19426 39040 19432 39052
rect 19484 39080 19490 39092
rect 20254 39080 20260 39092
rect 19484 39052 20260 39080
rect 19484 39040 19490 39052
rect 20254 39040 20260 39052
rect 20312 39040 20318 39092
rect 24486 39040 24492 39092
rect 24544 39080 24550 39092
rect 24673 39083 24731 39089
rect 24673 39080 24685 39083
rect 24544 39052 24685 39080
rect 24544 39040 24550 39052
rect 24673 39049 24685 39052
rect 24719 39049 24731 39083
rect 24673 39043 24731 39049
rect 24854 39040 24860 39092
rect 24912 39080 24918 39092
rect 25041 39083 25099 39089
rect 25041 39080 25053 39083
rect 24912 39052 25053 39080
rect 24912 39040 24918 39052
rect 25041 39049 25053 39052
rect 25087 39049 25099 39083
rect 26326 39080 26332 39092
rect 25041 39043 25099 39049
rect 25516 39052 26332 39080
rect 10888 39012 10916 39040
rect 9048 38916 9168 38944
rect 9324 38984 10916 39012
rect 8294 38836 8300 38888
rect 8352 38876 8358 38888
rect 9048 38885 9076 38916
rect 8573 38879 8631 38885
rect 8573 38876 8585 38879
rect 8352 38848 8585 38876
rect 8352 38836 8358 38848
rect 8573 38845 8585 38848
rect 8619 38845 8631 38879
rect 8573 38839 8631 38845
rect 9033 38879 9091 38885
rect 9033 38845 9045 38879
rect 9079 38845 9091 38879
rect 9033 38839 9091 38845
rect 9122 38836 9128 38888
rect 9180 38836 9186 38888
rect 9324 38885 9352 38984
rect 15562 38972 15568 39024
rect 15620 39012 15626 39024
rect 16393 39015 16451 39021
rect 16393 39012 16405 39015
rect 15620 38984 16405 39012
rect 15620 38972 15626 38984
rect 16393 38981 16405 38984
rect 16439 38981 16451 39015
rect 16393 38975 16451 38981
rect 17405 39015 17463 39021
rect 17405 38981 17417 39015
rect 17451 38981 17463 39015
rect 17405 38975 17463 38981
rect 9582 38904 9588 38956
rect 9640 38944 9646 38956
rect 10229 38947 10287 38953
rect 10229 38944 10241 38947
rect 9640 38916 10241 38944
rect 9640 38904 9646 38916
rect 10229 38913 10241 38916
rect 10275 38913 10287 38947
rect 10229 38907 10287 38913
rect 10962 38904 10968 38956
rect 11020 38944 11026 38956
rect 13630 38944 13636 38956
rect 11020 38916 13636 38944
rect 11020 38904 11026 38916
rect 13630 38904 13636 38916
rect 13688 38904 13694 38956
rect 16942 38904 16948 38956
rect 17000 38944 17006 38956
rect 17420 38944 17448 38975
rect 19518 38972 19524 39024
rect 19576 39012 19582 39024
rect 19886 39012 19892 39024
rect 19576 38984 19892 39012
rect 19576 38972 19582 38984
rect 19886 38972 19892 38984
rect 19944 38972 19950 39024
rect 23474 39012 23480 39024
rect 19996 38984 23480 39012
rect 19996 38944 20024 38984
rect 23474 38972 23480 38984
rect 23532 38972 23538 39024
rect 25406 38972 25412 39024
rect 25464 38972 25470 39024
rect 22922 38944 22928 38956
rect 17000 38916 17448 38944
rect 19720 38916 20024 38944
rect 20088 38916 22928 38944
rect 17000 38904 17006 38916
rect 9309 38879 9367 38885
rect 9309 38845 9321 38879
rect 9355 38845 9367 38879
rect 9309 38839 9367 38845
rect 9401 38879 9459 38885
rect 9401 38845 9413 38879
rect 9447 38876 9459 38879
rect 9674 38876 9680 38888
rect 9447 38848 9680 38876
rect 9447 38845 9459 38848
rect 9401 38839 9459 38845
rect 9674 38836 9680 38848
rect 9732 38836 9738 38888
rect 12345 38879 12403 38885
rect 12345 38845 12357 38879
rect 12391 38876 12403 38879
rect 12434 38876 12440 38888
rect 12391 38848 12440 38876
rect 12391 38845 12403 38848
rect 12345 38839 12403 38845
rect 12434 38836 12440 38848
rect 12492 38836 12498 38888
rect 15565 38879 15623 38885
rect 15565 38845 15577 38879
rect 15611 38876 15623 38879
rect 15654 38876 15660 38888
rect 15611 38848 15660 38876
rect 15611 38845 15623 38848
rect 15565 38839 15623 38845
rect 15654 38836 15660 38848
rect 15712 38836 15718 38888
rect 15749 38879 15807 38885
rect 15749 38845 15761 38879
rect 15795 38876 15807 38879
rect 16206 38876 16212 38888
rect 15795 38848 16212 38876
rect 15795 38845 15807 38848
rect 15749 38839 15807 38845
rect 16206 38836 16212 38848
rect 16264 38836 16270 38888
rect 16301 38879 16359 38885
rect 16301 38845 16313 38879
rect 16347 38876 16359 38879
rect 16482 38876 16488 38888
rect 16347 38848 16488 38876
rect 16347 38845 16359 38848
rect 16301 38839 16359 38845
rect 16482 38836 16488 38848
rect 16540 38876 16546 38888
rect 16540 38848 16988 38876
rect 16540 38836 16546 38848
rect 16960 38820 16988 38848
rect 17218 38836 17224 38888
rect 17276 38836 17282 38888
rect 17310 38836 17316 38888
rect 17368 38876 17374 38888
rect 19720 38876 19748 38916
rect 17368 38848 19748 38876
rect 17368 38836 17374 38848
rect 19794 38836 19800 38888
rect 19852 38876 19858 38888
rect 19981 38879 20039 38885
rect 19981 38876 19993 38879
rect 19852 38848 19993 38876
rect 19852 38836 19858 38848
rect 19981 38845 19993 38848
rect 20027 38845 20039 38879
rect 19981 38839 20039 38845
rect 9585 38811 9643 38817
rect 9585 38777 9597 38811
rect 9631 38808 9643 38811
rect 10042 38808 10048 38820
rect 9631 38780 10048 38808
rect 9631 38777 9643 38780
rect 9585 38771 9643 38777
rect 10042 38768 10048 38780
rect 10100 38768 10106 38820
rect 12161 38811 12219 38817
rect 12161 38777 12173 38811
rect 12207 38808 12219 38811
rect 12710 38808 12716 38820
rect 12207 38780 12716 38808
rect 12207 38777 12219 38780
rect 12161 38771 12219 38777
rect 12710 38768 12716 38780
rect 12768 38808 12774 38820
rect 12894 38808 12900 38820
rect 12768 38780 12900 38808
rect 12768 38768 12774 38780
rect 12894 38768 12900 38780
rect 12952 38768 12958 38820
rect 16942 38768 16948 38820
rect 17000 38768 17006 38820
rect 18414 38768 18420 38820
rect 18472 38808 18478 38820
rect 20088 38808 20116 38916
rect 22922 38904 22928 38916
rect 22980 38904 22986 38956
rect 25133 38947 25191 38953
rect 25133 38913 25145 38947
rect 25179 38944 25191 38947
rect 25424 38944 25452 38972
rect 25179 38916 25452 38944
rect 25179 38913 25191 38916
rect 25133 38907 25191 38913
rect 24857 38879 24915 38885
rect 24857 38845 24869 38879
rect 24903 38876 24915 38879
rect 25038 38876 25044 38888
rect 24903 38848 25044 38876
rect 24903 38845 24915 38848
rect 24857 38839 24915 38845
rect 25038 38836 25044 38848
rect 25096 38836 25102 38888
rect 25222 38836 25228 38888
rect 25280 38836 25286 38888
rect 25409 38879 25467 38885
rect 25409 38845 25421 38879
rect 25455 38876 25467 38879
rect 25516 38876 25544 39052
rect 26326 39040 26332 39052
rect 26384 39040 26390 39092
rect 26602 39040 26608 39092
rect 26660 39080 26666 39092
rect 27157 39083 27215 39089
rect 27157 39080 27169 39083
rect 26660 39052 27169 39080
rect 26660 39040 26666 39052
rect 27157 39049 27169 39052
rect 27203 39049 27215 39083
rect 27157 39043 27215 39049
rect 27338 39040 27344 39092
rect 27396 39080 27402 39092
rect 27396 39052 28856 39080
rect 27396 39040 27402 39052
rect 25590 38972 25596 39024
rect 25648 39012 25654 39024
rect 25648 38984 26004 39012
rect 25648 38972 25654 38984
rect 25866 38904 25872 38956
rect 25924 38904 25930 38956
rect 25976 38944 26004 38984
rect 26145 38947 26203 38953
rect 26145 38944 26157 38947
rect 25976 38916 26157 38944
rect 26145 38913 26157 38916
rect 26191 38913 26203 38947
rect 26145 38907 26203 38913
rect 26283 38947 26341 38953
rect 26283 38913 26295 38947
rect 26329 38944 26341 38947
rect 26602 38944 26608 38956
rect 26329 38916 26608 38944
rect 26329 38913 26341 38916
rect 26283 38907 26341 38913
rect 26602 38904 26608 38916
rect 26660 38904 26666 38956
rect 26786 38904 26792 38956
rect 26844 38944 26850 38956
rect 26844 38916 27292 38944
rect 26844 38904 26850 38916
rect 25455 38848 25544 38876
rect 25455 38845 25467 38848
rect 25409 38839 25467 38845
rect 26418 38836 26424 38888
rect 26476 38836 26482 38888
rect 27264 38876 27292 38916
rect 28828 38885 28856 39052
rect 29454 39040 29460 39092
rect 29512 39080 29518 39092
rect 29549 39083 29607 39089
rect 29549 39080 29561 39083
rect 29512 39052 29561 39080
rect 29512 39040 29518 39052
rect 29549 39049 29561 39052
rect 29595 39049 29607 39083
rect 29549 39043 29607 39049
rect 30190 39040 30196 39092
rect 30248 39040 30254 39092
rect 28902 38972 28908 39024
rect 28960 39012 28966 39024
rect 29733 39015 29791 39021
rect 29733 39012 29745 39015
rect 28960 38984 29745 39012
rect 28960 38972 28966 38984
rect 29733 38981 29745 38984
rect 29779 38981 29791 39015
rect 29733 38975 29791 38981
rect 28270 38879 28328 38885
rect 28270 38876 28282 38879
rect 27264 38848 28282 38876
rect 28270 38845 28282 38848
rect 28316 38845 28328 38879
rect 28270 38839 28328 38845
rect 28537 38879 28595 38885
rect 28537 38845 28549 38879
rect 28583 38876 28595 38879
rect 28721 38879 28779 38885
rect 28721 38876 28733 38879
rect 28583 38848 28733 38876
rect 28583 38845 28595 38848
rect 28537 38839 28595 38845
rect 28721 38845 28733 38848
rect 28767 38845 28779 38879
rect 28721 38839 28779 38845
rect 28813 38879 28871 38885
rect 28813 38845 28825 38879
rect 28859 38876 28871 38879
rect 29270 38876 29276 38888
rect 28859 38848 29276 38876
rect 28859 38845 28871 38848
rect 28813 38839 28871 38845
rect 29270 38836 29276 38848
rect 29328 38836 29334 38888
rect 29638 38836 29644 38888
rect 29696 38876 29702 38888
rect 30193 38879 30251 38885
rect 30193 38876 30205 38879
rect 29696 38848 30205 38876
rect 29696 38836 29702 38848
rect 30193 38845 30205 38848
rect 30239 38845 30251 38879
rect 30193 38839 30251 38845
rect 30374 38836 30380 38888
rect 30432 38836 30438 38888
rect 18472 38780 20116 38808
rect 18472 38768 18478 38780
rect 20346 38768 20352 38820
rect 20404 38808 20410 38820
rect 20441 38811 20499 38817
rect 20441 38808 20453 38811
rect 20404 38780 20453 38808
rect 20404 38768 20410 38780
rect 20441 38777 20453 38780
rect 20487 38777 20499 38811
rect 28074 38808 28080 38820
rect 20441 38771 20499 38777
rect 26896 38780 28080 38808
rect 8478 38700 8484 38752
rect 8536 38700 8542 38752
rect 9677 38743 9735 38749
rect 9677 38709 9689 38743
rect 9723 38740 9735 38743
rect 9858 38740 9864 38752
rect 9723 38712 9864 38740
rect 9723 38709 9735 38712
rect 9677 38703 9735 38709
rect 9858 38700 9864 38712
rect 9916 38700 9922 38752
rect 12529 38743 12587 38749
rect 12529 38709 12541 38743
rect 12575 38740 12587 38743
rect 14090 38740 14096 38752
rect 12575 38712 14096 38740
rect 12575 38709 12587 38712
rect 12529 38703 12587 38709
rect 14090 38700 14096 38712
rect 14148 38700 14154 38752
rect 15470 38700 15476 38752
rect 15528 38740 15534 38752
rect 15933 38743 15991 38749
rect 15933 38740 15945 38743
rect 15528 38712 15945 38740
rect 15528 38700 15534 38712
rect 15933 38709 15945 38712
rect 15979 38709 15991 38743
rect 15933 38703 15991 38709
rect 16206 38700 16212 38752
rect 16264 38700 16270 38752
rect 16666 38700 16672 38752
rect 16724 38740 16730 38752
rect 16761 38743 16819 38749
rect 16761 38740 16773 38743
rect 16724 38712 16773 38740
rect 16724 38700 16730 38712
rect 16761 38709 16773 38712
rect 16807 38709 16819 38743
rect 16761 38703 16819 38709
rect 16850 38700 16856 38752
rect 16908 38700 16914 38752
rect 19702 38700 19708 38752
rect 19760 38740 19766 38752
rect 19889 38743 19947 38749
rect 19889 38740 19901 38743
rect 19760 38712 19901 38740
rect 19760 38700 19766 38712
rect 19889 38709 19901 38712
rect 19935 38709 19947 38743
rect 19889 38703 19947 38709
rect 20162 38700 20168 38752
rect 20220 38700 20226 38752
rect 23842 38700 23848 38752
rect 23900 38740 23906 38752
rect 26418 38740 26424 38752
rect 23900 38712 26424 38740
rect 23900 38700 23906 38712
rect 26418 38700 26424 38712
rect 26476 38740 26482 38752
rect 26896 38740 26924 38780
rect 28074 38768 28080 38780
rect 28132 38768 28138 38820
rect 29178 38768 29184 38820
rect 29236 38808 29242 38820
rect 29365 38811 29423 38817
rect 29365 38808 29377 38811
rect 29236 38780 29377 38808
rect 29236 38768 29242 38780
rect 29365 38777 29377 38780
rect 29411 38777 29423 38811
rect 30558 38808 30564 38820
rect 29365 38771 29423 38777
rect 29656 38780 30564 38808
rect 26476 38712 26924 38740
rect 26476 38700 26482 38712
rect 26970 38700 26976 38752
rect 27028 38740 27034 38752
rect 27065 38743 27123 38749
rect 27065 38740 27077 38743
rect 27028 38712 27077 38740
rect 27028 38700 27034 38712
rect 27065 38709 27077 38712
rect 27111 38709 27123 38743
rect 28092 38740 28120 38768
rect 28810 38740 28816 38752
rect 28092 38712 28816 38740
rect 27065 38703 27123 38709
rect 28810 38700 28816 38712
rect 28868 38700 28874 38752
rect 29570 38743 29628 38749
rect 29570 38709 29582 38743
rect 29616 38740 29628 38743
rect 29656 38740 29684 38780
rect 30558 38768 30564 38780
rect 30616 38768 30622 38820
rect 29616 38712 29684 38740
rect 29616 38709 29628 38712
rect 29570 38703 29628 38709
rect 552 38650 31648 38672
rect 552 38598 4322 38650
rect 4374 38598 4386 38650
rect 4438 38598 4450 38650
rect 4502 38598 4514 38650
rect 4566 38598 4578 38650
rect 4630 38598 12096 38650
rect 12148 38598 12160 38650
rect 12212 38598 12224 38650
rect 12276 38598 12288 38650
rect 12340 38598 12352 38650
rect 12404 38598 19870 38650
rect 19922 38598 19934 38650
rect 19986 38598 19998 38650
rect 20050 38598 20062 38650
rect 20114 38598 20126 38650
rect 20178 38598 27644 38650
rect 27696 38598 27708 38650
rect 27760 38598 27772 38650
rect 27824 38598 27836 38650
rect 27888 38598 27900 38650
rect 27952 38598 31648 38650
rect 552 38576 31648 38598
rect 9493 38539 9551 38545
rect 9493 38505 9505 38539
rect 9539 38536 9551 38539
rect 9582 38536 9588 38548
rect 9539 38508 9588 38536
rect 9539 38505 9551 38508
rect 9493 38499 9551 38505
rect 9582 38496 9588 38508
rect 9640 38496 9646 38548
rect 14353 38539 14411 38545
rect 14353 38505 14365 38539
rect 14399 38536 14411 38539
rect 14645 38539 14703 38545
rect 14645 38536 14657 38539
rect 14399 38508 14657 38536
rect 14399 38505 14411 38508
rect 14353 38499 14411 38505
rect 14645 38505 14657 38508
rect 14691 38505 14703 38539
rect 14645 38499 14703 38505
rect 15013 38539 15071 38545
rect 15013 38505 15025 38539
rect 15059 38536 15071 38539
rect 15102 38536 15108 38548
rect 15059 38508 15108 38536
rect 15059 38505 15071 38508
rect 15013 38499 15071 38505
rect 15102 38496 15108 38508
rect 15160 38496 15166 38548
rect 15289 38539 15347 38545
rect 15289 38505 15301 38539
rect 15335 38536 15347 38539
rect 15654 38536 15660 38548
rect 15335 38508 15660 38536
rect 15335 38505 15347 38508
rect 15289 38499 15347 38505
rect 15654 38496 15660 38508
rect 15712 38496 15718 38548
rect 16390 38496 16396 38548
rect 16448 38536 16454 38548
rect 17497 38539 17555 38545
rect 17497 38536 17509 38539
rect 16448 38508 17509 38536
rect 16448 38496 16454 38508
rect 17497 38505 17509 38508
rect 17543 38505 17555 38539
rect 22278 38536 22284 38548
rect 17497 38499 17555 38505
rect 18800 38508 22284 38536
rect 8478 38468 8484 38480
rect 8128 38440 8484 38468
rect 8128 38409 8156 38440
rect 8478 38428 8484 38440
rect 8536 38428 8542 38480
rect 11330 38428 11336 38480
rect 11388 38468 11394 38480
rect 11882 38468 11888 38480
rect 11388 38440 11560 38468
rect 11388 38428 11394 38440
rect 8113 38403 8171 38409
rect 8113 38369 8125 38403
rect 8159 38369 8171 38403
rect 8113 38363 8171 38369
rect 8380 38403 8438 38409
rect 8380 38369 8392 38403
rect 8426 38400 8438 38403
rect 8426 38372 9628 38400
rect 8426 38369 8438 38372
rect 8380 38363 8438 38369
rect 9600 38341 9628 38372
rect 9858 38360 9864 38412
rect 9916 38360 9922 38412
rect 9953 38403 10011 38409
rect 9953 38369 9965 38403
rect 9999 38369 10011 38403
rect 9953 38363 10011 38369
rect 9585 38335 9643 38341
rect 9585 38301 9597 38335
rect 9631 38301 9643 38335
rect 9968 38332 9996 38363
rect 10042 38360 10048 38412
rect 10100 38360 10106 38412
rect 10226 38360 10232 38412
rect 10284 38360 10290 38412
rect 11532 38409 11560 38440
rect 11624 38440 11888 38468
rect 11624 38409 11652 38440
rect 11882 38428 11888 38440
rect 11940 38428 11946 38480
rect 13081 38471 13139 38477
rect 13081 38468 13093 38471
rect 12452 38440 13093 38468
rect 12452 38412 12480 38440
rect 13081 38437 13093 38440
rect 13127 38437 13139 38471
rect 13081 38431 13139 38437
rect 13446 38428 13452 38480
rect 13504 38468 13510 38480
rect 14553 38471 14611 38477
rect 13504 38440 13952 38468
rect 13504 38428 13510 38440
rect 11425 38403 11483 38409
rect 11425 38369 11437 38403
rect 11471 38369 11483 38403
rect 11425 38363 11483 38369
rect 11517 38403 11575 38409
rect 11517 38369 11529 38403
rect 11563 38369 11575 38403
rect 11517 38363 11575 38369
rect 11609 38403 11667 38409
rect 11609 38369 11621 38403
rect 11655 38369 11667 38403
rect 11609 38363 11667 38369
rect 11793 38403 11851 38409
rect 11793 38369 11805 38403
rect 11839 38400 11851 38403
rect 11839 38372 12020 38400
rect 11839 38369 11851 38372
rect 11793 38363 11851 38369
rect 10502 38332 10508 38344
rect 9585 38295 9643 38301
rect 9876 38304 10508 38332
rect 9876 38276 9904 38304
rect 10502 38292 10508 38304
rect 10560 38332 10566 38344
rect 10962 38332 10968 38344
rect 10560 38304 10968 38332
rect 10560 38292 10566 38304
rect 10962 38292 10968 38304
rect 11020 38292 11026 38344
rect 11440 38332 11468 38363
rect 11885 38335 11943 38341
rect 11885 38332 11897 38335
rect 11440 38304 11897 38332
rect 11885 38301 11897 38304
rect 11931 38301 11943 38335
rect 11885 38295 11943 38301
rect 9858 38224 9864 38276
rect 9916 38224 9922 38276
rect 10226 38224 10232 38276
rect 10284 38264 10290 38276
rect 11992 38264 12020 38372
rect 12434 38360 12440 38412
rect 12492 38360 12498 38412
rect 12989 38403 13047 38409
rect 12989 38369 13001 38403
rect 13035 38400 13047 38403
rect 13725 38403 13783 38409
rect 13725 38400 13737 38403
rect 13035 38372 13737 38400
rect 13035 38369 13047 38372
rect 12989 38363 13047 38369
rect 13725 38369 13737 38372
rect 13771 38369 13783 38403
rect 13725 38363 13783 38369
rect 13262 38292 13268 38344
rect 13320 38292 13326 38344
rect 13740 38332 13768 38363
rect 13814 38360 13820 38412
rect 13872 38360 13878 38412
rect 13924 38409 13952 38440
rect 14553 38437 14565 38471
rect 14599 38468 14611 38471
rect 15194 38468 15200 38480
rect 14599 38440 15200 38468
rect 14599 38437 14611 38440
rect 14553 38431 14611 38437
rect 15194 38428 15200 38440
rect 15252 38428 15258 38480
rect 13909 38403 13967 38409
rect 13909 38369 13921 38403
rect 13955 38369 13967 38403
rect 13909 38363 13967 38369
rect 14090 38360 14096 38412
rect 14148 38360 14154 38412
rect 14829 38403 14887 38409
rect 14829 38369 14841 38403
rect 14875 38400 14887 38403
rect 14918 38400 14924 38412
rect 14875 38372 14924 38400
rect 14875 38369 14887 38372
rect 14829 38363 14887 38369
rect 14844 38332 14872 38363
rect 14918 38360 14924 38372
rect 14976 38360 14982 38412
rect 15105 38403 15163 38409
rect 15105 38369 15117 38403
rect 15151 38400 15163 38403
rect 15473 38403 15531 38409
rect 15473 38400 15485 38403
rect 15151 38372 15485 38400
rect 15151 38369 15163 38372
rect 15105 38363 15163 38369
rect 15473 38369 15485 38372
rect 15519 38400 15531 38403
rect 16022 38400 16028 38412
rect 15519 38372 16028 38400
rect 15519 38369 15531 38372
rect 15473 38363 15531 38369
rect 16022 38360 16028 38372
rect 16080 38360 16086 38412
rect 16117 38403 16175 38409
rect 16117 38369 16129 38403
rect 16163 38400 16175 38403
rect 16206 38400 16212 38412
rect 16163 38372 16212 38400
rect 16163 38369 16175 38372
rect 16117 38363 16175 38369
rect 16206 38360 16212 38372
rect 16264 38360 16270 38412
rect 17678 38360 17684 38412
rect 17736 38400 17742 38412
rect 17865 38403 17923 38409
rect 17865 38400 17877 38403
rect 17736 38372 17877 38400
rect 17736 38360 17742 38372
rect 17865 38369 17877 38372
rect 17911 38369 17923 38403
rect 17865 38363 17923 38369
rect 18049 38403 18107 38409
rect 18049 38369 18061 38403
rect 18095 38400 18107 38403
rect 18414 38400 18420 38412
rect 18095 38372 18420 38400
rect 18095 38369 18107 38372
rect 18049 38363 18107 38369
rect 13740 38304 14872 38332
rect 15749 38335 15807 38341
rect 15749 38301 15761 38335
rect 15795 38301 15807 38335
rect 15749 38295 15807 38301
rect 10284 38236 12020 38264
rect 12621 38267 12679 38273
rect 10284 38224 10290 38236
rect 12621 38233 12633 38267
rect 12667 38264 12679 38267
rect 12986 38264 12992 38276
rect 12667 38236 12992 38264
rect 12667 38233 12679 38236
rect 12621 38227 12679 38233
rect 12986 38224 12992 38236
rect 13044 38224 13050 38276
rect 15764 38264 15792 38295
rect 15930 38292 15936 38344
rect 15988 38332 15994 38344
rect 16393 38335 16451 38341
rect 16393 38332 16405 38335
rect 15988 38304 16405 38332
rect 15988 38292 15994 38304
rect 16393 38301 16405 38304
rect 16439 38301 16451 38335
rect 16393 38295 16451 38301
rect 17494 38292 17500 38344
rect 17552 38332 17558 38344
rect 18064 38332 18092 38363
rect 18414 38360 18420 38372
rect 18472 38360 18478 38412
rect 18800 38409 18828 38508
rect 22278 38496 22284 38508
rect 22336 38496 22342 38548
rect 23566 38496 23572 38548
rect 23624 38496 23630 38548
rect 28445 38539 28503 38545
rect 28445 38505 28457 38539
rect 28491 38536 28503 38539
rect 28534 38536 28540 38548
rect 28491 38508 28540 38536
rect 28491 38505 28503 38508
rect 28445 38499 28503 38505
rect 28534 38496 28540 38508
rect 28592 38496 28598 38548
rect 20806 38468 20812 38480
rect 19904 38440 20812 38468
rect 18785 38403 18843 38409
rect 18785 38369 18797 38403
rect 18831 38369 18843 38403
rect 18785 38363 18843 38369
rect 19058 38360 19064 38412
rect 19116 38400 19122 38412
rect 19153 38403 19211 38409
rect 19153 38400 19165 38403
rect 19116 38372 19165 38400
rect 19116 38360 19122 38372
rect 19153 38369 19165 38372
rect 19199 38369 19211 38403
rect 19153 38363 19211 38369
rect 19337 38403 19395 38409
rect 19337 38369 19349 38403
rect 19383 38369 19395 38403
rect 19337 38363 19395 38369
rect 17552 38304 18092 38332
rect 18693 38335 18751 38341
rect 17552 38292 17558 38304
rect 18693 38301 18705 38335
rect 18739 38301 18751 38335
rect 18693 38295 18751 38301
rect 18877 38335 18935 38341
rect 18877 38301 18889 38335
rect 18923 38301 18935 38335
rect 18877 38295 18935 38301
rect 16114 38264 16120 38276
rect 15764 38236 16120 38264
rect 16114 38224 16120 38236
rect 16172 38224 16178 38276
rect 18509 38267 18567 38273
rect 18509 38264 18521 38267
rect 17052 38236 18521 38264
rect 10134 38156 10140 38208
rect 10192 38196 10198 38208
rect 10318 38196 10324 38208
rect 10192 38168 10324 38196
rect 10192 38156 10198 38168
rect 10318 38156 10324 38168
rect 10376 38156 10382 38208
rect 11149 38199 11207 38205
rect 11149 38165 11161 38199
rect 11195 38196 11207 38199
rect 11238 38196 11244 38208
rect 11195 38168 11244 38196
rect 11195 38165 11207 38168
rect 11149 38159 11207 38165
rect 11238 38156 11244 38168
rect 11296 38156 11302 38208
rect 12710 38156 12716 38208
rect 12768 38196 12774 38208
rect 13449 38199 13507 38205
rect 13449 38196 13461 38199
rect 12768 38168 13461 38196
rect 12768 38156 12774 38168
rect 13449 38165 13461 38168
rect 13495 38165 13507 38199
rect 13449 38159 13507 38165
rect 14182 38156 14188 38208
rect 14240 38156 14246 38208
rect 14366 38156 14372 38208
rect 14424 38156 14430 38208
rect 15654 38156 15660 38208
rect 15712 38156 15718 38208
rect 15746 38156 15752 38208
rect 15804 38196 15810 38208
rect 17052 38196 17080 38236
rect 18509 38233 18521 38236
rect 18555 38233 18567 38267
rect 18509 38227 18567 38233
rect 15804 38168 17080 38196
rect 15804 38156 15810 38168
rect 17862 38156 17868 38208
rect 17920 38196 17926 38208
rect 17957 38199 18015 38205
rect 17957 38196 17969 38199
rect 17920 38168 17969 38196
rect 17920 38156 17926 38168
rect 17957 38165 17969 38168
rect 18003 38165 18015 38199
rect 18708 38196 18736 38295
rect 18892 38264 18920 38295
rect 18966 38292 18972 38344
rect 19024 38292 19030 38344
rect 19352 38332 19380 38363
rect 19702 38360 19708 38412
rect 19760 38360 19766 38412
rect 19904 38400 19932 38440
rect 20806 38428 20812 38440
rect 20864 38428 20870 38480
rect 23477 38471 23535 38477
rect 23477 38437 23489 38471
rect 23523 38468 23535 38471
rect 25130 38468 25136 38480
rect 23523 38440 25136 38468
rect 23523 38437 23535 38440
rect 23477 38431 23535 38437
rect 25130 38428 25136 38440
rect 25188 38428 25194 38480
rect 27332 38471 27390 38477
rect 27332 38437 27344 38471
rect 27378 38468 27390 38471
rect 27982 38468 27988 38480
rect 27378 38440 27988 38468
rect 27378 38437 27390 38440
rect 27332 38431 27390 38437
rect 27982 38428 27988 38440
rect 28040 38428 28046 38480
rect 19978 38409 19984 38412
rect 19812 38372 19932 38400
rect 19812 38332 19840 38372
rect 19972 38363 19984 38409
rect 19978 38360 19984 38363
rect 20036 38360 20042 38412
rect 20530 38360 20536 38412
rect 20588 38400 20594 38412
rect 20588 38372 22131 38400
rect 20588 38360 20594 38372
rect 19352 38304 19840 38332
rect 22103 38332 22131 38372
rect 22370 38360 22376 38412
rect 22428 38400 22434 38412
rect 22465 38403 22523 38409
rect 22465 38400 22477 38403
rect 22428 38372 22477 38400
rect 22428 38360 22434 38372
rect 22465 38369 22477 38372
rect 22511 38400 22523 38403
rect 22649 38403 22707 38409
rect 22649 38400 22661 38403
rect 22511 38372 22661 38400
rect 22511 38369 22523 38372
rect 22465 38363 22523 38369
rect 22649 38369 22661 38372
rect 22695 38369 22707 38403
rect 22649 38363 22707 38369
rect 23750 38360 23756 38412
rect 23808 38360 23814 38412
rect 26878 38360 26884 38412
rect 26936 38400 26942 38412
rect 27065 38403 27123 38409
rect 27065 38400 27077 38403
rect 26936 38372 27077 38400
rect 26936 38360 26942 38372
rect 27065 38369 27077 38372
rect 27111 38369 27123 38403
rect 27065 38363 27123 38369
rect 29270 38360 29276 38412
rect 29328 38400 29334 38412
rect 29365 38403 29423 38409
rect 29365 38400 29377 38403
rect 29328 38372 29377 38400
rect 29328 38360 29334 38372
rect 29365 38369 29377 38372
rect 29411 38369 29423 38403
rect 29365 38363 29423 38369
rect 23934 38332 23940 38344
rect 22103 38304 23940 38332
rect 23934 38292 23940 38304
rect 23992 38292 23998 38344
rect 19245 38267 19303 38273
rect 19245 38264 19257 38267
rect 18892 38236 19257 38264
rect 19245 38233 19257 38236
rect 19291 38233 19303 38267
rect 22830 38264 22836 38276
rect 19245 38227 19303 38233
rect 20640 38236 22836 38264
rect 20640 38196 20668 38236
rect 22830 38224 22836 38236
rect 22888 38224 22894 38276
rect 18708 38168 20668 38196
rect 17957 38159 18015 38165
rect 20898 38156 20904 38208
rect 20956 38196 20962 38208
rect 21085 38199 21143 38205
rect 21085 38196 21097 38199
rect 20956 38168 21097 38196
rect 20956 38156 20962 38168
rect 21085 38165 21097 38168
rect 21131 38165 21143 38199
rect 21085 38159 21143 38165
rect 22186 38156 22192 38208
rect 22244 38196 22250 38208
rect 22373 38199 22431 38205
rect 22373 38196 22385 38199
rect 22244 38168 22385 38196
rect 22244 38156 22250 38168
rect 22373 38165 22385 38168
rect 22419 38165 22431 38199
rect 22373 38159 22431 38165
rect 29086 38156 29092 38208
rect 29144 38196 29150 38208
rect 29273 38199 29331 38205
rect 29273 38196 29285 38199
rect 29144 38168 29285 38196
rect 29144 38156 29150 38168
rect 29273 38165 29285 38168
rect 29319 38165 29331 38199
rect 29273 38159 29331 38165
rect 552 38106 31648 38128
rect 552 38054 3662 38106
rect 3714 38054 3726 38106
rect 3778 38054 3790 38106
rect 3842 38054 3854 38106
rect 3906 38054 3918 38106
rect 3970 38054 11436 38106
rect 11488 38054 11500 38106
rect 11552 38054 11564 38106
rect 11616 38054 11628 38106
rect 11680 38054 11692 38106
rect 11744 38054 19210 38106
rect 19262 38054 19274 38106
rect 19326 38054 19338 38106
rect 19390 38054 19402 38106
rect 19454 38054 19466 38106
rect 19518 38054 26984 38106
rect 27036 38054 27048 38106
rect 27100 38054 27112 38106
rect 27164 38054 27176 38106
rect 27228 38054 27240 38106
rect 27292 38054 31648 38106
rect 552 38032 31648 38054
rect 9674 37952 9680 38004
rect 9732 37952 9738 38004
rect 9876 37964 10916 37992
rect 8294 37884 8300 37936
rect 8352 37924 8358 37936
rect 9876 37924 9904 37964
rect 8352 37896 9904 37924
rect 8352 37884 8358 37896
rect 10134 37856 10140 37868
rect 9416 37828 10140 37856
rect 9416 37729 9444 37828
rect 10134 37816 10140 37828
rect 10192 37816 10198 37868
rect 10318 37816 10324 37868
rect 10376 37816 10382 37868
rect 10888 37800 10916 37964
rect 12434 37952 12440 38004
rect 12492 37992 12498 38004
rect 12529 37995 12587 38001
rect 12529 37992 12541 37995
rect 12492 37964 12541 37992
rect 12492 37952 12498 37964
rect 12529 37961 12541 37964
rect 12575 37961 12587 37995
rect 12529 37955 12587 37961
rect 13078 37952 13084 38004
rect 13136 37992 13142 38004
rect 13173 37995 13231 38001
rect 13173 37992 13185 37995
rect 13136 37964 13185 37992
rect 13136 37952 13142 37964
rect 13173 37961 13185 37964
rect 13219 37961 13231 37995
rect 13173 37955 13231 37961
rect 14918 37952 14924 38004
rect 14976 37992 14982 38004
rect 15197 37995 15255 38001
rect 15197 37992 15209 37995
rect 14976 37964 15209 37992
rect 14976 37952 14982 37964
rect 15197 37961 15209 37964
rect 15243 37961 15255 37995
rect 15197 37955 15255 37961
rect 15930 37952 15936 38004
rect 15988 37952 15994 38004
rect 16850 37952 16856 38004
rect 16908 37992 16914 38004
rect 17221 37995 17279 38001
rect 17221 37992 17233 37995
rect 16908 37964 17233 37992
rect 16908 37952 16914 37964
rect 17221 37961 17233 37964
rect 17267 37961 17279 37995
rect 18046 37992 18052 38004
rect 17221 37955 17279 37961
rect 17604 37964 18052 37992
rect 12894 37924 12900 37936
rect 12176 37896 12900 37924
rect 9490 37748 9496 37800
rect 9548 37788 9554 37800
rect 10045 37791 10103 37797
rect 10045 37788 10057 37791
rect 9548 37760 10057 37788
rect 9548 37748 9554 37760
rect 10045 37757 10057 37760
rect 10091 37757 10103 37791
rect 10045 37751 10103 37757
rect 10870 37748 10876 37800
rect 10928 37748 10934 37800
rect 10965 37791 11023 37797
rect 10965 37757 10977 37791
rect 11011 37788 11023 37791
rect 11149 37791 11207 37797
rect 11149 37788 11161 37791
rect 11011 37760 11161 37788
rect 11011 37757 11023 37760
rect 10965 37751 11023 37757
rect 11149 37757 11161 37760
rect 11195 37757 11207 37791
rect 11149 37751 11207 37757
rect 11238 37748 11244 37800
rect 11296 37788 11302 37800
rect 11405 37791 11463 37797
rect 11405 37788 11417 37791
rect 11296 37760 11417 37788
rect 11296 37748 11302 37760
rect 11405 37757 11417 37760
rect 11451 37757 11463 37791
rect 11405 37751 11463 37757
rect 9401 37723 9459 37729
rect 9401 37689 9413 37723
rect 9447 37689 9459 37723
rect 9401 37683 9459 37689
rect 9585 37723 9643 37729
rect 9585 37689 9597 37723
rect 9631 37720 9643 37723
rect 12176 37720 12204 37896
rect 12894 37884 12900 37896
rect 12952 37884 12958 37936
rect 16482 37884 16488 37936
rect 16540 37924 16546 37936
rect 17604 37924 17632 37964
rect 18046 37952 18052 37964
rect 18104 37992 18110 38004
rect 18417 37995 18475 38001
rect 18417 37992 18429 37995
rect 18104 37964 18429 37992
rect 18104 37952 18110 37964
rect 18417 37961 18429 37964
rect 18463 37992 18475 37995
rect 18874 37992 18880 38004
rect 18463 37964 18880 37992
rect 18463 37961 18475 37964
rect 18417 37955 18475 37961
rect 18874 37952 18880 37964
rect 18932 37952 18938 38004
rect 19797 37995 19855 38001
rect 19797 37961 19809 37995
rect 19843 37992 19855 37995
rect 19978 37992 19984 38004
rect 19843 37964 19984 37992
rect 19843 37961 19855 37964
rect 19797 37955 19855 37961
rect 19978 37952 19984 37964
rect 20036 37952 20042 38004
rect 20438 37952 20444 38004
rect 20496 37992 20502 38004
rect 20714 37992 20720 38004
rect 20496 37964 20720 37992
rect 20496 37952 20502 37964
rect 20714 37952 20720 37964
rect 20772 37952 20778 38004
rect 23290 37992 23296 38004
rect 22066 37964 23296 37992
rect 16540 37896 17632 37924
rect 16540 37884 16546 37896
rect 17678 37884 17684 37936
rect 17736 37924 17742 37936
rect 22066 37924 22094 37964
rect 23290 37952 23296 37964
rect 23348 37952 23354 38004
rect 23569 37995 23627 38001
rect 23569 37961 23581 37995
rect 23615 37992 23627 37995
rect 24026 37992 24032 38004
rect 23615 37964 24032 37992
rect 23615 37961 23627 37964
rect 23569 37955 23627 37961
rect 24026 37952 24032 37964
rect 24084 37992 24090 38004
rect 25866 37992 25872 38004
rect 24084 37964 25872 37992
rect 24084 37952 24090 37964
rect 25866 37952 25872 37964
rect 25924 37952 25930 38004
rect 17736 37896 22094 37924
rect 17736 37884 17742 37896
rect 13633 37859 13691 37865
rect 13633 37825 13645 37859
rect 13679 37856 13691 37859
rect 13817 37859 13875 37865
rect 13817 37856 13829 37859
rect 13679 37828 13829 37856
rect 13679 37825 13691 37828
rect 13633 37819 13691 37825
rect 13817 37825 13829 37828
rect 13863 37825 13875 37859
rect 13817 37819 13875 37825
rect 15212 37828 16988 37856
rect 12621 37791 12679 37797
rect 12621 37757 12633 37791
rect 12667 37757 12679 37791
rect 12621 37751 12679 37757
rect 12636 37720 12664 37751
rect 12710 37748 12716 37800
rect 12768 37748 12774 37800
rect 12802 37748 12808 37800
rect 12860 37788 12866 37800
rect 12897 37791 12955 37797
rect 12897 37788 12909 37791
rect 12860 37760 12909 37788
rect 12860 37748 12866 37760
rect 12897 37757 12909 37760
rect 12943 37757 12955 37791
rect 12897 37751 12955 37757
rect 12986 37748 12992 37800
rect 13044 37748 13050 37800
rect 13725 37791 13783 37797
rect 13725 37757 13737 37791
rect 13771 37788 13783 37791
rect 15212 37788 15240 37828
rect 16960 37800 16988 37828
rect 17862 37816 17868 37868
rect 17920 37816 17926 37868
rect 19334 37816 19340 37868
rect 19392 37816 19398 37868
rect 13771 37760 15240 37788
rect 15289 37791 15347 37797
rect 13771 37757 13783 37760
rect 13725 37751 13783 37757
rect 15289 37757 15301 37791
rect 15335 37788 15347 37791
rect 15378 37788 15384 37800
rect 15335 37760 15384 37788
rect 15335 37757 15347 37760
rect 15289 37751 15347 37757
rect 15378 37748 15384 37760
rect 15436 37748 15442 37800
rect 15470 37748 15476 37800
rect 15528 37748 15534 37800
rect 15562 37748 15568 37800
rect 15620 37748 15626 37800
rect 15657 37791 15715 37797
rect 15657 37757 15669 37791
rect 15703 37788 15715 37791
rect 15838 37788 15844 37800
rect 15703 37760 15844 37788
rect 15703 37757 15715 37760
rect 15657 37751 15715 37757
rect 15838 37748 15844 37760
rect 15896 37788 15902 37800
rect 16206 37788 16212 37800
rect 15896 37760 16212 37788
rect 15896 37748 15902 37760
rect 16206 37748 16212 37760
rect 16264 37748 16270 37800
rect 16942 37748 16948 37800
rect 17000 37748 17006 37800
rect 18233 37791 18291 37797
rect 18233 37757 18245 37791
rect 18279 37757 18291 37791
rect 18233 37751 18291 37757
rect 13906 37720 13912 37732
rect 9631 37692 12204 37720
rect 12406 37692 13912 37720
rect 9631 37689 9643 37692
rect 9585 37683 9643 37689
rect 9217 37655 9275 37661
rect 9217 37621 9229 37655
rect 9263 37652 9275 37655
rect 9490 37652 9496 37664
rect 9263 37624 9496 37652
rect 9263 37621 9275 37624
rect 9217 37615 9275 37621
rect 9490 37612 9496 37624
rect 9548 37612 9554 37664
rect 10594 37612 10600 37664
rect 10652 37652 10658 37664
rect 12406 37652 12434 37692
rect 13906 37680 13912 37692
rect 13964 37680 13970 37732
rect 14084 37723 14142 37729
rect 14084 37689 14096 37723
rect 14130 37720 14142 37723
rect 14182 37720 14188 37732
rect 14130 37692 14188 37720
rect 14130 37689 14142 37692
rect 14084 37683 14142 37689
rect 14182 37680 14188 37692
rect 14240 37680 14246 37732
rect 10652 37624 12434 37652
rect 15396 37652 15424 37748
rect 16390 37680 16396 37732
rect 16448 37720 16454 37732
rect 17681 37723 17739 37729
rect 17681 37720 17693 37723
rect 16448 37692 17693 37720
rect 16448 37680 16454 37692
rect 17681 37689 17693 37692
rect 17727 37689 17739 37723
rect 17681 37683 17739 37689
rect 16850 37652 16856 37664
rect 15396 37624 16856 37652
rect 10652 37612 10658 37624
rect 16850 37612 16856 37624
rect 16908 37612 16914 37664
rect 17589 37655 17647 37661
rect 17589 37621 17601 37655
rect 17635 37652 17647 37655
rect 17862 37652 17868 37664
rect 17635 37624 17868 37652
rect 17635 37621 17647 37624
rect 17589 37615 17647 37621
rect 17862 37612 17868 37624
rect 17920 37612 17926 37664
rect 18248 37652 18276 37751
rect 18322 37748 18328 37800
rect 18380 37788 18386 37800
rect 18966 37788 18972 37800
rect 18380 37760 18972 37788
rect 18380 37748 18386 37760
rect 18966 37748 18972 37760
rect 19024 37748 19030 37800
rect 19521 37791 19579 37797
rect 19521 37757 19533 37791
rect 19567 37788 19579 37791
rect 19720 37788 19748 37896
rect 19794 37816 19800 37868
rect 19852 37856 19858 37868
rect 19852 37828 21220 37856
rect 19852 37816 19858 37828
rect 19567 37760 19748 37788
rect 19567 37757 19579 37760
rect 19521 37751 19579 37757
rect 20070 37748 20076 37800
rect 20128 37748 20134 37800
rect 20162 37748 20168 37800
rect 20220 37748 20226 37800
rect 20257 37791 20315 37797
rect 20257 37757 20269 37791
rect 20303 37788 20315 37791
rect 20346 37788 20352 37800
rect 20303 37760 20352 37788
rect 20303 37757 20315 37760
rect 20257 37751 20315 37757
rect 20346 37748 20352 37760
rect 20404 37748 20410 37800
rect 20441 37791 20499 37797
rect 20441 37757 20453 37791
rect 20487 37788 20499 37791
rect 20530 37788 20536 37800
rect 20487 37760 20536 37788
rect 20487 37757 20499 37760
rect 20441 37751 20499 37757
rect 18782 37680 18788 37732
rect 18840 37680 18846 37732
rect 18874 37680 18880 37732
rect 18932 37680 18938 37732
rect 19610 37680 19616 37732
rect 19668 37720 19674 37732
rect 20456 37720 20484 37751
rect 20530 37748 20536 37760
rect 20588 37748 20594 37800
rect 20898 37748 20904 37800
rect 20956 37748 20962 37800
rect 21192 37788 21220 37828
rect 21266 37816 21272 37868
rect 21324 37856 21330 37868
rect 21913 37859 21971 37865
rect 21913 37856 21925 37859
rect 21324 37828 21925 37856
rect 21324 37816 21330 37828
rect 21913 37825 21925 37828
rect 21959 37825 21971 37859
rect 21913 37819 21971 37825
rect 22186 37816 22192 37868
rect 22244 37816 22250 37868
rect 29086 37816 29092 37868
rect 29144 37816 29150 37868
rect 31110 37856 31116 37868
rect 30392 37828 31116 37856
rect 22005 37791 22063 37797
rect 22005 37788 22017 37791
rect 21192 37760 22017 37788
rect 22005 37757 22017 37760
rect 22051 37788 22063 37791
rect 22278 37788 22284 37800
rect 22051 37760 22284 37788
rect 22051 37757 22063 37760
rect 22005 37751 22063 37757
rect 22278 37748 22284 37760
rect 22336 37748 22342 37800
rect 24946 37748 24952 37800
rect 25004 37748 25010 37800
rect 29356 37791 29414 37797
rect 29356 37757 29368 37791
rect 29402 37788 29414 37791
rect 30392 37788 30420 37828
rect 31110 37816 31116 37828
rect 31168 37816 31174 37868
rect 30653 37791 30711 37797
rect 30653 37788 30665 37791
rect 29402 37760 30420 37788
rect 30484 37760 30665 37788
rect 29402 37757 29414 37760
rect 29356 37751 29414 37757
rect 19668 37692 20484 37720
rect 19668 37680 19674 37692
rect 21634 37680 21640 37732
rect 21692 37680 21698 37732
rect 22456 37723 22514 37729
rect 22456 37689 22468 37723
rect 22502 37720 22514 37723
rect 23382 37720 23388 37732
rect 22502 37692 23388 37720
rect 22502 37689 22514 37692
rect 22456 37683 22514 37689
rect 23382 37680 23388 37692
rect 23440 37680 23446 37732
rect 30484 37664 30512 37760
rect 30653 37757 30665 37760
rect 30699 37757 30711 37791
rect 30653 37751 30711 37757
rect 19518 37652 19524 37664
rect 18248 37624 19524 37652
rect 19518 37612 19524 37624
rect 19576 37612 19582 37664
rect 20622 37612 20628 37664
rect 20680 37612 20686 37664
rect 21545 37655 21603 37661
rect 21545 37621 21557 37655
rect 21591 37652 21603 37655
rect 21818 37652 21824 37664
rect 21591 37624 21824 37652
rect 21591 37621 21603 37624
rect 21545 37615 21603 37621
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 30466 37612 30472 37664
rect 30524 37612 30530 37664
rect 31297 37655 31355 37661
rect 31297 37621 31309 37655
rect 31343 37652 31355 37655
rect 31343 37624 31708 37652
rect 31343 37621 31355 37624
rect 31297 37615 31355 37621
rect 552 37562 31648 37584
rect 552 37510 4322 37562
rect 4374 37510 4386 37562
rect 4438 37510 4450 37562
rect 4502 37510 4514 37562
rect 4566 37510 4578 37562
rect 4630 37510 12096 37562
rect 12148 37510 12160 37562
rect 12212 37510 12224 37562
rect 12276 37510 12288 37562
rect 12340 37510 12352 37562
rect 12404 37510 19870 37562
rect 19922 37510 19934 37562
rect 19986 37510 19998 37562
rect 20050 37510 20062 37562
rect 20114 37510 20126 37562
rect 20178 37510 27644 37562
rect 27696 37510 27708 37562
rect 27760 37510 27772 37562
rect 27824 37510 27836 37562
rect 27888 37510 27900 37562
rect 27952 37510 31648 37562
rect 552 37488 31648 37510
rect 8849 37451 8907 37457
rect 8849 37417 8861 37451
rect 8895 37448 8907 37451
rect 9122 37448 9128 37460
rect 8895 37420 9128 37448
rect 8895 37417 8907 37420
rect 8849 37411 8907 37417
rect 9122 37408 9128 37420
rect 9180 37408 9186 37460
rect 9950 37448 9956 37460
rect 9232 37420 9956 37448
rect 9122 37272 9128 37324
rect 9180 37272 9186 37324
rect 9232 37321 9260 37420
rect 9950 37408 9956 37420
rect 10008 37408 10014 37460
rect 10410 37408 10416 37460
rect 10468 37408 10474 37460
rect 14093 37451 14151 37457
rect 14093 37417 14105 37451
rect 14139 37448 14151 37451
rect 14366 37448 14372 37460
rect 14139 37420 14372 37448
rect 14139 37417 14151 37420
rect 14093 37411 14151 37417
rect 14366 37408 14372 37420
rect 14424 37408 14430 37460
rect 15654 37408 15660 37460
rect 15712 37448 15718 37460
rect 15933 37451 15991 37457
rect 15933 37448 15945 37451
rect 15712 37420 15945 37448
rect 15712 37408 15718 37420
rect 15933 37417 15945 37420
rect 15979 37448 15991 37451
rect 16482 37448 16488 37460
rect 15979 37420 16488 37448
rect 15979 37417 15991 37420
rect 15933 37411 15991 37417
rect 16482 37408 16488 37420
rect 16540 37408 16546 37460
rect 20346 37408 20352 37460
rect 20404 37408 20410 37460
rect 20441 37451 20499 37457
rect 20441 37417 20453 37451
rect 20487 37448 20499 37451
rect 20487 37420 21568 37448
rect 20487 37417 20499 37420
rect 20441 37411 20499 37417
rect 9766 37380 9772 37392
rect 9324 37352 9772 37380
rect 9324 37321 9352 37352
rect 9766 37340 9772 37352
rect 9824 37340 9830 37392
rect 10428 37380 10456 37408
rect 10336 37352 10456 37380
rect 10336 37324 10364 37352
rect 10870 37340 10876 37392
rect 10928 37380 10934 37392
rect 14277 37383 14335 37389
rect 14277 37380 14289 37383
rect 10928 37352 14289 37380
rect 10928 37340 10934 37352
rect 14277 37349 14289 37352
rect 14323 37349 14335 37383
rect 16117 37383 16175 37389
rect 16117 37380 16129 37383
rect 14277 37343 14335 37349
rect 15212 37352 16129 37380
rect 15212 37324 15240 37352
rect 16117 37349 16129 37352
rect 16163 37349 16175 37383
rect 16117 37343 16175 37349
rect 16500 37352 18276 37380
rect 9217 37315 9275 37321
rect 9217 37281 9229 37315
rect 9263 37281 9275 37315
rect 9217 37275 9275 37281
rect 9309 37315 9367 37321
rect 9309 37281 9321 37315
rect 9355 37281 9367 37315
rect 9309 37275 9367 37281
rect 9490 37272 9496 37324
rect 9548 37272 9554 37324
rect 10134 37272 10140 37324
rect 10192 37272 10198 37324
rect 10318 37272 10324 37324
rect 10376 37272 10382 37324
rect 10410 37272 10416 37324
rect 10468 37312 10474 37324
rect 10505 37315 10563 37321
rect 10505 37312 10517 37315
rect 10468 37284 10517 37312
rect 10468 37272 10474 37284
rect 10505 37281 10517 37284
rect 10551 37281 10563 37315
rect 10505 37275 10563 37281
rect 13541 37315 13599 37321
rect 13541 37281 13553 37315
rect 13587 37312 13599 37315
rect 14550 37312 14556 37324
rect 13587 37284 14556 37312
rect 13587 37281 13599 37284
rect 13541 37275 13599 37281
rect 14550 37272 14556 37284
rect 14608 37272 14614 37324
rect 15105 37315 15163 37321
rect 15105 37281 15117 37315
rect 15151 37312 15163 37315
rect 15194 37312 15200 37324
rect 15151 37284 15200 37312
rect 15151 37281 15163 37284
rect 15105 37275 15163 37281
rect 15194 37272 15200 37284
rect 15252 37272 15258 37324
rect 15749 37315 15807 37321
rect 15749 37281 15761 37315
rect 15795 37312 15807 37315
rect 16390 37312 16396 37324
rect 15795 37284 16396 37312
rect 15795 37281 15807 37284
rect 15749 37275 15807 37281
rect 16390 37272 16396 37284
rect 16448 37272 16454 37324
rect 13817 37247 13875 37253
rect 13817 37213 13829 37247
rect 13863 37244 13875 37247
rect 15286 37244 15292 37256
rect 13863 37216 15292 37244
rect 13863 37213 13875 37216
rect 13817 37207 13875 37213
rect 15286 37204 15292 37216
rect 15344 37204 15350 37256
rect 15473 37247 15531 37253
rect 15473 37213 15485 37247
rect 15519 37244 15531 37247
rect 15654 37244 15660 37256
rect 15519 37216 15660 37244
rect 15519 37213 15531 37216
rect 15473 37207 15531 37213
rect 15654 37204 15660 37216
rect 15712 37204 15718 37256
rect 15102 37136 15108 37188
rect 15160 37176 15166 37188
rect 16500 37176 16528 37352
rect 16942 37272 16948 37324
rect 17000 37272 17006 37324
rect 18248 37321 18276 37352
rect 18874 37340 18880 37392
rect 18932 37380 18938 37392
rect 19153 37383 19211 37389
rect 19153 37380 19165 37383
rect 18932 37352 19165 37380
rect 18932 37340 18938 37352
rect 19153 37349 19165 37352
rect 19199 37349 19211 37383
rect 19153 37343 19211 37349
rect 19720 37352 20760 37380
rect 19720 37321 19748 37352
rect 20732 37324 20760 37352
rect 18233 37315 18291 37321
rect 18233 37281 18245 37315
rect 18279 37312 18291 37315
rect 19613 37315 19671 37321
rect 19613 37312 19625 37315
rect 18279 37284 19625 37312
rect 18279 37281 18291 37284
rect 18233 37275 18291 37281
rect 19613 37281 19625 37284
rect 19659 37281 19671 37315
rect 19613 37275 19671 37281
rect 19705 37315 19763 37321
rect 19705 37281 19717 37315
rect 19751 37281 19763 37315
rect 19705 37275 19763 37281
rect 19981 37315 20039 37321
rect 19981 37281 19993 37315
rect 20027 37281 20039 37315
rect 19981 37275 20039 37281
rect 18325 37247 18383 37253
rect 18325 37213 18337 37247
rect 18371 37244 18383 37247
rect 19334 37244 19340 37256
rect 18371 37216 19340 37244
rect 18371 37213 18383 37216
rect 18325 37207 18383 37213
rect 19334 37204 19340 37216
rect 19392 37204 19398 37256
rect 19996 37244 20024 37275
rect 20162 37272 20168 37324
rect 20220 37272 20226 37324
rect 20714 37272 20720 37324
rect 20772 37272 20778 37324
rect 20809 37315 20867 37321
rect 20809 37281 20821 37315
rect 20855 37281 20867 37315
rect 20809 37275 20867 37281
rect 20438 37244 20444 37256
rect 19996 37216 20444 37244
rect 20438 37204 20444 37216
rect 20496 37204 20502 37256
rect 20530 37204 20536 37256
rect 20588 37244 20594 37256
rect 20824 37244 20852 37275
rect 20898 37272 20904 37324
rect 20956 37272 20962 37324
rect 21082 37272 21088 37324
rect 21140 37272 21146 37324
rect 21266 37272 21272 37324
rect 21324 37272 21330 37324
rect 21540 37321 21568 37420
rect 21634 37408 21640 37460
rect 21692 37448 21698 37460
rect 22649 37451 22707 37457
rect 22649 37448 22661 37451
rect 21692 37420 22661 37448
rect 21692 37408 21698 37420
rect 22649 37417 22661 37420
rect 22695 37417 22707 37451
rect 22649 37411 22707 37417
rect 23382 37408 23388 37460
rect 23440 37408 23446 37460
rect 24504 37420 26832 37448
rect 23474 37340 23480 37392
rect 23532 37380 23538 37392
rect 24504 37389 24532 37420
rect 24259 37383 24317 37389
rect 24259 37380 24271 37383
rect 23532 37352 24271 37380
rect 23532 37340 23538 37352
rect 24259 37349 24271 37352
rect 24305 37349 24317 37383
rect 24259 37343 24317 37349
rect 24489 37383 24547 37389
rect 24489 37349 24501 37383
rect 24535 37349 24547 37383
rect 24489 37343 24547 37349
rect 24946 37340 24952 37392
rect 25004 37380 25010 37392
rect 25593 37383 25651 37389
rect 25593 37380 25605 37383
rect 25004 37352 25605 37380
rect 25004 37340 25010 37352
rect 25593 37349 25605 37352
rect 25639 37380 25651 37383
rect 26804 37380 26832 37420
rect 28994 37408 29000 37460
rect 29052 37448 29058 37460
rect 30377 37451 30435 37457
rect 30377 37448 30389 37451
rect 29052 37420 30389 37448
rect 29052 37408 29058 37420
rect 30377 37417 30389 37420
rect 30423 37448 30435 37451
rect 30466 37448 30472 37460
rect 30423 37420 30472 37448
rect 30423 37417 30435 37420
rect 30377 37411 30435 37417
rect 30466 37408 30472 37420
rect 30524 37408 30530 37460
rect 30558 37408 30564 37460
rect 30616 37448 30622 37460
rect 31294 37448 31300 37460
rect 30616 37420 31300 37448
rect 30616 37408 30622 37420
rect 31294 37408 31300 37420
rect 31352 37408 31358 37460
rect 27338 37380 27344 37392
rect 25639 37352 26188 37380
rect 25639 37349 25651 37352
rect 25593 37343 25651 37349
rect 21525 37315 21583 37321
rect 21525 37281 21537 37315
rect 21571 37281 21583 37315
rect 21525 37275 21583 37281
rect 22370 37272 22376 37324
rect 22428 37312 22434 37324
rect 22741 37315 22799 37321
rect 22741 37312 22753 37315
rect 22428 37284 22753 37312
rect 22428 37272 22434 37284
rect 22741 37281 22753 37284
rect 22787 37281 22799 37315
rect 22741 37275 22799 37281
rect 23566 37272 23572 37324
rect 23624 37272 23630 37324
rect 23658 37272 23664 37324
rect 23716 37312 23722 37324
rect 24397 37315 24455 37321
rect 24397 37312 24409 37315
rect 23716 37284 24409 37312
rect 23716 37272 23722 37284
rect 24397 37281 24409 37284
rect 24443 37281 24455 37315
rect 24397 37275 24455 37281
rect 24578 37272 24584 37324
rect 24636 37272 24642 37324
rect 24857 37315 24915 37321
rect 24857 37281 24869 37315
rect 24903 37312 24915 37315
rect 25130 37312 25136 37324
rect 24903 37284 25136 37312
rect 24903 37281 24915 37284
rect 24857 37275 24915 37281
rect 25130 37272 25136 37284
rect 25188 37272 25194 37324
rect 26160 37321 26188 37352
rect 26804 37352 27344 37380
rect 26804 37321 26832 37352
rect 27338 37340 27344 37352
rect 27396 37380 27402 37392
rect 27617 37383 27675 37389
rect 27617 37380 27629 37383
rect 27396 37352 27629 37380
rect 27396 37340 27402 37352
rect 27617 37349 27629 37352
rect 27663 37349 27675 37383
rect 27617 37343 27675 37349
rect 30101 37383 30159 37389
rect 30101 37349 30113 37383
rect 30147 37380 30159 37383
rect 30576 37380 30604 37408
rect 30147 37352 30604 37380
rect 30745 37383 30803 37389
rect 30147 37349 30159 37352
rect 30101 37343 30159 37349
rect 30745 37349 30757 37383
rect 30791 37349 30803 37383
rect 31680 37380 31708 37624
rect 30745 37343 30803 37349
rect 31036 37352 31708 37380
rect 26145 37315 26203 37321
rect 26145 37281 26157 37315
rect 26191 37281 26203 37315
rect 26145 37275 26203 37281
rect 26789 37315 26847 37321
rect 26789 37281 26801 37315
rect 26835 37281 26847 37315
rect 26789 37275 26847 37281
rect 26878 37272 26884 37324
rect 26936 37272 26942 37324
rect 28994 37321 29000 37324
rect 28972 37315 29000 37321
rect 28972 37281 28984 37315
rect 28972 37275 29000 37281
rect 28994 37272 29000 37275
rect 29052 37272 29058 37324
rect 29086 37272 29092 37324
rect 29144 37272 29150 37324
rect 30190 37272 30196 37324
rect 30248 37312 30254 37324
rect 30285 37315 30343 37321
rect 30285 37312 30297 37315
rect 30248 37284 30297 37312
rect 30248 37272 30254 37284
rect 30285 37281 30297 37284
rect 30331 37281 30343 37315
rect 30285 37275 30343 37281
rect 30469 37315 30527 37321
rect 30469 37281 30481 37315
rect 30515 37281 30527 37315
rect 30760 37312 30788 37343
rect 31036 37321 31064 37352
rect 31021 37315 31079 37321
rect 30760 37284 30972 37312
rect 30469 37275 30527 37281
rect 20588 37216 20852 37244
rect 20588 37204 20594 37216
rect 22922 37204 22928 37256
rect 22980 37244 22986 37256
rect 23753 37247 23811 37253
rect 23753 37244 23765 37247
rect 22980 37216 23765 37244
rect 22980 37204 22986 37216
rect 23753 37213 23765 37216
rect 23799 37213 23811 37247
rect 23753 37207 23811 37213
rect 24121 37247 24179 37253
rect 24121 37213 24133 37247
rect 24167 37213 24179 37247
rect 24121 37207 24179 37213
rect 26421 37247 26479 37253
rect 26421 37213 26433 37247
rect 26467 37244 26479 37247
rect 26694 37244 26700 37256
rect 26467 37216 26700 37244
rect 26467 37213 26479 37216
rect 26421 37207 26479 37213
rect 18966 37176 18972 37188
rect 15160 37148 16528 37176
rect 18432 37148 18972 37176
rect 15160 37136 15166 37148
rect 9306 37068 9312 37120
rect 9364 37108 9370 37120
rect 9585 37111 9643 37117
rect 9585 37108 9597 37111
rect 9364 37080 9597 37108
rect 9364 37068 9370 37080
rect 9585 37077 9597 37080
rect 9631 37077 9643 37111
rect 9585 37071 9643 37077
rect 10686 37068 10692 37120
rect 10744 37068 10750 37120
rect 13722 37068 13728 37120
rect 13780 37068 13786 37120
rect 15562 37068 15568 37120
rect 15620 37108 15626 37120
rect 18322 37108 18328 37120
rect 15620 37080 18328 37108
rect 15620 37068 15626 37080
rect 18322 37068 18328 37080
rect 18380 37068 18386 37120
rect 18432 37117 18460 37148
rect 18966 37136 18972 37148
rect 19024 37176 19030 37188
rect 19153 37179 19211 37185
rect 19153 37176 19165 37179
rect 19024 37148 19165 37176
rect 19024 37136 19030 37148
rect 19153 37145 19165 37148
rect 19199 37176 19211 37179
rect 20622 37176 20628 37188
rect 19199 37148 20628 37176
rect 19199 37145 19211 37148
rect 19153 37139 19211 37145
rect 20622 37136 20628 37148
rect 20680 37136 20686 37188
rect 23290 37136 23296 37188
rect 23348 37176 23354 37188
rect 24136 37176 24164 37207
rect 26694 37204 26700 37216
rect 26752 37204 26758 37256
rect 28258 37204 28264 37256
rect 28316 37244 28322 37256
rect 28810 37244 28816 37256
rect 28316 37216 28816 37244
rect 28316 37204 28322 37216
rect 28810 37204 28816 37216
rect 28868 37204 28874 37256
rect 29825 37247 29883 37253
rect 29825 37213 29837 37247
rect 29871 37213 29883 37247
rect 29825 37207 29883 37213
rect 30009 37247 30067 37253
rect 30009 37213 30021 37247
rect 30055 37244 30067 37247
rect 30484 37244 30512 37275
rect 30055 37216 30512 37244
rect 30055 37213 30067 37216
rect 30009 37207 30067 37213
rect 23348 37148 24164 37176
rect 23348 37136 23354 37148
rect 26878 37136 26884 37188
rect 26936 37176 26942 37188
rect 27157 37179 27215 37185
rect 27157 37176 27169 37179
rect 26936 37148 27169 37176
rect 26936 37136 26942 37148
rect 27157 37145 27169 37148
rect 27203 37145 27215 37179
rect 27157 37139 27215 37145
rect 27341 37179 27399 37185
rect 27341 37145 27353 37179
rect 27387 37176 27399 37179
rect 27430 37176 27436 37188
rect 27387 37148 27436 37176
rect 27387 37145 27399 37148
rect 27341 37139 27399 37145
rect 27430 37136 27436 37148
rect 27488 37136 27494 37188
rect 29365 37179 29423 37185
rect 29365 37145 29377 37179
rect 29411 37145 29423 37179
rect 29365 37139 29423 37145
rect 18417 37111 18475 37117
rect 18417 37077 18429 37111
rect 18463 37077 18475 37111
rect 18417 37071 18475 37077
rect 18598 37068 18604 37120
rect 18656 37068 18662 37120
rect 19889 37111 19947 37117
rect 19889 37077 19901 37111
rect 19935 37108 19947 37111
rect 23474 37108 23480 37120
rect 19935 37080 23480 37108
rect 19935 37077 19947 37080
rect 19889 37071 19947 37077
rect 23474 37068 23480 37080
rect 23532 37068 23538 37120
rect 24765 37111 24823 37117
rect 24765 37077 24777 37111
rect 24811 37108 24823 37111
rect 24946 37108 24952 37120
rect 24811 37080 24952 37108
rect 24811 37077 24823 37080
rect 24765 37071 24823 37077
rect 24946 37068 24952 37080
rect 25004 37068 25010 37120
rect 25866 37068 25872 37120
rect 25924 37108 25930 37120
rect 26053 37111 26111 37117
rect 26053 37108 26065 37111
rect 25924 37080 26065 37108
rect 25924 37068 25930 37080
rect 26053 37077 26065 37080
rect 26099 37077 26111 37111
rect 26053 37071 26111 37077
rect 26786 37068 26792 37120
rect 26844 37108 26850 37120
rect 27065 37111 27123 37117
rect 27065 37108 27077 37111
rect 26844 37080 27077 37108
rect 26844 37068 26850 37080
rect 27065 37077 27077 37080
rect 27111 37077 27123 37111
rect 27065 37071 27123 37077
rect 27798 37068 27804 37120
rect 27856 37108 27862 37120
rect 28169 37111 28227 37117
rect 28169 37108 28181 37111
rect 27856 37080 28181 37108
rect 27856 37068 27862 37080
rect 28169 37077 28181 37080
rect 28215 37077 28227 37111
rect 28169 37071 28227 37077
rect 28718 37068 28724 37120
rect 28776 37108 28782 37120
rect 29380 37108 29408 37139
rect 28776 37080 29408 37108
rect 28776 37068 28782 37080
rect 29454 37068 29460 37120
rect 29512 37108 29518 37120
rect 29840 37108 29868 37207
rect 30300 37188 30328 37216
rect 30742 37204 30748 37256
rect 30800 37204 30806 37256
rect 30944 37244 30972 37284
rect 31021 37281 31033 37315
rect 31067 37281 31079 37315
rect 31021 37275 31079 37281
rect 31113 37315 31171 37321
rect 31113 37281 31125 37315
rect 31159 37281 31171 37315
rect 31113 37275 31171 37281
rect 31128 37244 31156 37275
rect 31294 37272 31300 37324
rect 31352 37272 31358 37324
rect 30944 37216 31156 37244
rect 30282 37136 30288 37188
rect 30340 37136 30346 37188
rect 30653 37179 30711 37185
rect 30653 37176 30665 37179
rect 30392 37148 30665 37176
rect 30392 37108 30420 37148
rect 30653 37145 30665 37148
rect 30699 37176 30711 37179
rect 31018 37176 31024 37188
rect 30699 37148 31024 37176
rect 30699 37145 30711 37148
rect 30653 37139 30711 37145
rect 31018 37136 31024 37148
rect 31076 37136 31082 37188
rect 31110 37136 31116 37188
rect 31168 37136 31174 37188
rect 29512 37080 30420 37108
rect 29512 37068 29518 37080
rect 30558 37068 30564 37120
rect 30616 37108 30622 37120
rect 30929 37111 30987 37117
rect 30929 37108 30941 37111
rect 30616 37080 30941 37108
rect 30616 37068 30622 37080
rect 30929 37077 30941 37080
rect 30975 37077 30987 37111
rect 30929 37071 30987 37077
rect 552 37018 31648 37040
rect 552 36966 3662 37018
rect 3714 36966 3726 37018
rect 3778 36966 3790 37018
rect 3842 36966 3854 37018
rect 3906 36966 3918 37018
rect 3970 36966 11436 37018
rect 11488 36966 11500 37018
rect 11552 36966 11564 37018
rect 11616 36966 11628 37018
rect 11680 36966 11692 37018
rect 11744 36966 19210 37018
rect 19262 36966 19274 37018
rect 19326 36966 19338 37018
rect 19390 36966 19402 37018
rect 19454 36966 19466 37018
rect 19518 36966 26984 37018
rect 27036 36966 27048 37018
rect 27100 36966 27112 37018
rect 27164 36966 27176 37018
rect 27228 36966 27240 37018
rect 27292 36966 31648 37018
rect 552 36944 31648 36966
rect 9769 36907 9827 36913
rect 9769 36873 9781 36907
rect 9815 36904 9827 36907
rect 10134 36904 10140 36916
rect 9815 36876 10140 36904
rect 9815 36873 9827 36876
rect 9769 36867 9827 36873
rect 10134 36864 10140 36876
rect 10192 36864 10198 36916
rect 12894 36904 12900 36916
rect 12406 36876 12900 36904
rect 8294 36768 8300 36780
rect 8036 36740 8300 36768
rect 8036 36709 8064 36740
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 10321 36771 10379 36777
rect 10321 36737 10333 36771
rect 10367 36768 10379 36771
rect 12406 36768 12434 36876
rect 12894 36864 12900 36876
rect 12952 36904 12958 36916
rect 13262 36904 13268 36916
rect 12952 36876 13268 36904
rect 12952 36864 12958 36876
rect 13262 36864 13268 36876
rect 13320 36864 13326 36916
rect 14550 36864 14556 36916
rect 14608 36904 14614 36916
rect 15102 36904 15108 36916
rect 14608 36876 15108 36904
rect 14608 36864 14614 36876
rect 15102 36864 15108 36876
rect 15160 36864 15166 36916
rect 16206 36864 16212 36916
rect 16264 36864 16270 36916
rect 17862 36864 17868 36916
rect 17920 36864 17926 36916
rect 18966 36864 18972 36916
rect 19024 36864 19030 36916
rect 20714 36864 20720 36916
rect 20772 36904 20778 36916
rect 20772 36876 20852 36904
rect 20772 36864 20778 36876
rect 13081 36839 13139 36845
rect 13081 36805 13093 36839
rect 13127 36805 13139 36839
rect 13081 36799 13139 36805
rect 10367 36740 12434 36768
rect 13096 36768 13124 36799
rect 13814 36796 13820 36848
rect 13872 36796 13878 36848
rect 15654 36836 15660 36848
rect 14476 36808 15660 36836
rect 13725 36771 13783 36777
rect 13725 36768 13737 36771
rect 13096 36740 13737 36768
rect 10367 36737 10379 36740
rect 10321 36731 10379 36737
rect 13725 36737 13737 36740
rect 13771 36768 13783 36771
rect 14476 36768 14504 36808
rect 15654 36796 15660 36808
rect 15712 36796 15718 36848
rect 16114 36796 16120 36848
rect 16172 36836 16178 36848
rect 20824 36836 20852 36876
rect 20898 36864 20904 36916
rect 20956 36904 20962 36916
rect 20993 36907 21051 36913
rect 20993 36904 21005 36907
rect 20956 36876 21005 36904
rect 20956 36864 20962 36876
rect 20993 36873 21005 36876
rect 21039 36873 21051 36907
rect 20993 36867 21051 36873
rect 21082 36864 21088 36916
rect 21140 36904 21146 36916
rect 22922 36904 22928 36916
rect 21140 36876 22928 36904
rect 21140 36864 21146 36876
rect 22922 36864 22928 36876
rect 22980 36864 22986 36916
rect 23566 36864 23572 36916
rect 23624 36904 23630 36916
rect 23661 36907 23719 36913
rect 23661 36904 23673 36907
rect 23624 36876 23673 36904
rect 23624 36864 23630 36876
rect 23661 36873 23673 36876
rect 23707 36873 23719 36907
rect 23661 36867 23719 36873
rect 27249 36907 27307 36913
rect 27249 36873 27261 36907
rect 27295 36904 27307 36907
rect 27338 36904 27344 36916
rect 27295 36876 27344 36904
rect 27295 36873 27307 36876
rect 27249 36867 27307 36873
rect 27338 36864 27344 36876
rect 27396 36864 27402 36916
rect 29641 36907 29699 36913
rect 29641 36873 29653 36907
rect 29687 36904 29699 36907
rect 30282 36904 30288 36916
rect 29687 36876 30288 36904
rect 29687 36873 29699 36876
rect 29641 36867 29699 36873
rect 30282 36864 30288 36876
rect 30340 36864 30346 36916
rect 21913 36839 21971 36845
rect 21913 36836 21925 36839
rect 16172 36808 16436 36836
rect 16172 36796 16178 36808
rect 16408 36780 16436 36808
rect 20824 36808 21925 36836
rect 13771 36740 14504 36768
rect 13771 36737 13783 36740
rect 13725 36731 13783 36737
rect 14550 36728 14556 36780
rect 14608 36728 14614 36780
rect 15562 36768 15568 36780
rect 14660 36740 15568 36768
rect 8021 36703 8079 36709
rect 8021 36669 8033 36703
rect 8067 36669 8079 36703
rect 8021 36663 8079 36669
rect 8113 36703 8171 36709
rect 8113 36669 8125 36703
rect 8159 36700 8171 36703
rect 8389 36703 8447 36709
rect 8389 36700 8401 36703
rect 8159 36672 8401 36700
rect 8159 36669 8171 36672
rect 8113 36663 8171 36669
rect 8389 36669 8401 36672
rect 8435 36669 8447 36703
rect 8389 36663 8447 36669
rect 9582 36660 9588 36712
rect 9640 36700 9646 36712
rect 10505 36703 10563 36709
rect 10505 36700 10517 36703
rect 9640 36672 10517 36700
rect 9640 36660 9646 36672
rect 10505 36669 10517 36672
rect 10551 36669 10563 36703
rect 11149 36703 11207 36709
rect 11149 36700 11161 36703
rect 10505 36663 10563 36669
rect 10888 36672 11161 36700
rect 8656 36635 8714 36641
rect 8656 36601 8668 36635
rect 8702 36632 8714 36635
rect 9030 36632 9036 36644
rect 8702 36604 9036 36632
rect 8702 36601 8714 36604
rect 8656 36595 8714 36601
rect 9030 36592 9036 36604
rect 9088 36592 9094 36644
rect 10410 36592 10416 36644
rect 10468 36592 10474 36644
rect 10888 36573 10916 36672
rect 11149 36669 11161 36672
rect 11195 36669 11207 36703
rect 11149 36663 11207 36669
rect 11238 36660 11244 36712
rect 11296 36660 11302 36712
rect 11422 36660 11428 36712
rect 11480 36660 11486 36712
rect 11517 36703 11575 36709
rect 11517 36669 11529 36703
rect 11563 36700 11575 36703
rect 12618 36700 12624 36712
rect 11563 36672 12624 36700
rect 11563 36669 11575 36672
rect 11517 36663 11575 36669
rect 11054 36592 11060 36644
rect 11112 36632 11118 36644
rect 11532 36632 11560 36663
rect 12618 36660 12624 36672
rect 12676 36660 12682 36712
rect 14001 36703 14059 36709
rect 14001 36669 14013 36703
rect 14047 36700 14059 36703
rect 14660 36700 14688 36740
rect 15120 36709 15148 36740
rect 15562 36728 15568 36740
rect 15620 36728 15626 36780
rect 15948 36740 16252 36768
rect 14047 36672 14688 36700
rect 14737 36703 14795 36709
rect 14047 36669 14059 36672
rect 14001 36663 14059 36669
rect 14737 36669 14749 36703
rect 14783 36700 14795 36703
rect 15013 36703 15071 36709
rect 14783 36672 14964 36700
rect 14783 36669 14795 36672
rect 14737 36663 14795 36669
rect 11112 36604 11560 36632
rect 13357 36635 13415 36641
rect 11112 36592 11118 36604
rect 13357 36601 13369 36635
rect 13403 36632 13415 36635
rect 14016 36632 14044 36663
rect 13403 36604 14044 36632
rect 13403 36601 13415 36604
rect 13357 36595 13415 36601
rect 14182 36592 14188 36644
rect 14240 36632 14246 36644
rect 14369 36635 14427 36641
rect 14369 36632 14381 36635
rect 14240 36604 14381 36632
rect 14240 36592 14246 36604
rect 14369 36601 14381 36604
rect 14415 36601 14427 36635
rect 14369 36595 14427 36601
rect 10873 36567 10931 36573
rect 10873 36533 10885 36567
rect 10919 36533 10931 36567
rect 10873 36527 10931 36533
rect 10962 36524 10968 36576
rect 11020 36524 11026 36576
rect 12897 36567 12955 36573
rect 12897 36533 12909 36567
rect 12943 36564 12955 36567
rect 12986 36564 12992 36576
rect 12943 36536 12992 36564
rect 12943 36533 12955 36536
rect 12897 36527 12955 36533
rect 12986 36524 12992 36536
rect 13044 36524 13050 36576
rect 14550 36524 14556 36576
rect 14608 36564 14614 36576
rect 14936 36564 14964 36672
rect 15013 36669 15025 36703
rect 15059 36669 15071 36703
rect 15013 36663 15071 36669
rect 15105 36703 15163 36709
rect 15105 36669 15117 36703
rect 15151 36669 15163 36703
rect 15105 36663 15163 36669
rect 15289 36703 15347 36709
rect 15289 36669 15301 36703
rect 15335 36700 15347 36703
rect 15654 36700 15660 36712
rect 15335 36672 15660 36700
rect 15335 36669 15347 36672
rect 15289 36663 15347 36669
rect 15028 36632 15056 36663
rect 15654 36660 15660 36672
rect 15712 36700 15718 36712
rect 15948 36700 15976 36740
rect 15712 36672 15976 36700
rect 15712 36660 15718 36672
rect 16022 36660 16028 36712
rect 16080 36700 16086 36712
rect 16117 36703 16175 36709
rect 16117 36700 16129 36703
rect 16080 36672 16129 36700
rect 16080 36660 16086 36672
rect 16117 36669 16129 36672
rect 16163 36669 16175 36703
rect 16224 36700 16252 36740
rect 16390 36728 16396 36780
rect 16448 36728 16454 36780
rect 18029 36771 18087 36777
rect 18029 36737 18041 36771
rect 18075 36768 18087 36771
rect 18690 36768 18696 36780
rect 18075 36740 18696 36768
rect 18075 36737 18087 36740
rect 18029 36731 18087 36737
rect 18690 36728 18696 36740
rect 18748 36728 18754 36780
rect 19058 36768 19064 36780
rect 18800 36740 19064 36768
rect 16224 36672 16436 36700
rect 16117 36663 16175 36669
rect 16206 36632 16212 36644
rect 15028 36604 16212 36632
rect 16206 36592 16212 36604
rect 16264 36592 16270 36644
rect 16408 36632 16436 36672
rect 16482 36660 16488 36712
rect 16540 36660 16546 36712
rect 18141 36703 18199 36709
rect 18141 36669 18153 36703
rect 18187 36700 18199 36703
rect 18800 36700 18828 36740
rect 19058 36728 19064 36740
rect 19116 36728 19122 36780
rect 20824 36768 20852 36808
rect 21913 36805 21925 36808
rect 21959 36805 21971 36839
rect 27356 36836 27384 36864
rect 27356 36808 27936 36836
rect 21913 36799 21971 36805
rect 19168 36740 20852 36768
rect 18187 36672 18828 36700
rect 18877 36703 18935 36709
rect 18187 36669 18199 36672
rect 18141 36663 18199 36669
rect 18877 36669 18889 36703
rect 18923 36700 18935 36703
rect 19168 36700 19196 36740
rect 22830 36728 22836 36780
rect 22888 36768 22894 36780
rect 22888 36740 23336 36768
rect 22888 36728 22894 36740
rect 18923 36672 19196 36700
rect 18923 36669 18935 36672
rect 18877 36663 18935 36669
rect 17954 36632 17960 36644
rect 16408 36604 17960 36632
rect 17954 36592 17960 36604
rect 18012 36592 18018 36644
rect 18417 36635 18475 36641
rect 18417 36601 18429 36635
rect 18463 36601 18475 36635
rect 18417 36595 18475 36601
rect 18509 36635 18567 36641
rect 18509 36601 18521 36635
rect 18555 36601 18567 36635
rect 18509 36595 18567 36601
rect 15562 36564 15568 36576
rect 14608 36536 15568 36564
rect 14608 36524 14614 36536
rect 15562 36524 15568 36536
rect 15620 36564 15626 36576
rect 16114 36564 16120 36576
rect 15620 36536 16120 36564
rect 15620 36524 15626 36536
rect 16114 36524 16120 36536
rect 16172 36524 16178 36576
rect 18138 36524 18144 36576
rect 18196 36564 18202 36576
rect 18432 36564 18460 36595
rect 18196 36536 18460 36564
rect 18524 36564 18552 36595
rect 18782 36592 18788 36644
rect 18840 36632 18846 36644
rect 18892 36632 18920 36663
rect 19242 36660 19248 36712
rect 19300 36660 19306 36712
rect 19337 36703 19395 36709
rect 19337 36669 19349 36703
rect 19383 36669 19395 36703
rect 21085 36703 21143 36709
rect 21085 36700 21097 36703
rect 19337 36663 19395 36669
rect 20548 36672 21097 36700
rect 18840 36604 18920 36632
rect 18840 36592 18846 36604
rect 18966 36592 18972 36644
rect 19024 36632 19030 36644
rect 19352 36632 19380 36663
rect 20548 36644 20576 36672
rect 21085 36669 21097 36672
rect 21131 36669 21143 36703
rect 21085 36663 21143 36669
rect 21450 36660 21456 36712
rect 21508 36700 21514 36712
rect 21729 36703 21787 36709
rect 21729 36700 21741 36703
rect 21508 36672 21741 36700
rect 21508 36660 21514 36672
rect 21729 36669 21741 36672
rect 21775 36669 21787 36703
rect 21729 36663 21787 36669
rect 21910 36660 21916 36712
rect 21968 36700 21974 36712
rect 22097 36703 22155 36709
rect 22097 36700 22109 36703
rect 21968 36672 22109 36700
rect 21968 36660 21974 36672
rect 22097 36669 22109 36672
rect 22143 36669 22155 36703
rect 22097 36663 22155 36669
rect 23014 36660 23020 36712
rect 23072 36660 23078 36712
rect 23308 36709 23336 36740
rect 23934 36728 23940 36780
rect 23992 36768 23998 36780
rect 23992 36740 24532 36768
rect 23992 36728 23998 36740
rect 23293 36703 23351 36709
rect 23293 36669 23305 36703
rect 23339 36669 23351 36703
rect 23293 36663 23351 36669
rect 23477 36703 23535 36709
rect 23477 36669 23489 36703
rect 23523 36700 23535 36703
rect 23658 36700 23664 36712
rect 23523 36672 23664 36700
rect 23523 36669 23535 36672
rect 23477 36663 23535 36669
rect 23658 36660 23664 36672
rect 23716 36660 23722 36712
rect 24118 36660 24124 36712
rect 24176 36660 24182 36712
rect 24394 36660 24400 36712
rect 24452 36660 24458 36712
rect 24504 36700 24532 36740
rect 25866 36728 25872 36780
rect 25924 36728 25930 36780
rect 27798 36728 27804 36780
rect 27856 36728 27862 36780
rect 27908 36777 27936 36808
rect 27893 36771 27951 36777
rect 27893 36737 27905 36771
rect 27939 36737 27951 36771
rect 27893 36731 27951 36737
rect 24504 36672 24808 36700
rect 24780 36644 24808 36672
rect 29178 36660 29184 36712
rect 29236 36660 29242 36712
rect 29273 36703 29331 36709
rect 29273 36669 29285 36703
rect 29319 36700 29331 36703
rect 29917 36703 29975 36709
rect 29917 36700 29929 36703
rect 29319 36672 29929 36700
rect 29319 36669 29331 36672
rect 29273 36663 29331 36669
rect 29917 36669 29929 36672
rect 29963 36669 29975 36703
rect 29917 36663 29975 36669
rect 19024 36604 19380 36632
rect 19024 36592 19030 36604
rect 20346 36592 20352 36644
rect 20404 36592 20410 36644
rect 20530 36592 20536 36644
rect 20588 36592 20594 36644
rect 20622 36592 20628 36644
rect 20680 36592 20686 36644
rect 20806 36592 20812 36644
rect 20864 36632 20870 36644
rect 23175 36635 23233 36641
rect 20864 36604 21588 36632
rect 20864 36592 20870 36604
rect 18693 36567 18751 36573
rect 18693 36564 18705 36567
rect 18524 36536 18705 36564
rect 18196 36524 18202 36536
rect 18693 36533 18705 36536
rect 18739 36533 18751 36567
rect 18693 36527 18751 36533
rect 20254 36524 20260 36576
rect 20312 36564 20318 36576
rect 21560 36573 21588 36604
rect 23175 36601 23187 36635
rect 23221 36632 23233 36635
rect 23385 36635 23443 36641
rect 23221 36601 23244 36632
rect 23175 36595 23244 36601
rect 23385 36601 23397 36635
rect 23431 36632 23443 36635
rect 24026 36632 24032 36644
rect 23431 36604 24032 36632
rect 23431 36601 23443 36604
rect 23385 36595 23443 36601
rect 21269 36567 21327 36573
rect 21269 36564 21281 36567
rect 20312 36536 21281 36564
rect 20312 36524 20318 36536
rect 21269 36533 21281 36536
rect 21315 36533 21327 36567
rect 21269 36527 21327 36533
rect 21545 36567 21603 36573
rect 21545 36533 21557 36567
rect 21591 36533 21603 36567
rect 23216 36564 23244 36595
rect 24026 36592 24032 36604
rect 24084 36592 24090 36644
rect 24305 36635 24363 36641
rect 24305 36601 24317 36635
rect 24351 36632 24363 36635
rect 24642 36635 24700 36641
rect 24642 36632 24654 36635
rect 24351 36604 24654 36632
rect 24351 36601 24363 36604
rect 24305 36595 24363 36601
rect 24642 36601 24654 36604
rect 24688 36601 24700 36635
rect 24642 36595 24700 36601
rect 24762 36592 24768 36644
rect 24820 36592 24826 36644
rect 25222 36592 25228 36644
rect 25280 36632 25286 36644
rect 26114 36635 26172 36641
rect 26114 36632 26126 36635
rect 25280 36604 26126 36632
rect 25280 36592 25286 36604
rect 26114 36601 26126 36604
rect 26160 36601 26172 36635
rect 26114 36595 26172 36601
rect 26602 36592 26608 36644
rect 26660 36632 26666 36644
rect 26660 36604 27384 36632
rect 26660 36592 26666 36604
rect 23474 36564 23480 36576
rect 23216 36536 23480 36564
rect 21545 36527 21603 36533
rect 23474 36524 23480 36536
rect 23532 36524 23538 36576
rect 25774 36524 25780 36576
rect 25832 36524 25838 36576
rect 27356 36573 27384 36604
rect 29454 36592 29460 36644
rect 29512 36592 29518 36644
rect 30006 36592 30012 36644
rect 30064 36632 30070 36644
rect 30162 36635 30220 36641
rect 30162 36632 30174 36635
rect 30064 36604 30174 36632
rect 30064 36592 30070 36604
rect 30162 36601 30174 36604
rect 30208 36601 30220 36635
rect 30162 36595 30220 36601
rect 27341 36567 27399 36573
rect 27341 36533 27353 36567
rect 27387 36533 27399 36567
rect 27341 36527 27399 36533
rect 27709 36567 27767 36573
rect 27709 36533 27721 36567
rect 27755 36564 27767 36567
rect 28074 36564 28080 36576
rect 27755 36536 28080 36564
rect 27755 36533 27767 36536
rect 27709 36527 27767 36533
rect 28074 36524 28080 36536
rect 28132 36524 28138 36576
rect 29638 36524 29644 36576
rect 29696 36573 29702 36576
rect 29696 36567 29715 36573
rect 29703 36533 29715 36567
rect 29696 36527 29715 36533
rect 29825 36567 29883 36573
rect 29825 36533 29837 36567
rect 29871 36564 29883 36567
rect 30558 36564 30564 36576
rect 29871 36536 30564 36564
rect 29871 36533 29883 36536
rect 29825 36527 29883 36533
rect 29696 36524 29702 36527
rect 30558 36524 30564 36536
rect 30616 36524 30622 36576
rect 31297 36567 31355 36573
rect 31297 36533 31309 36567
rect 31343 36564 31355 36567
rect 31343 36536 31708 36564
rect 31343 36533 31355 36536
rect 31297 36527 31355 36533
rect 552 36474 31648 36496
rect 552 36422 4322 36474
rect 4374 36422 4386 36474
rect 4438 36422 4450 36474
rect 4502 36422 4514 36474
rect 4566 36422 4578 36474
rect 4630 36422 12096 36474
rect 12148 36422 12160 36474
rect 12212 36422 12224 36474
rect 12276 36422 12288 36474
rect 12340 36422 12352 36474
rect 12404 36422 19870 36474
rect 19922 36422 19934 36474
rect 19986 36422 19998 36474
rect 20050 36422 20062 36474
rect 20114 36422 20126 36474
rect 20178 36422 27644 36474
rect 27696 36422 27708 36474
rect 27760 36422 27772 36474
rect 27824 36422 27836 36474
rect 27888 36422 27900 36474
rect 27952 36422 31648 36474
rect 552 36400 31648 36422
rect 9030 36320 9036 36372
rect 9088 36320 9094 36372
rect 9858 36360 9864 36372
rect 9416 36332 9864 36360
rect 9306 36184 9312 36236
rect 9364 36184 9370 36236
rect 9416 36233 9444 36332
rect 9858 36320 9864 36332
rect 9916 36320 9922 36372
rect 10045 36363 10103 36369
rect 10045 36329 10057 36363
rect 10091 36360 10103 36363
rect 11422 36360 11428 36372
rect 10091 36332 11428 36360
rect 10091 36329 10103 36332
rect 10045 36323 10103 36329
rect 11422 36320 11428 36332
rect 11480 36320 11486 36372
rect 13170 36320 13176 36372
rect 13228 36320 13234 36372
rect 14550 36320 14556 36372
rect 14608 36320 14614 36372
rect 16022 36320 16028 36372
rect 16080 36360 16086 36372
rect 16209 36363 16267 36369
rect 16209 36360 16221 36363
rect 16080 36332 16221 36360
rect 16080 36320 16086 36332
rect 16209 36329 16221 36332
rect 16255 36329 16267 36363
rect 16209 36323 16267 36329
rect 17954 36320 17960 36372
rect 18012 36360 18018 36372
rect 18966 36360 18972 36372
rect 18012 36332 18972 36360
rect 18012 36320 18018 36332
rect 18966 36320 18972 36332
rect 19024 36320 19030 36372
rect 20438 36360 20444 36372
rect 19536 36332 20444 36360
rect 10962 36292 10968 36304
rect 9508 36264 10968 36292
rect 9508 36233 9536 36264
rect 10962 36252 10968 36264
rect 11020 36252 11026 36304
rect 11238 36252 11244 36304
rect 11296 36292 11302 36304
rect 14568 36292 14596 36320
rect 16761 36295 16819 36301
rect 16761 36292 16773 36295
rect 11296 36264 12112 36292
rect 11296 36252 11302 36264
rect 9401 36227 9459 36233
rect 9401 36193 9413 36227
rect 9447 36193 9459 36227
rect 9401 36187 9459 36193
rect 9493 36227 9551 36233
rect 9493 36193 9505 36227
rect 9539 36193 9551 36227
rect 9493 36187 9551 36193
rect 9677 36227 9735 36233
rect 9677 36193 9689 36227
rect 9723 36224 9735 36227
rect 10226 36224 10232 36236
rect 9723 36196 10232 36224
rect 9723 36193 9735 36196
rect 9677 36187 9735 36193
rect 10226 36184 10232 36196
rect 10284 36184 10290 36236
rect 10321 36227 10379 36233
rect 10321 36193 10333 36227
rect 10367 36193 10379 36227
rect 10321 36187 10379 36193
rect 10413 36227 10471 36233
rect 10413 36193 10425 36227
rect 10459 36193 10471 36227
rect 10413 36187 10471 36193
rect 9582 36116 9588 36168
rect 9640 36156 9646 36168
rect 10336 36156 10364 36187
rect 9640 36128 10364 36156
rect 9640 36116 9646 36128
rect 10428 36088 10456 36187
rect 10502 36184 10508 36236
rect 10560 36184 10566 36236
rect 10686 36184 10692 36236
rect 10744 36184 10750 36236
rect 11974 36184 11980 36236
rect 12032 36184 12038 36236
rect 12084 36233 12112 36264
rect 13924 36264 14596 36292
rect 16316 36264 16773 36292
rect 12069 36227 12127 36233
rect 12069 36193 12081 36227
rect 12115 36224 12127 36227
rect 12158 36224 12164 36236
rect 12115 36196 12164 36224
rect 12115 36193 12127 36196
rect 12069 36187 12127 36193
rect 12158 36184 12164 36196
rect 12216 36184 12222 36236
rect 12253 36227 12311 36233
rect 12253 36193 12265 36227
rect 12299 36193 12311 36227
rect 12253 36187 12311 36193
rect 12345 36227 12403 36233
rect 12345 36193 12357 36227
rect 12391 36224 12403 36227
rect 12618 36224 12624 36236
rect 12391 36196 12624 36224
rect 12391 36193 12403 36196
rect 12345 36187 12403 36193
rect 11238 36116 11244 36168
rect 11296 36156 11302 36168
rect 11514 36156 11520 36168
rect 11296 36128 11520 36156
rect 11296 36116 11302 36128
rect 11514 36116 11520 36128
rect 11572 36116 11578 36168
rect 11882 36116 11888 36168
rect 11940 36116 11946 36168
rect 12268 36156 12296 36187
rect 12618 36184 12624 36196
rect 12676 36224 12682 36236
rect 12802 36224 12808 36236
rect 12676 36196 12808 36224
rect 12676 36184 12682 36196
rect 12802 36184 12808 36196
rect 12860 36184 12866 36236
rect 12894 36184 12900 36236
rect 12952 36184 12958 36236
rect 13357 36227 13415 36233
rect 13357 36193 13369 36227
rect 13403 36224 13415 36227
rect 13814 36224 13820 36236
rect 13403 36196 13820 36224
rect 13403 36193 13415 36196
rect 13357 36187 13415 36193
rect 12710 36156 12716 36168
rect 12268 36128 12716 36156
rect 12710 36116 12716 36128
rect 12768 36116 12774 36168
rect 11900 36088 11928 36116
rect 13372 36088 13400 36187
rect 13814 36184 13820 36196
rect 13872 36184 13878 36236
rect 13924 36233 13952 36264
rect 13909 36227 13967 36233
rect 13909 36193 13921 36227
rect 13955 36193 13967 36227
rect 14369 36227 14427 36233
rect 14369 36224 14381 36227
rect 13909 36187 13967 36193
rect 14016 36196 14381 36224
rect 13541 36159 13599 36165
rect 13541 36125 13553 36159
rect 13587 36156 13599 36159
rect 14016 36156 14044 36196
rect 14369 36193 14381 36196
rect 14415 36193 14427 36227
rect 14369 36187 14427 36193
rect 14645 36227 14703 36233
rect 14645 36193 14657 36227
rect 14691 36224 14703 36227
rect 15470 36224 15476 36236
rect 14691 36196 15476 36224
rect 14691 36193 14703 36196
rect 14645 36187 14703 36193
rect 13587 36128 14044 36156
rect 14093 36159 14151 36165
rect 13587 36125 13599 36128
rect 13541 36119 13599 36125
rect 14093 36125 14105 36159
rect 14139 36156 14151 36159
rect 14274 36156 14280 36168
rect 14139 36128 14280 36156
rect 14139 36125 14151 36128
rect 14093 36119 14151 36125
rect 14274 36116 14280 36128
rect 14332 36116 14338 36168
rect 14384 36156 14412 36187
rect 15470 36184 15476 36196
rect 15528 36184 15534 36236
rect 16117 36227 16175 36233
rect 16117 36193 16129 36227
rect 16163 36224 16175 36227
rect 16206 36224 16212 36236
rect 16163 36196 16212 36224
rect 16163 36193 16175 36196
rect 16117 36187 16175 36193
rect 16206 36184 16212 36196
rect 16264 36184 16270 36236
rect 16316 36233 16344 36264
rect 16761 36261 16773 36264
rect 16807 36292 16819 36295
rect 18874 36292 18880 36304
rect 16807 36264 18880 36292
rect 16807 36261 16819 36264
rect 16761 36255 16819 36261
rect 18874 36252 18880 36264
rect 18932 36252 18938 36304
rect 19536 36301 19564 36332
rect 20438 36320 20444 36332
rect 20496 36360 20502 36372
rect 20622 36360 20628 36372
rect 20496 36332 20628 36360
rect 20496 36320 20502 36332
rect 20622 36320 20628 36332
rect 20680 36320 20686 36372
rect 23474 36320 23480 36372
rect 23532 36320 23538 36372
rect 23750 36320 23756 36372
rect 23808 36360 23814 36372
rect 23845 36363 23903 36369
rect 23845 36360 23857 36363
rect 23808 36332 23857 36360
rect 23808 36320 23814 36332
rect 23845 36329 23857 36332
rect 23891 36329 23903 36363
rect 23845 36323 23903 36329
rect 24118 36320 24124 36372
rect 24176 36320 24182 36372
rect 24394 36320 24400 36372
rect 24452 36360 24458 36372
rect 25317 36363 25375 36369
rect 25317 36360 25329 36363
rect 24452 36332 25329 36360
rect 24452 36320 24458 36332
rect 25317 36329 25329 36332
rect 25363 36329 25375 36363
rect 26694 36360 26700 36372
rect 25317 36323 25375 36329
rect 25976 36332 26700 36360
rect 19521 36295 19579 36301
rect 19521 36261 19533 36295
rect 19567 36261 19579 36295
rect 19521 36255 19579 36261
rect 19610 36252 19616 36304
rect 19668 36292 19674 36304
rect 19889 36295 19947 36301
rect 19668 36264 19840 36292
rect 19668 36252 19674 36264
rect 16301 36227 16359 36233
rect 16301 36193 16313 36227
rect 16347 36193 16359 36227
rect 16301 36187 16359 36193
rect 16390 36184 16396 36236
rect 16448 36224 16454 36236
rect 16577 36227 16635 36233
rect 16577 36224 16589 36227
rect 16448 36196 16589 36224
rect 16448 36184 16454 36196
rect 16577 36193 16589 36196
rect 16623 36193 16635 36227
rect 16577 36187 16635 36193
rect 15286 36156 15292 36168
rect 14384 36128 15292 36156
rect 15286 36116 15292 36128
rect 15344 36156 15350 36168
rect 15344 36128 16436 36156
rect 15344 36116 15350 36128
rect 10428 36060 12434 36088
rect 11793 36023 11851 36029
rect 11793 35989 11805 36023
rect 11839 36020 11851 36023
rect 11882 36020 11888 36032
rect 11839 35992 11888 36020
rect 11839 35989 11851 35992
rect 11793 35983 11851 35989
rect 11882 35980 11888 35992
rect 11940 35980 11946 36032
rect 12406 36020 12434 36060
rect 12544 36060 13400 36088
rect 12544 36020 12572 36060
rect 13630 36048 13636 36100
rect 13688 36088 13694 36100
rect 13998 36088 14004 36100
rect 13688 36060 14004 36088
rect 13688 36048 13694 36060
rect 13998 36048 14004 36060
rect 14056 36048 14062 36100
rect 16408 36032 16436 36128
rect 16482 36116 16488 36168
rect 16540 36116 16546 36168
rect 16592 36156 16620 36187
rect 16850 36184 16856 36236
rect 16908 36184 16914 36236
rect 17954 36184 17960 36236
rect 18012 36184 18018 36236
rect 18414 36224 18420 36236
rect 18064 36196 18420 36224
rect 18064 36156 18092 36196
rect 18414 36184 18420 36196
rect 18472 36224 18478 36236
rect 18782 36224 18788 36236
rect 18472 36196 18788 36224
rect 18472 36184 18478 36196
rect 18782 36184 18788 36196
rect 18840 36184 18846 36236
rect 19705 36227 19763 36233
rect 19705 36193 19717 36227
rect 19751 36193 19763 36227
rect 19812 36224 19840 36264
rect 19889 36261 19901 36295
rect 19935 36292 19947 36295
rect 23359 36295 23417 36301
rect 19935 36264 20208 36292
rect 19935 36261 19947 36264
rect 19889 36255 19947 36261
rect 20180 36233 20208 36264
rect 23359 36261 23371 36295
rect 23405 36292 23417 36295
rect 23492 36292 23520 36320
rect 24136 36292 24164 36320
rect 24673 36295 24731 36301
rect 24673 36292 24685 36295
rect 23405 36264 23796 36292
rect 24136 36264 24685 36292
rect 23405 36261 23417 36264
rect 23359 36255 23417 36261
rect 19981 36227 20039 36233
rect 19981 36224 19993 36227
rect 19812 36196 19993 36224
rect 19705 36187 19763 36193
rect 19981 36193 19993 36196
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 20165 36227 20223 36233
rect 20165 36193 20177 36227
rect 20211 36193 20223 36227
rect 20165 36187 20223 36193
rect 16592 36128 18092 36156
rect 18138 36116 18144 36168
rect 18196 36156 18202 36168
rect 18233 36159 18291 36165
rect 18233 36156 18245 36159
rect 18196 36128 18245 36156
rect 18196 36116 18202 36128
rect 18233 36125 18245 36128
rect 18279 36125 18291 36159
rect 18233 36119 18291 36125
rect 18322 36116 18328 36168
rect 18380 36156 18386 36168
rect 18506 36156 18512 36168
rect 18380 36128 18512 36156
rect 18380 36116 18386 36128
rect 18506 36116 18512 36128
rect 18564 36156 18570 36168
rect 19242 36156 19248 36168
rect 18564 36128 19248 36156
rect 18564 36116 18570 36128
rect 19242 36116 19248 36128
rect 19300 36156 19306 36168
rect 19720 36156 19748 36187
rect 20254 36184 20260 36236
rect 20312 36184 20318 36236
rect 20349 36227 20407 36233
rect 20349 36193 20361 36227
rect 20395 36224 20407 36227
rect 20806 36224 20812 36236
rect 20395 36196 20812 36224
rect 20395 36193 20407 36196
rect 20349 36187 20407 36193
rect 19300 36128 19748 36156
rect 19300 36116 19306 36128
rect 16500 36088 16528 36116
rect 19518 36088 19524 36100
rect 16500 36060 19524 36088
rect 12406 35992 12572 36020
rect 12618 35980 12624 36032
rect 12676 35980 12682 36032
rect 13906 35980 13912 36032
rect 13964 36020 13970 36032
rect 14185 36023 14243 36029
rect 14185 36020 14197 36023
rect 13964 35992 14197 36020
rect 13964 35980 13970 35992
rect 14185 35989 14197 35992
rect 14231 36020 14243 36023
rect 14734 36020 14740 36032
rect 14231 35992 14740 36020
rect 14231 35989 14243 35992
rect 14185 35983 14243 35989
rect 14734 35980 14740 35992
rect 14792 35980 14798 36032
rect 16390 35980 16396 36032
rect 16448 35980 16454 36032
rect 16482 35980 16488 36032
rect 16540 36020 16546 36032
rect 18432 36029 18460 36060
rect 19518 36048 19524 36060
rect 19576 36048 19582 36100
rect 17037 36023 17095 36029
rect 17037 36020 17049 36023
rect 16540 35992 17049 36020
rect 16540 35980 16546 35992
rect 17037 35989 17049 35992
rect 17083 35989 17095 36023
rect 17037 35983 17095 35989
rect 18417 36023 18475 36029
rect 18417 35989 18429 36023
rect 18463 35989 18475 36023
rect 18417 35983 18475 35989
rect 18601 36023 18659 36029
rect 18601 35989 18613 36023
rect 18647 36020 18659 36023
rect 18690 36020 18696 36032
rect 18647 35992 18696 36020
rect 18647 35989 18659 35992
rect 18601 35983 18659 35989
rect 18690 35980 18696 35992
rect 18748 35980 18754 36032
rect 18966 35980 18972 36032
rect 19024 36020 19030 36032
rect 20364 36020 20392 36187
rect 20806 36184 20812 36196
rect 20864 36184 20870 36236
rect 21542 36184 21548 36236
rect 21600 36184 21606 36236
rect 22097 36227 22155 36233
rect 22097 36193 22109 36227
rect 22143 36224 22155 36227
rect 22370 36224 22376 36236
rect 22143 36196 22376 36224
rect 22143 36193 22155 36196
rect 22097 36187 22155 36193
rect 22370 36184 22376 36196
rect 22428 36184 22434 36236
rect 22554 36184 22560 36236
rect 22612 36184 22618 36236
rect 23474 36184 23480 36236
rect 23532 36184 23538 36236
rect 23569 36227 23627 36233
rect 23569 36193 23581 36227
rect 23615 36193 23627 36227
rect 23569 36187 23627 36193
rect 23198 36116 23204 36168
rect 23256 36116 23262 36168
rect 23584 36156 23612 36187
rect 23658 36184 23664 36236
rect 23716 36184 23722 36236
rect 23768 36224 23796 36264
rect 24673 36261 24685 36264
rect 24719 36261 24731 36295
rect 24673 36255 24731 36261
rect 25133 36295 25191 36301
rect 25133 36261 25145 36295
rect 25179 36292 25191 36295
rect 25222 36292 25228 36304
rect 25179 36264 25228 36292
rect 25179 36261 25191 36264
rect 25133 36255 25191 36261
rect 25222 36252 25228 36264
rect 25280 36252 25286 36304
rect 25774 36252 25780 36304
rect 25832 36292 25838 36304
rect 25976 36292 26004 36332
rect 26694 36320 26700 36332
rect 26752 36320 26758 36372
rect 30006 36320 30012 36372
rect 30064 36320 30070 36372
rect 30282 36320 30288 36372
rect 30340 36360 30346 36372
rect 30340 36332 30880 36360
rect 30340 36320 30346 36332
rect 30193 36295 30251 36301
rect 25832 36264 26004 36292
rect 25832 36252 25838 36264
rect 24118 36224 24124 36236
rect 23768 36196 24124 36224
rect 24118 36184 24124 36196
rect 24176 36233 24182 36236
rect 24176 36227 24225 36233
rect 24176 36193 24179 36227
rect 24213 36193 24225 36227
rect 24176 36187 24225 36193
rect 24305 36227 24363 36233
rect 24305 36193 24317 36227
rect 24351 36193 24363 36227
rect 24305 36187 24363 36193
rect 24397 36227 24455 36233
rect 24397 36193 24409 36227
rect 24443 36193 24455 36227
rect 24397 36187 24455 36193
rect 24489 36227 24547 36233
rect 24489 36193 24501 36227
rect 24535 36224 24547 36227
rect 24578 36224 24584 36236
rect 24535 36196 24584 36224
rect 24535 36193 24547 36196
rect 24489 36187 24547 36193
rect 24176 36184 24182 36187
rect 23842 36156 23848 36168
rect 23584 36128 23848 36156
rect 23842 36116 23848 36128
rect 23900 36116 23906 36168
rect 24026 36116 24032 36168
rect 24084 36116 24090 36168
rect 22278 36048 22284 36100
rect 22336 36048 22342 36100
rect 22830 36048 22836 36100
rect 22888 36088 22894 36100
rect 24320 36088 24348 36187
rect 22888 36060 24348 36088
rect 24412 36088 24440 36187
rect 24578 36184 24584 36196
rect 24636 36184 24642 36236
rect 24762 36184 24768 36236
rect 24820 36184 24826 36236
rect 24946 36184 24952 36236
rect 25004 36184 25010 36236
rect 25406 36184 25412 36236
rect 25464 36184 25470 36236
rect 25792 36088 25820 36252
rect 25976 36233 26004 36264
rect 26252 36264 26924 36292
rect 26252 36233 26280 36264
rect 26896 36236 26924 36264
rect 30193 36261 30205 36295
rect 30239 36292 30251 36295
rect 30653 36295 30711 36301
rect 30653 36292 30665 36295
rect 30239 36264 30665 36292
rect 30239 36261 30251 36264
rect 30193 36255 30251 36261
rect 30653 36261 30665 36264
rect 30699 36261 30711 36295
rect 30653 36255 30711 36261
rect 30852 36292 30880 36332
rect 31018 36320 31024 36372
rect 31076 36360 31082 36372
rect 31294 36360 31300 36372
rect 31076 36332 31300 36360
rect 31076 36320 31082 36332
rect 31294 36320 31300 36332
rect 31352 36320 31358 36372
rect 31680 36292 31708 36536
rect 30852 36264 31708 36292
rect 25869 36227 25927 36233
rect 25869 36193 25881 36227
rect 25915 36193 25927 36227
rect 25869 36187 25927 36193
rect 25961 36227 26019 36233
rect 25961 36193 25973 36227
rect 26007 36193 26019 36227
rect 25961 36187 26019 36193
rect 26237 36227 26295 36233
rect 26237 36193 26249 36227
rect 26283 36193 26295 36227
rect 26237 36187 26295 36193
rect 25884 36156 25912 36187
rect 26418 36184 26424 36236
rect 26476 36184 26482 36236
rect 26602 36224 26608 36236
rect 26528 36196 26608 36224
rect 26528 36156 26556 36196
rect 26602 36184 26608 36196
rect 26660 36184 26666 36236
rect 26694 36184 26700 36236
rect 26752 36184 26758 36236
rect 26786 36184 26792 36236
rect 26844 36184 26850 36236
rect 26878 36184 26884 36236
rect 26936 36224 26942 36236
rect 26973 36227 27031 36233
rect 26973 36224 26985 36227
rect 26936 36196 26985 36224
rect 26936 36184 26942 36196
rect 26973 36193 26985 36196
rect 27019 36193 27031 36227
rect 26973 36187 27031 36193
rect 30558 36184 30564 36236
rect 30616 36184 30622 36236
rect 30852 36233 30880 36264
rect 30837 36227 30895 36233
rect 30837 36193 30849 36227
rect 30883 36193 30895 36227
rect 30837 36187 30895 36193
rect 31113 36227 31171 36233
rect 31113 36193 31125 36227
rect 31159 36193 31171 36227
rect 31113 36187 31171 36193
rect 25884 36128 26556 36156
rect 24412 36060 25820 36088
rect 26145 36091 26203 36097
rect 22888 36048 22894 36060
rect 26145 36057 26157 36091
rect 26191 36088 26203 36091
rect 26804 36088 26832 36184
rect 29638 36116 29644 36168
rect 29696 36156 29702 36168
rect 30282 36156 30288 36168
rect 29696 36128 30288 36156
rect 29696 36116 29702 36128
rect 30282 36116 30288 36128
rect 30340 36156 30346 36168
rect 31128 36156 31156 36187
rect 30340 36128 31156 36156
rect 30340 36116 30346 36128
rect 26191 36060 26832 36088
rect 26191 36057 26203 36060
rect 26145 36051 26203 36057
rect 19024 35992 20392 36020
rect 19024 35980 19030 35992
rect 20622 35980 20628 36032
rect 20680 35980 20686 36032
rect 21361 36023 21419 36029
rect 21361 35989 21373 36023
rect 21407 36020 21419 36023
rect 21450 36020 21456 36032
rect 21407 35992 21456 36020
rect 21407 35989 21419 35992
rect 21361 35983 21419 35989
rect 21450 35980 21456 35992
rect 21508 35980 21514 36032
rect 21818 35980 21824 36032
rect 21876 36020 21882 36032
rect 22005 36023 22063 36029
rect 22005 36020 22017 36023
rect 21876 35992 22017 36020
rect 21876 35980 21882 35992
rect 22005 35989 22017 35992
rect 22051 35989 22063 36023
rect 22005 35983 22063 35989
rect 25682 35980 25688 36032
rect 25740 35980 25746 36032
rect 26786 35980 26792 36032
rect 26844 36020 26850 36032
rect 27065 36023 27123 36029
rect 27065 36020 27077 36023
rect 26844 35992 27077 36020
rect 26844 35980 26850 35992
rect 27065 35989 27077 35992
rect 27111 35989 27123 36023
rect 27065 35983 27123 35989
rect 29546 35980 29552 36032
rect 29604 36020 29610 36032
rect 30193 36023 30251 36029
rect 30193 36020 30205 36023
rect 29604 35992 30205 36020
rect 29604 35980 29610 35992
rect 30193 35989 30205 35992
rect 30239 36020 30251 36023
rect 30742 36020 30748 36032
rect 30239 35992 30748 36020
rect 30239 35989 30251 35992
rect 30193 35983 30251 35989
rect 30742 35980 30748 35992
rect 30800 35980 30806 36032
rect 552 35930 31648 35952
rect 552 35878 3662 35930
rect 3714 35878 3726 35930
rect 3778 35878 3790 35930
rect 3842 35878 3854 35930
rect 3906 35878 3918 35930
rect 3970 35878 11436 35930
rect 11488 35878 11500 35930
rect 11552 35878 11564 35930
rect 11616 35878 11628 35930
rect 11680 35878 11692 35930
rect 11744 35878 19210 35930
rect 19262 35878 19274 35930
rect 19326 35878 19338 35930
rect 19390 35878 19402 35930
rect 19454 35878 19466 35930
rect 19518 35878 26984 35930
rect 27036 35878 27048 35930
rect 27100 35878 27112 35930
rect 27164 35878 27176 35930
rect 27228 35878 27240 35930
rect 27292 35878 31648 35930
rect 552 35856 31648 35878
rect 10042 35776 10048 35828
rect 10100 35816 10106 35828
rect 12618 35816 12624 35828
rect 10100 35788 12624 35816
rect 10100 35776 10106 35788
rect 12618 35776 12624 35788
rect 12676 35776 12682 35828
rect 12710 35776 12716 35828
rect 12768 35776 12774 35828
rect 12802 35776 12808 35828
rect 12860 35816 12866 35828
rect 14642 35816 14648 35828
rect 12860 35788 14648 35816
rect 12860 35776 12866 35788
rect 14642 35776 14648 35788
rect 14700 35776 14706 35828
rect 17126 35816 17132 35828
rect 14752 35788 17132 35816
rect 12250 35708 12256 35760
rect 12308 35748 12314 35760
rect 14752 35748 14780 35788
rect 15746 35748 15752 35760
rect 12308 35720 14780 35748
rect 15212 35720 15752 35748
rect 12308 35708 12314 35720
rect 8294 35640 8300 35692
rect 8352 35680 8358 35692
rect 8352 35652 11008 35680
rect 8352 35640 8358 35652
rect 9490 35572 9496 35624
rect 9548 35572 9554 35624
rect 9677 35615 9735 35621
rect 9677 35581 9689 35615
rect 9723 35581 9735 35615
rect 9677 35575 9735 35581
rect 9692 35544 9720 35575
rect 9766 35572 9772 35624
rect 9824 35572 9830 35624
rect 9861 35615 9919 35621
rect 9861 35581 9873 35615
rect 9907 35612 9919 35615
rect 10134 35612 10140 35624
rect 9907 35584 10140 35612
rect 9907 35581 9919 35584
rect 9861 35575 9919 35581
rect 10134 35572 10140 35584
rect 10192 35572 10198 35624
rect 10980 35621 11008 35652
rect 12802 35640 12808 35692
rect 12860 35680 12866 35692
rect 13446 35680 13452 35692
rect 12860 35652 13452 35680
rect 12860 35640 12866 35652
rect 10965 35615 11023 35621
rect 10965 35581 10977 35615
rect 11011 35581 11023 35615
rect 10965 35575 11023 35581
rect 11057 35615 11115 35621
rect 11057 35581 11069 35615
rect 11103 35612 11115 35615
rect 11241 35615 11299 35621
rect 11241 35612 11253 35615
rect 11103 35584 11253 35612
rect 11103 35581 11115 35584
rect 11057 35575 11115 35581
rect 11241 35581 11253 35584
rect 11287 35581 11299 35615
rect 12989 35615 13047 35621
rect 12989 35612 13001 35615
rect 11241 35575 11299 35581
rect 12406 35584 13001 35612
rect 10502 35544 10508 35556
rect 9692 35516 10508 35544
rect 10502 35504 10508 35516
rect 10560 35504 10566 35556
rect 11514 35553 11520 35556
rect 11508 35507 11520 35553
rect 11514 35504 11520 35507
rect 11572 35504 11578 35556
rect 11698 35504 11704 35556
rect 11756 35544 11762 35556
rect 12406 35544 12434 35584
rect 12989 35581 13001 35584
rect 13035 35581 13047 35615
rect 12989 35575 13047 35581
rect 13078 35572 13084 35624
rect 13136 35572 13142 35624
rect 13188 35621 13216 35652
rect 13446 35640 13452 35652
rect 13504 35680 13510 35692
rect 15010 35680 15016 35692
rect 13504 35652 15016 35680
rect 13504 35640 13510 35652
rect 15010 35640 15016 35652
rect 15068 35640 15074 35692
rect 15212 35621 15240 35720
rect 15746 35708 15752 35720
rect 15804 35708 15810 35760
rect 15856 35680 15884 35788
rect 17126 35776 17132 35788
rect 17184 35776 17190 35828
rect 21542 35776 21548 35828
rect 21600 35816 21606 35828
rect 21729 35819 21787 35825
rect 21729 35816 21741 35819
rect 21600 35788 21741 35816
rect 21600 35776 21606 35788
rect 21729 35785 21741 35788
rect 21775 35785 21787 35819
rect 21729 35779 21787 35785
rect 22554 35776 22560 35828
rect 22612 35816 22618 35828
rect 23201 35819 23259 35825
rect 23201 35816 23213 35819
rect 22612 35788 23213 35816
rect 22612 35776 22618 35788
rect 23201 35785 23213 35788
rect 23247 35785 23259 35819
rect 23201 35779 23259 35785
rect 23658 35776 23664 35828
rect 23716 35816 23722 35828
rect 24029 35819 24087 35825
rect 24029 35816 24041 35819
rect 23716 35788 24041 35816
rect 23716 35776 23722 35788
rect 24029 35785 24041 35788
rect 24075 35816 24087 35819
rect 24578 35816 24584 35828
rect 24075 35788 24584 35816
rect 24075 35785 24087 35788
rect 24029 35779 24087 35785
rect 24578 35776 24584 35788
rect 24636 35776 24642 35828
rect 26510 35776 26516 35828
rect 26568 35816 26574 35828
rect 27154 35816 27160 35828
rect 26568 35788 27160 35816
rect 26568 35776 26574 35788
rect 27154 35776 27160 35788
rect 27212 35816 27218 35828
rect 28353 35819 28411 35825
rect 28353 35816 28365 35819
rect 27212 35788 28365 35816
rect 27212 35776 27218 35788
rect 28353 35785 28365 35788
rect 28399 35816 28411 35819
rect 28442 35816 28448 35828
rect 28399 35788 28448 35816
rect 28399 35785 28411 35788
rect 28353 35779 28411 35785
rect 28442 35776 28448 35788
rect 28500 35776 28506 35828
rect 16482 35748 16488 35760
rect 15396 35652 15884 35680
rect 15948 35720 16488 35748
rect 13173 35615 13231 35621
rect 13173 35581 13185 35615
rect 13219 35581 13231 35615
rect 13173 35575 13231 35581
rect 13357 35615 13415 35621
rect 13357 35581 13369 35615
rect 13403 35612 13415 35615
rect 13909 35615 13967 35621
rect 13909 35612 13921 35615
rect 13403 35584 13921 35612
rect 13403 35581 13415 35584
rect 13357 35575 13415 35581
rect 13909 35581 13921 35584
rect 13955 35581 13967 35615
rect 13909 35575 13967 35581
rect 15197 35615 15255 35621
rect 15197 35581 15209 35615
rect 15243 35581 15255 35615
rect 15197 35575 15255 35581
rect 15286 35572 15292 35624
rect 15344 35612 15350 35624
rect 15396 35621 15424 35652
rect 15381 35615 15439 35621
rect 15381 35612 15393 35615
rect 15344 35584 15393 35612
rect 15344 35572 15350 35584
rect 15381 35581 15393 35584
rect 15427 35581 15439 35615
rect 15381 35575 15439 35581
rect 15470 35572 15476 35624
rect 15528 35572 15534 35624
rect 15565 35615 15623 35621
rect 15565 35581 15577 35615
rect 15611 35581 15623 35615
rect 15565 35575 15623 35581
rect 13262 35544 13268 35556
rect 11756 35516 12434 35544
rect 12636 35516 13268 35544
rect 11756 35504 11762 35516
rect 10137 35479 10195 35485
rect 10137 35445 10149 35479
rect 10183 35476 10195 35479
rect 10318 35476 10324 35488
rect 10183 35448 10324 35476
rect 10183 35445 10195 35448
rect 10137 35439 10195 35445
rect 10318 35436 10324 35448
rect 10376 35436 10382 35488
rect 11606 35436 11612 35488
rect 11664 35476 11670 35488
rect 12636 35485 12664 35516
rect 13262 35504 13268 35516
rect 13320 35504 13326 35556
rect 13538 35504 13544 35556
rect 13596 35504 13602 35556
rect 13722 35504 13728 35556
rect 13780 35544 13786 35556
rect 15580 35544 15608 35575
rect 15654 35572 15660 35624
rect 15712 35612 15718 35624
rect 15948 35621 15976 35720
rect 16482 35708 16488 35720
rect 16540 35708 16546 35760
rect 16022 35640 16028 35692
rect 16080 35680 16086 35692
rect 16301 35683 16359 35689
rect 16301 35680 16313 35683
rect 16080 35652 16313 35680
rect 16080 35640 16086 35652
rect 16301 35649 16313 35652
rect 16347 35649 16359 35683
rect 16301 35643 16359 35649
rect 16408 35652 16896 35680
rect 15933 35615 15991 35621
rect 15933 35612 15945 35615
rect 15712 35584 15945 35612
rect 15712 35572 15718 35584
rect 15933 35581 15945 35584
rect 15979 35581 15991 35615
rect 15933 35575 15991 35581
rect 16117 35615 16175 35621
rect 16117 35581 16129 35615
rect 16163 35581 16175 35615
rect 16117 35575 16175 35581
rect 13780 35516 15608 35544
rect 15841 35547 15899 35553
rect 13780 35504 13786 35516
rect 15841 35513 15853 35547
rect 15887 35544 15899 35547
rect 16132 35544 16160 35575
rect 16206 35572 16212 35624
rect 16264 35572 16270 35624
rect 15887 35516 16160 35544
rect 15887 35513 15899 35516
rect 15841 35507 15899 35513
rect 12621 35479 12679 35485
rect 12621 35476 12633 35479
rect 11664 35448 12633 35476
rect 11664 35436 11670 35448
rect 12621 35445 12633 35448
rect 12667 35445 12679 35479
rect 12621 35439 12679 35445
rect 12894 35436 12900 35488
rect 12952 35476 12958 35488
rect 15470 35476 15476 35488
rect 12952 35448 15476 35476
rect 12952 35436 12958 35448
rect 15470 35436 15476 35448
rect 15528 35476 15534 35488
rect 16408 35476 16436 35652
rect 16482 35572 16488 35624
rect 16540 35572 16546 35624
rect 16758 35572 16764 35624
rect 16816 35572 16822 35624
rect 16868 35612 16896 35652
rect 21818 35640 21824 35692
rect 21876 35640 21882 35692
rect 26878 35640 26884 35692
rect 26936 35680 26942 35692
rect 26936 35652 27936 35680
rect 26936 35640 26942 35652
rect 16868 35584 17172 35612
rect 16669 35547 16727 35553
rect 16669 35513 16681 35547
rect 16715 35544 16727 35547
rect 17006 35547 17064 35553
rect 17006 35544 17018 35547
rect 16715 35516 17018 35544
rect 16715 35513 16727 35516
rect 16669 35507 16727 35513
rect 17006 35513 17018 35516
rect 17052 35513 17064 35547
rect 17144 35544 17172 35584
rect 18598 35572 18604 35624
rect 18656 35612 18662 35624
rect 19061 35615 19119 35621
rect 19061 35612 19073 35615
rect 18656 35584 19073 35612
rect 18656 35572 18662 35584
rect 19061 35581 19073 35584
rect 19107 35581 19119 35615
rect 19061 35575 19119 35581
rect 19794 35572 19800 35624
rect 19852 35612 19858 35624
rect 20622 35621 20628 35624
rect 20073 35615 20131 35621
rect 20073 35612 20085 35615
rect 19852 35584 20085 35612
rect 19852 35572 19858 35584
rect 20073 35581 20085 35584
rect 20119 35581 20131 35615
rect 20073 35575 20131 35581
rect 20165 35615 20223 35621
rect 20165 35581 20177 35615
rect 20211 35612 20223 35615
rect 20349 35615 20407 35621
rect 20349 35612 20361 35615
rect 20211 35584 20361 35612
rect 20211 35581 20223 35584
rect 20165 35575 20223 35581
rect 20349 35581 20361 35584
rect 20395 35581 20407 35615
rect 20616 35612 20628 35621
rect 20583 35584 20628 35612
rect 20349 35575 20407 35581
rect 20616 35575 20628 35584
rect 20622 35572 20628 35575
rect 20680 35572 20686 35624
rect 23845 35615 23903 35621
rect 23845 35612 23857 35615
rect 20824 35584 23857 35612
rect 20824 35556 20852 35584
rect 23845 35581 23857 35584
rect 23891 35612 23903 35615
rect 23934 35612 23940 35624
rect 23891 35584 23940 35612
rect 23891 35581 23903 35584
rect 23845 35575 23903 35581
rect 23934 35572 23940 35584
rect 23992 35572 23998 35624
rect 24029 35615 24087 35621
rect 24029 35581 24041 35615
rect 24075 35612 24087 35615
rect 24118 35612 24124 35624
rect 24075 35584 24124 35612
rect 24075 35581 24087 35584
rect 24029 35575 24087 35581
rect 24118 35572 24124 35584
rect 24176 35572 24182 35624
rect 26694 35572 26700 35624
rect 26752 35612 26758 35624
rect 27801 35615 27859 35621
rect 27801 35612 27813 35615
rect 26752 35584 27813 35612
rect 26752 35572 26758 35584
rect 27801 35581 27813 35584
rect 27847 35581 27859 35615
rect 27908 35612 27936 35652
rect 27982 35640 27988 35692
rect 28040 35680 28046 35692
rect 28902 35680 28908 35692
rect 28040 35652 28908 35680
rect 28040 35640 28046 35652
rect 28902 35640 28908 35652
rect 28960 35640 28966 35692
rect 28077 35615 28135 35621
rect 28077 35612 28089 35615
rect 27908 35584 28089 35612
rect 27801 35575 27859 35581
rect 28077 35581 28089 35584
rect 28123 35612 28135 35615
rect 29638 35612 29644 35624
rect 28123 35584 29644 35612
rect 28123 35581 28135 35584
rect 28077 35575 28135 35581
rect 29638 35572 29644 35584
rect 29696 35572 29702 35624
rect 17144 35516 18828 35544
rect 17006 35507 17064 35513
rect 18800 35488 18828 35516
rect 20806 35504 20812 35556
rect 20864 35504 20870 35556
rect 22088 35547 22146 35553
rect 22088 35513 22100 35547
rect 22134 35544 22146 35547
rect 22186 35544 22192 35556
rect 22134 35516 22192 35544
rect 22134 35513 22146 35516
rect 22088 35507 22146 35513
rect 22186 35504 22192 35516
rect 22244 35504 22250 35556
rect 25314 35504 25320 35556
rect 25372 35544 25378 35556
rect 28261 35547 28319 35553
rect 28261 35544 28273 35547
rect 25372 35516 28273 35544
rect 25372 35504 25378 35516
rect 28261 35513 28273 35516
rect 28307 35513 28319 35547
rect 28261 35507 28319 35513
rect 15528 35448 16436 35476
rect 15528 35436 15534 35448
rect 16482 35436 16488 35488
rect 16540 35476 16546 35488
rect 18138 35476 18144 35488
rect 16540 35448 18144 35476
rect 16540 35436 16546 35448
rect 18138 35436 18144 35448
rect 18196 35436 18202 35488
rect 18782 35436 18788 35488
rect 18840 35476 18846 35488
rect 18969 35479 19027 35485
rect 18969 35476 18981 35479
rect 18840 35448 18981 35476
rect 18840 35436 18846 35448
rect 18969 35445 18981 35448
rect 19015 35445 19027 35479
rect 18969 35439 19027 35445
rect 19702 35436 19708 35488
rect 19760 35476 19766 35488
rect 20254 35476 20260 35488
rect 19760 35448 20260 35476
rect 19760 35436 19766 35448
rect 20254 35436 20260 35448
rect 20312 35436 20318 35488
rect 27246 35436 27252 35488
rect 27304 35476 27310 35488
rect 27617 35479 27675 35485
rect 27617 35476 27629 35479
rect 27304 35448 27629 35476
rect 27304 35436 27310 35448
rect 27617 35445 27629 35448
rect 27663 35445 27675 35479
rect 27617 35439 27675 35445
rect 27982 35436 27988 35488
rect 28040 35436 28046 35488
rect 28442 35436 28448 35488
rect 28500 35476 28506 35488
rect 30834 35476 30840 35488
rect 28500 35448 30840 35476
rect 28500 35436 28506 35448
rect 30834 35436 30840 35448
rect 30892 35436 30898 35488
rect 552 35386 31648 35408
rect 552 35334 4322 35386
rect 4374 35334 4386 35386
rect 4438 35334 4450 35386
rect 4502 35334 4514 35386
rect 4566 35334 4578 35386
rect 4630 35334 12096 35386
rect 12148 35334 12160 35386
rect 12212 35334 12224 35386
rect 12276 35334 12288 35386
rect 12340 35334 12352 35386
rect 12404 35334 19870 35386
rect 19922 35334 19934 35386
rect 19986 35334 19998 35386
rect 20050 35334 20062 35386
rect 20114 35334 20126 35386
rect 20178 35334 27644 35386
rect 27696 35334 27708 35386
rect 27760 35334 27772 35386
rect 27824 35334 27836 35386
rect 27888 35334 27900 35386
rect 27952 35334 31648 35386
rect 552 35312 31648 35334
rect 9953 35275 10011 35281
rect 9953 35241 9965 35275
rect 9999 35272 10011 35275
rect 10134 35272 10140 35284
rect 9999 35244 10140 35272
rect 9999 35241 10011 35244
rect 9953 35235 10011 35241
rect 10134 35232 10140 35244
rect 10192 35232 10198 35284
rect 11425 35275 11483 35281
rect 11425 35241 11437 35275
rect 11471 35272 11483 35275
rect 11514 35272 11520 35284
rect 11471 35244 11520 35272
rect 11471 35241 11483 35244
rect 11425 35235 11483 35241
rect 11514 35232 11520 35244
rect 11572 35232 11578 35284
rect 11974 35232 11980 35284
rect 12032 35272 12038 35284
rect 12161 35275 12219 35281
rect 12161 35272 12173 35275
rect 12032 35244 12173 35272
rect 12032 35232 12038 35244
rect 12161 35241 12173 35244
rect 12207 35241 12219 35275
rect 15470 35272 15476 35284
rect 12161 35235 12219 35241
rect 13280 35244 15476 35272
rect 12618 35164 12624 35216
rect 12676 35204 12682 35216
rect 12676 35176 12940 35204
rect 12676 35164 12682 35176
rect 10042 35136 10048 35148
rect 9692 35108 10048 35136
rect 9692 35077 9720 35108
rect 10042 35096 10048 35108
rect 10100 35096 10106 35148
rect 11606 35096 11612 35148
rect 11664 35136 11670 35148
rect 11701 35139 11759 35145
rect 11701 35136 11713 35139
rect 11664 35108 11713 35136
rect 11664 35096 11670 35108
rect 11701 35105 11713 35108
rect 11747 35105 11759 35139
rect 11701 35099 11759 35105
rect 11793 35139 11851 35145
rect 11793 35105 11805 35139
rect 11839 35105 11851 35139
rect 11793 35099 11851 35105
rect 9677 35071 9735 35077
rect 9677 35037 9689 35071
rect 9723 35037 9735 35071
rect 9677 35031 9735 35037
rect 9766 35028 9772 35080
rect 9824 35068 9830 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9824 35040 9873 35068
rect 9824 35028 9830 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 11238 35028 11244 35080
rect 11296 35068 11302 35080
rect 11808 35068 11836 35099
rect 11882 35096 11888 35148
rect 11940 35096 11946 35148
rect 12066 35096 12072 35148
rect 12124 35096 12130 35148
rect 12158 35096 12164 35148
rect 12216 35136 12222 35148
rect 12529 35139 12587 35145
rect 12529 35136 12541 35139
rect 12216 35108 12541 35136
rect 12216 35096 12222 35108
rect 12529 35105 12541 35108
rect 12575 35105 12587 35139
rect 12529 35099 12587 35105
rect 12621 35071 12679 35077
rect 11296 35040 11928 35068
rect 11296 35028 11302 35040
rect 11900 35000 11928 35040
rect 12621 35037 12633 35071
rect 12667 35068 12679 35071
rect 12710 35068 12716 35080
rect 12667 35040 12716 35068
rect 12667 35037 12679 35040
rect 12621 35031 12679 35037
rect 12710 35028 12716 35040
rect 12768 35028 12774 35080
rect 12805 35071 12863 35077
rect 12805 35037 12817 35071
rect 12851 35068 12863 35071
rect 12912 35068 12940 35176
rect 13280 35145 13308 35244
rect 15470 35232 15476 35244
rect 15528 35232 15534 35284
rect 16206 35232 16212 35284
rect 16264 35272 16270 35284
rect 16577 35275 16635 35281
rect 16577 35272 16589 35275
rect 16264 35244 16589 35272
rect 16264 35232 16270 35244
rect 16577 35241 16589 35244
rect 16623 35241 16635 35275
rect 16577 35235 16635 35241
rect 16758 35232 16764 35284
rect 16816 35272 16822 35284
rect 16945 35275 17003 35281
rect 16945 35272 16957 35275
rect 16816 35244 16957 35272
rect 16816 35232 16822 35244
rect 16945 35241 16957 35244
rect 16991 35241 17003 35275
rect 16945 35235 17003 35241
rect 19061 35275 19119 35281
rect 19061 35241 19073 35275
rect 19107 35272 19119 35275
rect 19794 35272 19800 35284
rect 19107 35244 19800 35272
rect 19107 35241 19119 35244
rect 19061 35235 19119 35241
rect 19794 35232 19800 35244
rect 19852 35232 19858 35284
rect 22186 35232 22192 35284
rect 22244 35232 22250 35284
rect 22465 35275 22523 35281
rect 22465 35241 22477 35275
rect 22511 35241 22523 35275
rect 22465 35235 22523 35241
rect 14093 35207 14151 35213
rect 14093 35204 14105 35207
rect 13556 35176 14105 35204
rect 13265 35139 13323 35145
rect 13265 35105 13277 35139
rect 13311 35105 13323 35139
rect 13265 35099 13323 35105
rect 13354 35096 13360 35148
rect 13412 35096 13418 35148
rect 13556 35145 13584 35176
rect 14093 35173 14105 35176
rect 14139 35173 14151 35207
rect 14093 35167 14151 35173
rect 15010 35164 15016 35216
rect 15068 35204 15074 35216
rect 18417 35207 18475 35213
rect 15068 35176 16252 35204
rect 15068 35164 15074 35176
rect 13541 35139 13599 35145
rect 13541 35105 13553 35139
rect 13587 35105 13599 35139
rect 13541 35099 13599 35105
rect 13630 35096 13636 35148
rect 13688 35096 13694 35148
rect 13722 35096 13728 35148
rect 13780 35096 13786 35148
rect 14274 35096 14280 35148
rect 14332 35096 14338 35148
rect 14369 35139 14427 35145
rect 14369 35105 14381 35139
rect 14415 35136 14427 35139
rect 14415 35108 14504 35136
rect 14415 35105 14427 35108
rect 14369 35099 14427 35105
rect 12851 35040 12940 35068
rect 12851 35037 12863 35040
rect 12805 35031 12863 35037
rect 13630 35000 13636 35012
rect 11900 34972 13636 35000
rect 13630 34960 13636 34972
rect 13688 34960 13694 35012
rect 10042 34892 10048 34944
rect 10100 34932 10106 34944
rect 10321 34935 10379 34941
rect 10321 34932 10333 34935
rect 10100 34904 10333 34932
rect 10100 34892 10106 34904
rect 10321 34901 10333 34904
rect 10367 34901 10379 34935
rect 10321 34895 10379 34901
rect 11698 34892 11704 34944
rect 11756 34932 11762 34944
rect 11882 34932 11888 34944
rect 11756 34904 11888 34932
rect 11756 34892 11762 34904
rect 11882 34892 11888 34904
rect 11940 34932 11946 34944
rect 12158 34932 12164 34944
rect 11940 34904 12164 34932
rect 11940 34892 11946 34904
rect 12158 34892 12164 34904
rect 12216 34892 12222 34944
rect 13081 34935 13139 34941
rect 13081 34901 13093 34935
rect 13127 34932 13139 34935
rect 13446 34932 13452 34944
rect 13127 34904 13452 34932
rect 13127 34901 13139 34904
rect 13081 34895 13139 34901
rect 13446 34892 13452 34904
rect 13504 34892 13510 34944
rect 13906 34892 13912 34944
rect 13964 34932 13970 34944
rect 14001 34935 14059 34941
rect 14001 34932 14013 34935
rect 13964 34904 14013 34932
rect 13964 34892 13970 34904
rect 14001 34901 14013 34904
rect 14047 34901 14059 34935
rect 14476 34932 14504 35108
rect 14550 35096 14556 35148
rect 14608 35096 14614 35148
rect 14642 35096 14648 35148
rect 14700 35096 14706 35148
rect 14734 35096 14740 35148
rect 14792 35096 14798 35148
rect 15102 35096 15108 35148
rect 15160 35136 15166 35148
rect 16224 35145 16252 35176
rect 18417 35173 18429 35207
rect 18463 35204 18475 35207
rect 18690 35204 18696 35216
rect 18463 35176 18696 35204
rect 18463 35173 18475 35176
rect 18417 35167 18475 35173
rect 18690 35164 18696 35176
rect 18748 35204 18754 35216
rect 21821 35207 21879 35213
rect 18748 35176 19748 35204
rect 18748 35164 18754 35176
rect 16117 35139 16175 35145
rect 16117 35136 16129 35139
rect 15160 35108 16129 35136
rect 15160 35096 15166 35108
rect 16117 35105 16129 35108
rect 16163 35105 16175 35139
rect 16117 35099 16175 35105
rect 16209 35139 16267 35145
rect 16209 35105 16221 35139
rect 16255 35105 16267 35139
rect 16209 35099 16267 35105
rect 16390 35096 16396 35148
rect 16448 35096 16454 35148
rect 16942 35096 16948 35148
rect 17000 35136 17006 35148
rect 17037 35139 17095 35145
rect 17037 35136 17049 35139
rect 17000 35108 17049 35136
rect 17000 35096 17006 35108
rect 17037 35105 17049 35108
rect 17083 35105 17095 35139
rect 17037 35099 17095 35105
rect 18782 35096 18788 35148
rect 18840 35096 18846 35148
rect 19720 35145 19748 35176
rect 21821 35173 21833 35207
rect 21867 35204 21879 35207
rect 21910 35204 21916 35216
rect 21867 35176 21916 35204
rect 21867 35173 21879 35176
rect 21821 35167 21879 35173
rect 21910 35164 21916 35176
rect 21968 35164 21974 35216
rect 22037 35207 22095 35213
rect 22037 35173 22049 35207
rect 22083 35204 22095 35207
rect 22480 35204 22508 35235
rect 22554 35232 22560 35284
rect 22612 35272 22618 35284
rect 22833 35275 22891 35281
rect 22833 35272 22845 35275
rect 22612 35244 22845 35272
rect 22612 35232 22618 35244
rect 22833 35241 22845 35244
rect 22879 35241 22891 35275
rect 22833 35235 22891 35241
rect 25314 35232 25320 35284
rect 25372 35232 25378 35284
rect 26973 35275 27031 35281
rect 26973 35241 26985 35275
rect 27019 35272 27031 35275
rect 27019 35244 27108 35272
rect 27019 35241 27031 35244
rect 26973 35235 27031 35241
rect 22083 35176 22508 35204
rect 22083 35173 22095 35176
rect 22037 35167 22095 35173
rect 26694 35164 26700 35216
rect 26752 35164 26758 35216
rect 26878 35164 26884 35216
rect 26936 35164 26942 35216
rect 27080 35213 27108 35244
rect 27246 35232 27252 35284
rect 27304 35281 27310 35284
rect 27304 35275 27323 35281
rect 27311 35241 27323 35275
rect 27304 35235 27323 35241
rect 27525 35275 27583 35281
rect 27525 35241 27537 35275
rect 27571 35272 27583 35275
rect 28074 35272 28080 35284
rect 27571 35244 28080 35272
rect 27571 35241 27583 35244
rect 27525 35235 27583 35241
rect 27304 35232 27310 35235
rect 28074 35232 28080 35244
rect 28132 35232 28138 35284
rect 29178 35232 29184 35284
rect 29236 35272 29242 35284
rect 30009 35275 30067 35281
rect 30009 35272 30021 35275
rect 29236 35244 30021 35272
rect 29236 35232 29242 35244
rect 30009 35241 30021 35244
rect 30055 35272 30067 35275
rect 30282 35272 30288 35284
rect 30055 35244 30288 35272
rect 30055 35241 30067 35244
rect 30009 35235 30067 35241
rect 30282 35232 30288 35244
rect 30340 35272 30346 35284
rect 30340 35244 30512 35272
rect 30340 35232 30346 35244
rect 27065 35207 27123 35213
rect 27065 35173 27077 35207
rect 27111 35173 27123 35207
rect 29825 35207 29883 35213
rect 29825 35204 29837 35207
rect 27065 35167 27123 35173
rect 29564 35176 29837 35204
rect 18877 35139 18935 35145
rect 18877 35105 18889 35139
rect 18923 35136 18935 35139
rect 19521 35139 19579 35145
rect 19521 35136 19533 35139
rect 18923 35108 19533 35136
rect 18923 35105 18935 35108
rect 18877 35099 18935 35105
rect 19521 35105 19533 35108
rect 19567 35105 19579 35139
rect 19521 35099 19579 35105
rect 19705 35139 19763 35145
rect 19705 35105 19717 35139
rect 19751 35105 19763 35139
rect 19705 35099 19763 35105
rect 19797 35139 19855 35145
rect 19797 35105 19809 35139
rect 19843 35136 19855 35139
rect 19843 35108 20668 35136
rect 19843 35105 19855 35108
rect 19797 35099 19855 35105
rect 14660 35000 14688 35096
rect 18046 35028 18052 35080
rect 18104 35068 18110 35080
rect 18892 35068 18920 35099
rect 18104 35040 18920 35068
rect 19536 35068 19564 35099
rect 20640 35068 20668 35108
rect 20714 35096 20720 35148
rect 20772 35136 20778 35148
rect 24581 35139 24639 35145
rect 24581 35136 24593 35139
rect 20772 35108 24593 35136
rect 20772 35096 20778 35108
rect 24581 35105 24593 35108
rect 24627 35105 24639 35139
rect 24581 35099 24639 35105
rect 24765 35139 24823 35145
rect 24765 35105 24777 35139
rect 24811 35136 24823 35139
rect 24854 35136 24860 35148
rect 24811 35108 24860 35136
rect 24811 35105 24823 35108
rect 24765 35099 24823 35105
rect 20806 35068 20812 35080
rect 19536 35040 19840 35068
rect 20640 35040 20812 35068
rect 18104 35028 18110 35040
rect 14921 35003 14979 35009
rect 14921 35000 14933 35003
rect 14660 34972 14933 35000
rect 14921 34969 14933 34972
rect 14967 34969 14979 35003
rect 14921 34963 14979 34969
rect 16022 34960 16028 35012
rect 16080 35000 16086 35012
rect 17402 35000 17408 35012
rect 16080 34972 17408 35000
rect 16080 34960 16086 34972
rect 17402 34960 17408 34972
rect 17460 34960 17466 35012
rect 18874 35000 18880 35012
rect 18800 34972 18880 35000
rect 15286 34932 15292 34944
rect 14476 34904 15292 34932
rect 14001 34895 14059 34901
rect 15286 34892 15292 34904
rect 15344 34892 15350 34944
rect 15470 34892 15476 34944
rect 15528 34932 15534 34944
rect 17218 34932 17224 34944
rect 15528 34904 17224 34932
rect 15528 34892 15534 34904
rect 17218 34892 17224 34904
rect 17276 34892 17282 34944
rect 18800 34941 18828 34972
rect 18874 34960 18880 34972
rect 18932 35000 18938 35012
rect 19613 35003 19671 35009
rect 19613 35000 19625 35003
rect 18932 34972 19625 35000
rect 18932 34960 18938 34972
rect 19613 34969 19625 34972
rect 19659 35000 19671 35003
rect 19702 35000 19708 35012
rect 19659 34972 19708 35000
rect 19659 34969 19671 34972
rect 19613 34963 19671 34969
rect 19702 34960 19708 34972
rect 19760 34960 19766 35012
rect 19812 35000 19840 35040
rect 20806 35028 20812 35040
rect 20864 35028 20870 35080
rect 22922 35028 22928 35080
rect 22980 35028 22986 35080
rect 23109 35071 23167 35077
rect 23109 35037 23121 35071
rect 23155 35068 23167 35071
rect 23842 35068 23848 35080
rect 23155 35040 23848 35068
rect 23155 35037 23167 35040
rect 23109 35031 23167 35037
rect 23842 35028 23848 35040
rect 23900 35028 23906 35080
rect 24596 35068 24624 35099
rect 24854 35096 24860 35108
rect 24912 35096 24918 35148
rect 25225 35139 25283 35145
rect 25225 35105 25237 35139
rect 25271 35105 25283 35139
rect 25225 35099 25283 35105
rect 25409 35139 25467 35145
rect 25409 35105 25421 35139
rect 25455 35136 25467 35139
rect 25682 35136 25688 35148
rect 25455 35108 25688 35136
rect 25455 35105 25467 35108
rect 25409 35099 25467 35105
rect 25038 35068 25044 35080
rect 24596 35040 25044 35068
rect 25038 35028 25044 35040
rect 25096 35068 25102 35080
rect 25240 35068 25268 35099
rect 25682 35096 25688 35108
rect 25740 35096 25746 35148
rect 26973 35139 27031 35145
rect 26973 35105 26985 35139
rect 27019 35105 27031 35139
rect 26973 35099 27031 35105
rect 25096 35040 25268 35068
rect 26988 35068 27016 35099
rect 28166 35096 28172 35148
rect 28224 35096 28230 35148
rect 28350 35145 28356 35148
rect 28307 35139 28356 35145
rect 28307 35105 28319 35139
rect 28353 35105 28356 35139
rect 28307 35099 28356 35105
rect 28350 35096 28356 35099
rect 28408 35096 28414 35148
rect 29564 35136 29592 35176
rect 29825 35173 29837 35176
rect 29871 35204 29883 35207
rect 30190 35204 30196 35216
rect 29871 35176 30196 35204
rect 29871 35173 29883 35176
rect 29825 35167 29883 35173
rect 30190 35164 30196 35176
rect 30248 35164 30254 35216
rect 29638 35136 29644 35148
rect 29104 35108 29592 35136
rect 27982 35068 27988 35080
rect 26988 35040 27988 35068
rect 25096 35028 25102 35040
rect 27982 35028 27988 35040
rect 28040 35028 28046 35080
rect 28445 35071 28503 35077
rect 28445 35037 28457 35071
rect 28491 35068 28503 35071
rect 29104 35068 29132 35108
rect 29636 35096 29644 35136
rect 29696 35096 29702 35148
rect 29730 35096 29736 35148
rect 29788 35096 29794 35148
rect 30484 35145 30512 35244
rect 30745 35207 30803 35213
rect 30745 35173 30757 35207
rect 30791 35204 30803 35207
rect 30837 35207 30895 35213
rect 30837 35204 30849 35207
rect 30791 35176 30849 35204
rect 30791 35173 30803 35176
rect 30745 35167 30803 35173
rect 30837 35173 30849 35176
rect 30883 35173 30895 35207
rect 30837 35167 30895 35173
rect 30101 35139 30159 35145
rect 30101 35105 30113 35139
rect 30147 35105 30159 35139
rect 30101 35099 30159 35105
rect 30469 35139 30527 35145
rect 30469 35105 30481 35139
rect 30515 35105 30527 35139
rect 30469 35099 30527 35105
rect 28491 35040 29132 35068
rect 29181 35071 29239 35077
rect 28491 35037 28503 35040
rect 28445 35031 28503 35037
rect 29181 35037 29193 35071
rect 29227 35037 29239 35071
rect 29181 35031 29239 35037
rect 29365 35071 29423 35077
rect 29365 35037 29377 35071
rect 29411 35068 29423 35071
rect 29636 35068 29664 35096
rect 30116 35068 30144 35099
rect 29411 35040 29664 35068
rect 29748 35040 30144 35068
rect 29411 35037 29423 35040
rect 29365 35031 29423 35037
rect 22738 35000 22744 35012
rect 19812 34972 22744 35000
rect 22738 34960 22744 34972
rect 22796 35000 22802 35012
rect 24026 35000 24032 35012
rect 22796 34972 24032 35000
rect 22796 34960 22802 34972
rect 24026 34960 24032 34972
rect 24084 34960 24090 35012
rect 24765 35003 24823 35009
rect 24765 34969 24777 35003
rect 24811 35000 24823 35003
rect 24811 34972 27844 35000
rect 24811 34969 24823 34972
rect 24765 34963 24823 34969
rect 18785 34935 18843 34941
rect 18785 34901 18797 34935
rect 18831 34901 18843 34935
rect 18785 34895 18843 34901
rect 19337 34935 19395 34941
rect 19337 34901 19349 34935
rect 19383 34932 19395 34935
rect 19886 34932 19892 34944
rect 19383 34904 19892 34932
rect 19383 34901 19395 34904
rect 19337 34895 19395 34901
rect 19886 34892 19892 34904
rect 19944 34892 19950 34944
rect 22005 34935 22063 34941
rect 22005 34901 22017 34935
rect 22051 34932 22063 34935
rect 22094 34932 22100 34944
rect 22051 34904 22100 34932
rect 22051 34901 22063 34904
rect 22005 34895 22063 34901
rect 22094 34892 22100 34904
rect 22152 34892 22158 34944
rect 27154 34892 27160 34944
rect 27212 34932 27218 34944
rect 27249 34935 27307 34941
rect 27249 34932 27261 34935
rect 27212 34904 27261 34932
rect 27212 34892 27218 34904
rect 27249 34901 27261 34904
rect 27295 34901 27307 34935
rect 27249 34895 27307 34901
rect 27338 34892 27344 34944
rect 27396 34932 27402 34944
rect 27433 34935 27491 34941
rect 27433 34932 27445 34935
rect 27396 34904 27445 34932
rect 27396 34892 27402 34904
rect 27433 34901 27445 34904
rect 27479 34901 27491 34935
rect 27816 34932 27844 34972
rect 28718 34960 28724 35012
rect 28776 34960 28782 35012
rect 28902 34960 28908 35012
rect 28960 35000 28966 35012
rect 29196 35000 29224 35031
rect 29457 35003 29515 35009
rect 29457 35000 29469 35003
rect 28960 34972 29469 35000
rect 28960 34960 28966 34972
rect 29457 34969 29469 34972
rect 29503 34969 29515 35003
rect 29457 34963 29515 34969
rect 27982 34932 27988 34944
rect 27816 34904 27988 34932
rect 27433 34895 27491 34901
rect 27982 34892 27988 34904
rect 28040 34892 28046 34944
rect 28626 34892 28632 34944
rect 28684 34932 28690 34944
rect 29748 34932 29776 35040
rect 29914 34960 29920 35012
rect 29972 35000 29978 35012
rect 30193 35003 30251 35009
rect 30193 35000 30205 35003
rect 29972 34972 30205 35000
rect 29972 34960 29978 34972
rect 30193 34969 30205 34972
rect 30239 34969 30251 35003
rect 30484 35000 30512 35099
rect 30558 35096 30564 35148
rect 30616 35136 30622 35148
rect 31113 35139 31171 35145
rect 31113 35136 31125 35139
rect 30616 35108 31125 35136
rect 30616 35096 30622 35108
rect 31113 35105 31125 35108
rect 31159 35105 31171 35139
rect 31113 35099 31171 35105
rect 30834 35028 30840 35080
rect 30892 35028 30898 35080
rect 31021 35003 31079 35009
rect 31021 35000 31033 35003
rect 30484 34972 31033 35000
rect 30193 34963 30251 34969
rect 31021 34969 31033 34972
rect 31067 34969 31079 35003
rect 31021 34963 31079 34969
rect 28684 34904 29776 34932
rect 28684 34892 28690 34904
rect 30282 34892 30288 34944
rect 30340 34932 30346 34944
rect 30745 34935 30803 34941
rect 30745 34932 30757 34935
rect 30340 34904 30757 34932
rect 30340 34892 30346 34904
rect 30745 34901 30757 34904
rect 30791 34901 30803 34935
rect 30745 34895 30803 34901
rect 552 34842 31648 34864
rect 552 34790 3662 34842
rect 3714 34790 3726 34842
rect 3778 34790 3790 34842
rect 3842 34790 3854 34842
rect 3906 34790 3918 34842
rect 3970 34790 11436 34842
rect 11488 34790 11500 34842
rect 11552 34790 11564 34842
rect 11616 34790 11628 34842
rect 11680 34790 11692 34842
rect 11744 34790 19210 34842
rect 19262 34790 19274 34842
rect 19326 34790 19338 34842
rect 19390 34790 19402 34842
rect 19454 34790 19466 34842
rect 19518 34790 26984 34842
rect 27036 34790 27048 34842
rect 27100 34790 27112 34842
rect 27164 34790 27176 34842
rect 27228 34790 27240 34842
rect 27292 34790 31648 34842
rect 552 34768 31648 34790
rect 9674 34688 9680 34740
rect 9732 34728 9738 34740
rect 9769 34731 9827 34737
rect 9769 34728 9781 34731
rect 9732 34700 9781 34728
rect 9732 34688 9738 34700
rect 9769 34697 9781 34700
rect 9815 34728 9827 34731
rect 10410 34728 10416 34740
rect 9815 34700 10416 34728
rect 9815 34697 9827 34700
rect 9769 34691 9827 34697
rect 10410 34688 10416 34700
rect 10468 34688 10474 34740
rect 11790 34688 11796 34740
rect 11848 34728 11854 34740
rect 12066 34728 12072 34740
rect 11848 34700 12072 34728
rect 11848 34688 11854 34700
rect 12066 34688 12072 34700
rect 12124 34688 12130 34740
rect 13357 34731 13415 34737
rect 13357 34697 13369 34731
rect 13403 34728 13415 34731
rect 14550 34728 14556 34740
rect 13403 34700 14556 34728
rect 13403 34697 13415 34700
rect 13357 34691 13415 34697
rect 14550 34688 14556 34700
rect 14608 34688 14614 34740
rect 14734 34688 14740 34740
rect 14792 34728 14798 34740
rect 16482 34728 16488 34740
rect 14792 34700 15148 34728
rect 14792 34688 14798 34700
rect 12434 34660 12440 34672
rect 10152 34632 12440 34660
rect 8113 34595 8171 34601
rect 8113 34561 8125 34595
rect 8159 34592 8171 34595
rect 8389 34595 8447 34601
rect 8389 34592 8401 34595
rect 8159 34564 8401 34592
rect 8159 34561 8171 34564
rect 8113 34555 8171 34561
rect 8389 34561 8401 34564
rect 8435 34561 8447 34595
rect 8389 34555 8447 34561
rect 8205 34527 8263 34533
rect 8205 34493 8217 34527
rect 8251 34524 8263 34527
rect 9122 34524 9128 34536
rect 8251 34496 9128 34524
rect 8251 34493 8263 34496
rect 8205 34487 8263 34493
rect 9122 34484 9128 34496
rect 9180 34524 9186 34536
rect 9180 34496 9674 34524
rect 9180 34484 9186 34496
rect 8656 34459 8714 34465
rect 8656 34425 8668 34459
rect 8702 34456 8714 34459
rect 8846 34456 8852 34468
rect 8702 34428 8852 34456
rect 8702 34425 8714 34428
rect 8656 34419 8714 34425
rect 8846 34416 8852 34428
rect 8904 34416 8910 34468
rect 9646 34456 9674 34496
rect 10042 34484 10048 34536
rect 10100 34484 10106 34536
rect 10152 34533 10180 34632
rect 12434 34620 12440 34632
rect 12492 34660 12498 34672
rect 13446 34660 13452 34672
rect 12492 34632 13452 34660
rect 12492 34620 12498 34632
rect 13446 34620 13452 34632
rect 13504 34620 13510 34672
rect 15013 34663 15071 34669
rect 15013 34629 15025 34663
rect 15059 34629 15071 34663
rect 15120 34660 15148 34700
rect 15396 34700 16488 34728
rect 15396 34660 15424 34700
rect 16316 34669 16344 34700
rect 16482 34688 16488 34700
rect 16540 34688 16546 34740
rect 19058 34728 19064 34740
rect 17696 34700 19064 34728
rect 15120 34632 15424 34660
rect 16301 34663 16359 34669
rect 15013 34623 15071 34629
rect 16301 34629 16313 34663
rect 16347 34629 16359 34663
rect 16301 34623 16359 34629
rect 12529 34595 12587 34601
rect 10244 34564 12480 34592
rect 10137 34527 10195 34533
rect 10137 34493 10149 34527
rect 10183 34493 10195 34527
rect 10137 34487 10195 34493
rect 10244 34456 10272 34564
rect 10321 34527 10379 34533
rect 10321 34493 10333 34527
rect 10367 34493 10379 34527
rect 10321 34487 10379 34493
rect 10413 34527 10471 34533
rect 10413 34493 10425 34527
rect 10459 34526 10471 34527
rect 10459 34524 10548 34526
rect 11054 34524 11060 34536
rect 10459 34498 11060 34524
rect 10459 34493 10471 34498
rect 10520 34496 11060 34498
rect 10413 34487 10471 34493
rect 9646 34428 10272 34456
rect 10348 34400 10376 34487
rect 11054 34484 11060 34496
rect 11112 34484 11118 34536
rect 12452 34533 12480 34564
rect 12529 34561 12541 34595
rect 12575 34592 12587 34595
rect 13633 34595 13691 34601
rect 13633 34592 13645 34595
rect 12575 34564 13645 34592
rect 12575 34561 12587 34564
rect 12529 34555 12587 34561
rect 13633 34561 13645 34564
rect 13679 34561 13691 34595
rect 13633 34555 13691 34561
rect 15028 34592 15056 34623
rect 15749 34595 15807 34601
rect 15749 34592 15761 34595
rect 15028 34564 15761 34592
rect 12437 34527 12495 34533
rect 12437 34493 12449 34527
rect 12483 34493 12495 34527
rect 12437 34487 12495 34493
rect 12713 34527 12771 34533
rect 12713 34493 12725 34527
rect 12759 34524 12771 34527
rect 12802 34524 12808 34536
rect 12759 34496 12808 34524
rect 12759 34493 12771 34496
rect 12713 34487 12771 34493
rect 12802 34484 12808 34496
rect 12860 34484 12866 34536
rect 12894 34484 12900 34536
rect 12952 34484 12958 34536
rect 12989 34527 13047 34533
rect 12989 34493 13001 34527
rect 13035 34493 13047 34527
rect 12989 34487 13047 34493
rect 13081 34527 13139 34533
rect 13081 34493 13093 34527
rect 13127 34524 13139 34527
rect 13262 34524 13268 34536
rect 13127 34496 13268 34524
rect 13127 34493 13139 34496
rect 13081 34487 13139 34493
rect 13004 34456 13032 34487
rect 13262 34484 13268 34496
rect 13320 34484 13326 34536
rect 13906 34533 13912 34536
rect 13900 34524 13912 34533
rect 13867 34496 13912 34524
rect 13900 34487 13912 34496
rect 13906 34484 13912 34487
rect 13964 34484 13970 34536
rect 13170 34456 13176 34468
rect 13004 34428 13176 34456
rect 13170 34416 13176 34428
rect 13228 34416 13234 34468
rect 13722 34416 13728 34468
rect 13780 34456 13786 34468
rect 15028 34456 15056 34564
rect 15749 34561 15761 34564
rect 15795 34561 15807 34595
rect 15749 34555 15807 34561
rect 15908 34595 15966 34601
rect 15908 34561 15920 34595
rect 15954 34592 15966 34595
rect 16666 34592 16672 34604
rect 15954 34564 16672 34592
rect 15954 34561 15966 34564
rect 15908 34555 15966 34561
rect 16666 34552 16672 34564
rect 16724 34552 16730 34604
rect 16945 34595 17003 34601
rect 16945 34561 16957 34595
rect 16991 34592 17003 34595
rect 17696 34592 17724 34700
rect 19058 34688 19064 34700
rect 19116 34688 19122 34740
rect 20714 34688 20720 34740
rect 20772 34688 20778 34740
rect 22094 34728 22100 34740
rect 21192 34700 22100 34728
rect 18417 34663 18475 34669
rect 18417 34629 18429 34663
rect 18463 34660 18475 34663
rect 18463 34632 19104 34660
rect 18463 34629 18475 34632
rect 18417 34623 18475 34629
rect 18046 34592 18052 34604
rect 16991 34564 17724 34592
rect 17788 34564 18052 34592
rect 16991 34561 17003 34564
rect 16945 34555 17003 34561
rect 15102 34484 15108 34536
rect 15160 34484 15166 34536
rect 16022 34484 16028 34536
rect 16080 34484 16086 34536
rect 16761 34527 16819 34533
rect 16761 34493 16773 34527
rect 16807 34524 16819 34527
rect 17788 34524 17816 34564
rect 18046 34552 18052 34564
rect 18104 34552 18110 34604
rect 18138 34552 18144 34604
rect 18196 34592 18202 34604
rect 18785 34595 18843 34601
rect 18785 34592 18797 34595
rect 18196 34564 18797 34592
rect 18196 34552 18202 34564
rect 18785 34561 18797 34564
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 18966 34552 18972 34604
rect 19024 34552 19030 34604
rect 19076 34601 19104 34632
rect 21192 34601 21220 34700
rect 22066 34688 22100 34700
rect 22152 34688 22158 34740
rect 22557 34731 22615 34737
rect 22557 34697 22569 34731
rect 22603 34728 22615 34731
rect 22922 34728 22928 34740
rect 22603 34700 22928 34728
rect 22603 34697 22615 34700
rect 22557 34691 22615 34697
rect 22922 34688 22928 34700
rect 22980 34688 22986 34740
rect 23934 34688 23940 34740
rect 23992 34688 23998 34740
rect 24121 34731 24179 34737
rect 24121 34697 24133 34731
rect 24167 34728 24179 34731
rect 25682 34728 25688 34740
rect 24167 34700 25688 34728
rect 24167 34697 24179 34700
rect 24121 34691 24179 34697
rect 25682 34688 25688 34700
rect 25740 34688 25746 34740
rect 26694 34688 26700 34740
rect 26752 34728 26758 34740
rect 28350 34728 28356 34740
rect 26752 34700 28356 34728
rect 26752 34688 26758 34700
rect 28350 34688 28356 34700
rect 28408 34728 28414 34740
rect 29638 34728 29644 34740
rect 28408 34700 29644 34728
rect 28408 34688 28414 34700
rect 29638 34688 29644 34700
rect 29696 34688 29702 34740
rect 29730 34688 29736 34740
rect 29788 34728 29794 34740
rect 30190 34728 30196 34740
rect 29788 34700 30196 34728
rect 29788 34688 29794 34700
rect 30190 34688 30196 34700
rect 30248 34728 30254 34740
rect 30377 34731 30435 34737
rect 30377 34728 30389 34731
rect 30248 34700 30389 34728
rect 30248 34688 30254 34700
rect 30377 34697 30389 34700
rect 30423 34697 30435 34731
rect 30377 34691 30435 34697
rect 30558 34688 30564 34740
rect 30616 34728 30622 34740
rect 30653 34731 30711 34737
rect 30653 34728 30665 34731
rect 30616 34700 30665 34728
rect 30616 34688 30622 34700
rect 30653 34697 30665 34700
rect 30699 34697 30711 34731
rect 30653 34691 30711 34697
rect 22066 34660 22094 34688
rect 22830 34660 22836 34672
rect 22066 34632 22836 34660
rect 22830 34620 22836 34632
rect 22888 34620 22894 34672
rect 24946 34620 24952 34672
rect 25004 34660 25010 34672
rect 25041 34663 25099 34669
rect 25041 34660 25053 34663
rect 25004 34632 25053 34660
rect 25004 34620 25010 34632
rect 25041 34629 25053 34632
rect 25087 34629 25099 34663
rect 25041 34623 25099 34629
rect 19061 34595 19119 34601
rect 19061 34561 19073 34595
rect 19107 34561 19119 34595
rect 21177 34595 21235 34601
rect 21177 34592 21189 34595
rect 19061 34555 19119 34561
rect 20824 34564 21189 34592
rect 16807 34496 17816 34524
rect 16807 34493 16819 34496
rect 16761 34487 16819 34493
rect 17954 34484 17960 34536
rect 18012 34524 18018 34536
rect 18325 34527 18383 34533
rect 18325 34524 18337 34527
rect 18012 34496 18337 34524
rect 18012 34484 18018 34496
rect 18325 34493 18337 34496
rect 18371 34493 18383 34527
rect 18325 34487 18383 34493
rect 18693 34527 18751 34533
rect 18693 34493 18705 34527
rect 18739 34524 18751 34527
rect 19317 34527 19375 34533
rect 19317 34524 19329 34527
rect 18739 34496 18920 34524
rect 18739 34493 18751 34496
rect 18693 34487 18751 34493
rect 13780 34428 15056 34456
rect 13780 34416 13786 34428
rect 9306 34348 9312 34400
rect 9364 34388 9370 34400
rect 9861 34391 9919 34397
rect 9861 34388 9873 34391
rect 9364 34360 9873 34388
rect 9364 34348 9370 34360
rect 9861 34357 9873 34360
rect 9907 34357 9919 34391
rect 9861 34351 9919 34357
rect 10318 34348 10324 34400
rect 10376 34348 10382 34400
rect 13906 34348 13912 34400
rect 13964 34388 13970 34400
rect 14182 34388 14188 34400
rect 13964 34360 14188 34388
rect 13964 34348 13970 34360
rect 14182 34348 14188 34360
rect 14240 34388 14246 34400
rect 18230 34388 18236 34400
rect 14240 34360 18236 34388
rect 14240 34348 14246 34360
rect 18230 34348 18236 34360
rect 18288 34348 18294 34400
rect 18892 34388 18920 34496
rect 18984 34496 19329 34524
rect 18984 34465 19012 34496
rect 19317 34493 19329 34496
rect 19363 34493 19375 34527
rect 19317 34487 19375 34493
rect 19610 34484 19616 34536
rect 19668 34524 19674 34536
rect 19886 34524 19892 34536
rect 19668 34496 19892 34524
rect 19668 34484 19674 34496
rect 19886 34484 19892 34496
rect 19944 34484 19950 34536
rect 20824 34533 20852 34564
rect 21177 34561 21189 34564
rect 21223 34561 21235 34595
rect 25406 34592 25412 34604
rect 21177 34555 21235 34561
rect 22296 34564 24164 34592
rect 20625 34527 20683 34533
rect 20625 34493 20637 34527
rect 20671 34493 20683 34527
rect 20625 34487 20683 34493
rect 20809 34527 20867 34533
rect 20809 34493 20821 34527
rect 20855 34493 20867 34527
rect 20809 34487 20867 34493
rect 20901 34527 20959 34533
rect 20901 34493 20913 34527
rect 20947 34524 20959 34527
rect 21082 34524 21088 34536
rect 20947 34496 21088 34524
rect 20947 34493 20959 34496
rect 20901 34487 20959 34493
rect 18969 34459 19027 34465
rect 18969 34425 18981 34459
rect 19015 34425 19027 34459
rect 18969 34419 19027 34425
rect 19518 34416 19524 34468
rect 19576 34456 19582 34468
rect 20640 34456 20668 34487
rect 21082 34484 21088 34496
rect 21140 34484 21146 34536
rect 22002 34484 22008 34536
rect 22060 34524 22066 34536
rect 22296 34533 22324 34564
rect 22097 34527 22155 34533
rect 22097 34524 22109 34527
rect 22060 34496 22109 34524
rect 22060 34484 22066 34496
rect 22097 34493 22109 34496
rect 22143 34493 22155 34527
rect 22097 34487 22155 34493
rect 22281 34527 22339 34533
rect 22281 34493 22293 34527
rect 22327 34493 22339 34527
rect 22281 34487 22339 34493
rect 22370 34484 22376 34536
rect 22428 34524 22434 34536
rect 23293 34527 23351 34533
rect 23293 34524 23305 34527
rect 22428 34496 23305 34524
rect 22428 34484 22434 34496
rect 23293 34493 23305 34496
rect 23339 34524 23351 34527
rect 23474 34524 23480 34536
rect 23339 34496 23480 34524
rect 23339 34493 23351 34496
rect 23293 34487 23351 34493
rect 23474 34484 23480 34496
rect 23532 34524 23538 34536
rect 23661 34527 23719 34533
rect 23661 34524 23673 34527
rect 23532 34496 23673 34524
rect 23532 34484 23538 34496
rect 23661 34493 23673 34496
rect 23707 34493 23719 34527
rect 23661 34487 23719 34493
rect 24136 34468 24164 34564
rect 24688 34564 25412 34592
rect 24688 34533 24716 34564
rect 25406 34552 25412 34564
rect 25464 34592 25470 34604
rect 25961 34595 26019 34601
rect 25961 34592 25973 34595
rect 25464 34564 25973 34592
rect 25464 34552 25470 34564
rect 25961 34561 25973 34564
rect 26007 34592 26019 34595
rect 26234 34592 26240 34604
rect 26007 34564 26240 34592
rect 26007 34561 26019 34564
rect 25961 34555 26019 34561
rect 26234 34552 26240 34564
rect 26292 34592 26298 34604
rect 26292 34564 27108 34592
rect 26292 34552 26298 34564
rect 24673 34527 24731 34533
rect 24673 34493 24685 34527
rect 24719 34493 24731 34527
rect 24673 34487 24731 34493
rect 24762 34484 24768 34536
rect 24820 34484 24826 34536
rect 25038 34484 25044 34536
rect 25096 34484 25102 34536
rect 26712 34533 26740 34564
rect 26697 34527 26755 34533
rect 26697 34493 26709 34527
rect 26743 34493 26755 34527
rect 26697 34487 26755 34493
rect 26789 34527 26847 34533
rect 26789 34493 26801 34527
rect 26835 34524 26847 34527
rect 26973 34527 27031 34533
rect 26973 34524 26985 34527
rect 26835 34496 26985 34524
rect 26835 34493 26847 34496
rect 26789 34487 26847 34493
rect 26973 34493 26985 34496
rect 27019 34493 27031 34527
rect 27080 34524 27108 34564
rect 28626 34524 28632 34536
rect 27080 34496 28632 34524
rect 26973 34487 27031 34493
rect 28626 34484 28632 34496
rect 28684 34484 28690 34536
rect 28721 34527 28779 34533
rect 28721 34493 28733 34527
rect 28767 34524 28779 34527
rect 28997 34527 29055 34533
rect 28997 34524 29009 34527
rect 28767 34496 29009 34524
rect 28767 34493 28779 34496
rect 28721 34487 28779 34493
rect 28997 34493 29009 34496
rect 29043 34493 29055 34527
rect 28997 34487 29055 34493
rect 31294 34484 31300 34536
rect 31352 34484 31358 34536
rect 19576 34428 21956 34456
rect 19576 34416 19582 34428
rect 19794 34388 19800 34400
rect 18892 34360 19800 34388
rect 19794 34348 19800 34360
rect 19852 34348 19858 34400
rect 20441 34391 20499 34397
rect 20441 34357 20453 34391
rect 20487 34388 20499 34391
rect 21082 34388 21088 34400
rect 20487 34360 21088 34388
rect 20487 34357 20499 34360
rect 20441 34351 20499 34357
rect 21082 34348 21088 34360
rect 21140 34348 21146 34400
rect 21928 34397 21956 34428
rect 22554 34416 22560 34468
rect 22612 34416 22618 34468
rect 24118 34416 24124 34468
rect 24176 34416 24182 34468
rect 24305 34459 24363 34465
rect 24305 34425 24317 34459
rect 24351 34456 24363 34459
rect 24486 34456 24492 34468
rect 24351 34428 24492 34456
rect 24351 34425 24363 34428
rect 24305 34419 24363 34425
rect 24486 34416 24492 34428
rect 24544 34416 24550 34468
rect 25130 34416 25136 34468
rect 25188 34416 25194 34468
rect 27240 34459 27298 34465
rect 27240 34425 27252 34459
rect 27286 34456 27298 34459
rect 27338 34456 27344 34468
rect 27286 34428 27344 34456
rect 27286 34425 27298 34428
rect 27240 34419 27298 34425
rect 27338 34416 27344 34428
rect 27396 34416 27402 34468
rect 29270 34465 29276 34468
rect 29264 34419 29276 34465
rect 29270 34416 29276 34419
rect 29328 34416 29334 34468
rect 21913 34391 21971 34397
rect 21913 34357 21925 34391
rect 21959 34357 21971 34391
rect 21913 34351 21971 34357
rect 22370 34348 22376 34400
rect 22428 34348 22434 34400
rect 23566 34348 23572 34400
rect 23624 34348 23630 34400
rect 24578 34348 24584 34400
rect 24636 34348 24642 34400
rect 24857 34391 24915 34397
rect 24857 34357 24869 34391
rect 24903 34388 24915 34391
rect 25590 34388 25596 34400
rect 24903 34360 25596 34388
rect 24903 34357 24915 34360
rect 24857 34351 24915 34357
rect 25590 34348 25596 34360
rect 25648 34348 25654 34400
rect 552 34298 31648 34320
rect 552 34246 4322 34298
rect 4374 34246 4386 34298
rect 4438 34246 4450 34298
rect 4502 34246 4514 34298
rect 4566 34246 4578 34298
rect 4630 34246 12096 34298
rect 12148 34246 12160 34298
rect 12212 34246 12224 34298
rect 12276 34246 12288 34298
rect 12340 34246 12352 34298
rect 12404 34246 19870 34298
rect 19922 34246 19934 34298
rect 19986 34246 19998 34298
rect 20050 34246 20062 34298
rect 20114 34246 20126 34298
rect 20178 34246 27644 34298
rect 27696 34246 27708 34298
rect 27760 34246 27772 34298
rect 27824 34246 27836 34298
rect 27888 34246 27900 34298
rect 27952 34246 31648 34298
rect 552 34224 31648 34246
rect 8846 34144 8852 34196
rect 8904 34144 8910 34196
rect 9490 34144 9496 34196
rect 9548 34184 9554 34196
rect 9585 34187 9643 34193
rect 9585 34184 9597 34187
rect 9548 34156 9597 34184
rect 9548 34144 9554 34156
rect 9585 34153 9597 34156
rect 9631 34153 9643 34187
rect 11330 34184 11336 34196
rect 9585 34147 9643 34153
rect 9876 34156 11336 34184
rect 9876 34116 9904 34156
rect 11330 34144 11336 34156
rect 11388 34184 11394 34196
rect 11790 34184 11796 34196
rect 11388 34156 11796 34184
rect 11388 34144 11394 34156
rect 11790 34144 11796 34156
rect 11848 34144 11854 34196
rect 12894 34144 12900 34196
rect 12952 34184 12958 34196
rect 12952 34156 13676 34184
rect 12952 34144 12958 34156
rect 9508 34088 9904 34116
rect 9953 34119 10011 34125
rect 9125 34051 9183 34057
rect 9125 34017 9137 34051
rect 9171 34017 9183 34051
rect 9125 34011 9183 34017
rect 9140 33980 9168 34011
rect 9214 34008 9220 34060
rect 9272 34008 9278 34060
rect 9306 34008 9312 34060
rect 9364 34008 9370 34060
rect 9508 34057 9536 34088
rect 9953 34085 9965 34119
rect 9999 34116 10011 34119
rect 10226 34116 10232 34128
rect 9999 34088 10232 34116
rect 9999 34085 10011 34088
rect 9953 34079 10011 34085
rect 10226 34076 10232 34088
rect 10284 34116 10290 34128
rect 11149 34119 11207 34125
rect 11149 34116 11161 34119
rect 10284 34088 11161 34116
rect 10284 34076 10290 34088
rect 11149 34085 11161 34088
rect 11195 34116 11207 34119
rect 12434 34116 12440 34128
rect 11195 34088 12440 34116
rect 11195 34085 11207 34088
rect 11149 34079 11207 34085
rect 12434 34076 12440 34088
rect 12492 34116 12498 34128
rect 13173 34119 13231 34125
rect 13173 34116 13185 34119
rect 12492 34088 13185 34116
rect 12492 34076 12498 34088
rect 13173 34085 13185 34088
rect 13219 34116 13231 34119
rect 13265 34119 13323 34125
rect 13265 34116 13277 34119
rect 13219 34088 13277 34116
rect 13219 34085 13231 34088
rect 13173 34079 13231 34085
rect 13265 34085 13277 34088
rect 13311 34116 13323 34119
rect 13538 34116 13544 34128
rect 13311 34088 13544 34116
rect 13311 34085 13323 34088
rect 13265 34079 13323 34085
rect 13538 34076 13544 34088
rect 13596 34076 13602 34128
rect 13648 34125 13676 34156
rect 14274 34144 14280 34196
rect 14332 34184 14338 34196
rect 14461 34187 14519 34193
rect 14461 34184 14473 34187
rect 14332 34156 14473 34184
rect 14332 34144 14338 34156
rect 14461 34153 14473 34156
rect 14507 34153 14519 34187
rect 14461 34147 14519 34153
rect 14936 34156 16712 34184
rect 13633 34119 13691 34125
rect 13633 34085 13645 34119
rect 13679 34116 13691 34119
rect 14936 34116 14964 34156
rect 13679 34088 14964 34116
rect 15381 34119 15439 34125
rect 13679 34085 13691 34088
rect 13633 34079 13691 34085
rect 15381 34085 15393 34119
rect 15427 34116 15439 34119
rect 15427 34088 15884 34116
rect 15427 34085 15439 34088
rect 15381 34079 15439 34085
rect 9493 34051 9551 34057
rect 9493 34017 9505 34051
rect 9539 34017 9551 34051
rect 9493 34011 9551 34017
rect 9766 34008 9772 34060
rect 9824 34008 9830 34060
rect 11333 34051 11391 34057
rect 11333 34017 11345 34051
rect 11379 34048 11391 34051
rect 11882 34048 11888 34060
rect 11379 34020 11888 34048
rect 11379 34017 11391 34020
rect 11333 34011 11391 34017
rect 11882 34008 11888 34020
rect 11940 34008 11946 34060
rect 12986 34008 12992 34060
rect 13044 34008 13050 34060
rect 13449 34051 13507 34057
rect 13449 34017 13461 34051
rect 13495 34048 13507 34051
rect 14093 34051 14151 34057
rect 14093 34048 14105 34051
rect 13495 34020 14105 34048
rect 13495 34017 13507 34020
rect 13449 34011 13507 34017
rect 13556 33992 13584 34020
rect 14093 34017 14105 34020
rect 14139 34048 14151 34051
rect 14734 34048 14740 34060
rect 14139 34020 14740 34048
rect 14139 34017 14151 34020
rect 14093 34011 14151 34017
rect 14734 34008 14740 34020
rect 14792 34008 14798 34060
rect 14829 34051 14887 34057
rect 14829 34017 14841 34051
rect 14875 34048 14887 34051
rect 14875 34020 14964 34048
rect 14875 34017 14887 34020
rect 14829 34011 14887 34017
rect 9674 33980 9680 33992
rect 9140 33952 9680 33980
rect 9674 33940 9680 33952
rect 9732 33940 9738 33992
rect 13538 33940 13544 33992
rect 13596 33940 13602 33992
rect 13906 33940 13912 33992
rect 13964 33940 13970 33992
rect 14001 33983 14059 33989
rect 14001 33949 14013 33983
rect 14047 33949 14059 33983
rect 14001 33943 14059 33949
rect 9306 33872 9312 33924
rect 9364 33912 9370 33924
rect 11238 33912 11244 33924
rect 9364 33884 11244 33912
rect 9364 33872 9370 33884
rect 11238 33872 11244 33884
rect 11296 33872 11302 33924
rect 12066 33872 12072 33924
rect 12124 33912 12130 33924
rect 12710 33912 12716 33924
rect 12124 33884 12716 33912
rect 12124 33872 12130 33884
rect 12710 33872 12716 33884
rect 12768 33912 12774 33924
rect 13262 33912 13268 33924
rect 12768 33884 13268 33912
rect 12768 33872 12774 33884
rect 13262 33872 13268 33884
rect 13320 33912 13326 33924
rect 14016 33912 14044 33943
rect 13320 33884 14044 33912
rect 13320 33872 13326 33884
rect 11517 33847 11575 33853
rect 11517 33813 11529 33847
rect 11563 33844 11575 33847
rect 11790 33844 11796 33856
rect 11563 33816 11796 33844
rect 11563 33813 11575 33816
rect 11517 33807 11575 33813
rect 11790 33804 11796 33816
rect 11848 33804 11854 33856
rect 12802 33804 12808 33856
rect 12860 33844 12866 33856
rect 14936 33853 14964 34020
rect 15470 34008 15476 34060
rect 15528 34008 15534 34060
rect 15562 34008 15568 34060
rect 15620 34048 15626 34060
rect 15856 34057 15884 34088
rect 15687 34051 15745 34057
rect 15687 34048 15699 34051
rect 15620 34020 15699 34048
rect 15620 34008 15626 34020
rect 15687 34017 15699 34020
rect 15733 34017 15745 34051
rect 15687 34011 15745 34017
rect 15841 34051 15899 34057
rect 15841 34017 15853 34051
rect 15887 34048 15899 34051
rect 16298 34048 16304 34060
rect 15887 34020 16304 34048
rect 15887 34017 15899 34020
rect 15841 34011 15899 34017
rect 16298 34008 16304 34020
rect 16356 34008 16362 34060
rect 16485 34051 16543 34057
rect 16485 34017 16497 34051
rect 16531 34017 16543 34051
rect 16485 34011 16543 34017
rect 15105 33915 15163 33921
rect 15105 33881 15117 33915
rect 15151 33912 15163 33915
rect 15580 33912 15608 34008
rect 15151 33884 15608 33912
rect 16500 33912 16528 34011
rect 16574 34008 16580 34060
rect 16632 34008 16638 34060
rect 16684 34048 16712 34156
rect 18138 34144 18144 34196
rect 18196 34144 18202 34196
rect 18230 34144 18236 34196
rect 18288 34144 18294 34196
rect 18966 34144 18972 34196
rect 19024 34184 19030 34196
rect 19245 34187 19303 34193
rect 19245 34184 19257 34187
rect 19024 34156 19257 34184
rect 19024 34144 19030 34156
rect 19245 34153 19257 34156
rect 19291 34153 19303 34187
rect 19245 34147 19303 34153
rect 21637 34187 21695 34193
rect 21637 34153 21649 34187
rect 21683 34184 21695 34187
rect 22278 34184 22284 34196
rect 21683 34156 22284 34184
rect 21683 34153 21695 34156
rect 21637 34147 21695 34153
rect 22278 34144 22284 34156
rect 22336 34144 22342 34196
rect 25130 34184 25136 34196
rect 22388 34156 25136 34184
rect 16758 34076 16764 34128
rect 16816 34116 16822 34128
rect 16853 34119 16911 34125
rect 16853 34116 16865 34119
rect 16816 34088 16865 34116
rect 16816 34076 16822 34088
rect 16853 34085 16865 34088
rect 16899 34116 16911 34119
rect 22094 34116 22100 34128
rect 16899 34088 22100 34116
rect 16899 34085 16911 34088
rect 16853 34079 16911 34085
rect 22094 34076 22100 34088
rect 22152 34116 22158 34128
rect 22388 34116 22416 34156
rect 25130 34144 25136 34156
rect 25188 34144 25194 34196
rect 29181 34187 29239 34193
rect 29181 34153 29193 34187
rect 29227 34184 29239 34187
rect 29270 34184 29276 34196
rect 29227 34156 29276 34184
rect 29227 34153 29239 34156
rect 29181 34147 29239 34153
rect 29270 34144 29276 34156
rect 29328 34144 29334 34196
rect 31294 34144 31300 34196
rect 31352 34144 31358 34196
rect 23566 34116 23572 34128
rect 22152 34088 22416 34116
rect 22480 34088 23572 34116
rect 22152 34076 22158 34088
rect 18325 34051 18383 34057
rect 18325 34048 18337 34051
rect 16684 34020 18337 34048
rect 18325 34017 18337 34020
rect 18371 34017 18383 34051
rect 18325 34011 18383 34017
rect 18417 34051 18475 34057
rect 18417 34017 18429 34051
rect 18463 34017 18475 34051
rect 18417 34011 18475 34017
rect 16592 33980 16620 34008
rect 17589 33983 17647 33989
rect 17589 33980 17601 33983
rect 16592 33952 17601 33980
rect 17589 33949 17601 33952
rect 17635 33980 17647 33983
rect 17954 33980 17960 33992
rect 17635 33952 17960 33980
rect 17635 33949 17647 33952
rect 17589 33943 17647 33949
rect 17954 33940 17960 33952
rect 18012 33940 18018 33992
rect 18046 33940 18052 33992
rect 18104 33980 18110 33992
rect 18432 33980 18460 34011
rect 18506 34008 18512 34060
rect 18564 34008 18570 34060
rect 18874 34008 18880 34060
rect 18932 34008 18938 34060
rect 19061 34051 19119 34057
rect 19061 34017 19073 34051
rect 19107 34048 19119 34051
rect 19150 34048 19156 34060
rect 19107 34020 19156 34048
rect 19107 34017 19119 34020
rect 19061 34011 19119 34017
rect 19150 34008 19156 34020
rect 19208 34008 19214 34060
rect 19521 34051 19579 34057
rect 19521 34017 19533 34051
rect 19567 34048 19579 34051
rect 19610 34048 19616 34060
rect 19567 34020 19616 34048
rect 19567 34017 19579 34020
rect 19521 34011 19579 34017
rect 19610 34008 19616 34020
rect 19668 34008 19674 34060
rect 19702 34008 19708 34060
rect 19760 34008 19766 34060
rect 19794 34008 19800 34060
rect 19852 34008 19858 34060
rect 22480 34057 22508 34088
rect 23566 34076 23572 34088
rect 23624 34076 23630 34128
rect 26418 34076 26424 34128
rect 26476 34116 26482 34128
rect 26786 34116 26792 34128
rect 26476 34088 26792 34116
rect 26476 34076 26482 34088
rect 26786 34076 26792 34088
rect 26844 34116 26850 34128
rect 27338 34116 27344 34128
rect 26844 34088 27344 34116
rect 26844 34076 26850 34088
rect 27338 34076 27344 34088
rect 27396 34076 27402 34128
rect 27709 34119 27767 34125
rect 27709 34085 27721 34119
rect 27755 34116 27767 34119
rect 27982 34116 27988 34128
rect 27755 34088 27988 34116
rect 27755 34085 27767 34088
rect 27709 34079 27767 34085
rect 27982 34076 27988 34088
rect 28040 34076 28046 34128
rect 28997 34119 29055 34125
rect 28997 34085 29009 34119
rect 29043 34116 29055 34119
rect 29638 34116 29644 34128
rect 29043 34088 29316 34116
rect 29043 34085 29055 34088
rect 28997 34079 29055 34085
rect 22465 34051 22523 34057
rect 22465 34017 22477 34051
rect 22511 34017 22523 34051
rect 22465 34011 22523 34017
rect 22554 34008 22560 34060
rect 22612 34048 22618 34060
rect 22721 34051 22779 34057
rect 22721 34048 22733 34051
rect 22612 34020 22733 34048
rect 22612 34008 22618 34020
rect 22721 34017 22733 34020
rect 22767 34017 22779 34051
rect 22721 34011 22779 34017
rect 24578 34008 24584 34060
rect 24636 34008 24642 34060
rect 24854 34057 24860 34060
rect 24848 34011 24860 34057
rect 24854 34008 24860 34011
rect 24912 34008 24918 34060
rect 26234 34008 26240 34060
rect 26292 34008 26298 34060
rect 27157 34051 27215 34057
rect 27157 34048 27169 34051
rect 26344 34020 27169 34048
rect 18969 33983 19027 33989
rect 18969 33980 18981 33983
rect 18104 33952 18368 33980
rect 18432 33952 18981 33980
rect 18104 33940 18110 33952
rect 16942 33912 16948 33924
rect 16500 33884 16948 33912
rect 15151 33881 15163 33884
rect 15105 33875 15163 33881
rect 16942 33872 16948 33884
rect 17000 33872 17006 33924
rect 18340 33912 18368 33952
rect 18892 33924 18920 33952
rect 18969 33949 18981 33952
rect 19015 33949 19027 33983
rect 19720 33980 19748 34008
rect 18969 33943 19027 33949
rect 19628 33952 19748 33980
rect 18340 33884 18828 33912
rect 18800 33856 18828 33884
rect 18874 33872 18880 33924
rect 18932 33872 18938 33924
rect 19628 33856 19656 33952
rect 21726 33940 21732 33992
rect 21784 33940 21790 33992
rect 21818 33940 21824 33992
rect 21876 33940 21882 33992
rect 25682 33940 25688 33992
rect 25740 33980 25746 33992
rect 26344 33980 26372 34020
rect 27157 34017 27169 34020
rect 27203 34017 27215 34051
rect 27157 34011 27215 34017
rect 28629 34051 28687 34057
rect 28629 34017 28641 34051
rect 28675 34048 28687 34051
rect 29178 34048 29184 34060
rect 28675 34020 29184 34048
rect 28675 34017 28687 34020
rect 28629 34011 28687 34017
rect 29178 34008 29184 34020
rect 29236 34008 29242 34060
rect 29288 33989 29316 34088
rect 29472 34088 29644 34116
rect 29472 34057 29500 34088
rect 29638 34076 29644 34088
rect 29696 34076 29702 34128
rect 30184 34119 30242 34125
rect 30184 34085 30196 34119
rect 30230 34116 30242 34119
rect 30282 34116 30288 34128
rect 30230 34088 30288 34116
rect 30230 34085 30242 34088
rect 30184 34079 30242 34085
rect 30282 34076 30288 34088
rect 30340 34076 30346 34128
rect 29457 34051 29515 34057
rect 29457 34017 29469 34051
rect 29503 34017 29515 34051
rect 29457 34011 29515 34017
rect 29730 34008 29736 34060
rect 29788 34008 29794 34060
rect 29914 34008 29920 34060
rect 29972 34008 29978 34060
rect 25740 33952 26372 33980
rect 26973 33983 27031 33989
rect 25740 33940 25746 33952
rect 26973 33949 26985 33983
rect 27019 33949 27031 33983
rect 26973 33943 27031 33949
rect 29273 33983 29331 33989
rect 29273 33949 29285 33983
rect 29319 33949 29331 33983
rect 29273 33943 29331 33949
rect 25590 33872 25596 33924
rect 25648 33912 25654 33924
rect 25961 33915 26019 33921
rect 25961 33912 25973 33915
rect 25648 33884 25973 33912
rect 25648 33872 25654 33884
rect 25961 33881 25973 33884
rect 26007 33912 26019 33915
rect 26510 33912 26516 33924
rect 26007 33884 26516 33912
rect 26007 33881 26019 33884
rect 25961 33875 26019 33881
rect 26510 33872 26516 33884
rect 26568 33912 26574 33924
rect 26988 33912 27016 33943
rect 29546 33940 29552 33992
rect 29604 33940 29610 33992
rect 29641 33983 29699 33989
rect 29641 33949 29653 33983
rect 29687 33949 29699 33983
rect 29641 33943 29699 33949
rect 26568 33884 27016 33912
rect 27893 33915 27951 33921
rect 26568 33872 26574 33884
rect 27893 33881 27905 33915
rect 27939 33912 27951 33915
rect 27982 33912 27988 33924
rect 27939 33884 27988 33912
rect 27939 33881 27951 33884
rect 27893 33875 27951 33881
rect 27982 33872 27988 33884
rect 28040 33872 28046 33924
rect 28902 33872 28908 33924
rect 28960 33912 28966 33924
rect 29656 33912 29684 33943
rect 28960 33884 29684 33912
rect 28960 33872 28966 33884
rect 14645 33847 14703 33853
rect 14645 33844 14657 33847
rect 12860 33816 14657 33844
rect 12860 33804 12866 33816
rect 14645 33813 14657 33816
rect 14691 33813 14703 33847
rect 14645 33807 14703 33813
rect 14921 33847 14979 33853
rect 14921 33813 14933 33847
rect 14967 33844 14979 33847
rect 15378 33844 15384 33856
rect 14967 33816 15384 33844
rect 14967 33813 14979 33816
rect 14921 33807 14979 33813
rect 15378 33804 15384 33816
rect 15436 33804 15442 33856
rect 16114 33804 16120 33856
rect 16172 33844 16178 33856
rect 16301 33847 16359 33853
rect 16301 33844 16313 33847
rect 16172 33816 16313 33844
rect 16172 33804 16178 33816
rect 16301 33813 16313 33816
rect 16347 33813 16359 33847
rect 16301 33807 16359 33813
rect 16669 33847 16727 33853
rect 16669 33813 16681 33847
rect 16715 33844 16727 33847
rect 16850 33844 16856 33856
rect 16715 33816 16856 33844
rect 16715 33813 16727 33816
rect 16669 33807 16727 33813
rect 16850 33804 16856 33816
rect 16908 33804 16914 33856
rect 18598 33804 18604 33856
rect 18656 33844 18662 33856
rect 18693 33847 18751 33853
rect 18693 33844 18705 33847
rect 18656 33816 18705 33844
rect 18656 33804 18662 33816
rect 18693 33813 18705 33816
rect 18739 33813 18751 33847
rect 18693 33807 18751 33813
rect 18782 33804 18788 33856
rect 18840 33844 18846 33856
rect 19518 33844 19524 33856
rect 18840 33816 19524 33844
rect 18840 33804 18846 33816
rect 19518 33804 19524 33816
rect 19576 33804 19582 33856
rect 19610 33804 19616 33856
rect 19668 33804 19674 33856
rect 19705 33847 19763 33853
rect 19705 33813 19717 33847
rect 19751 33844 19763 33847
rect 20714 33844 20720 33856
rect 19751 33816 20720 33844
rect 19751 33813 19763 33816
rect 19705 33807 19763 33813
rect 20714 33804 20720 33816
rect 20772 33804 20778 33856
rect 21266 33804 21272 33856
rect 21324 33804 21330 33856
rect 22278 33804 22284 33856
rect 22336 33844 22342 33856
rect 23106 33844 23112 33856
rect 22336 33816 23112 33844
rect 22336 33804 22342 33816
rect 23106 33804 23112 33816
rect 23164 33804 23170 33856
rect 23845 33847 23903 33853
rect 23845 33813 23857 33847
rect 23891 33844 23903 33847
rect 24394 33844 24400 33856
rect 23891 33816 24400 33844
rect 23891 33813 23903 33816
rect 23845 33807 23903 33813
rect 24394 33804 24400 33816
rect 24452 33804 24458 33856
rect 26142 33804 26148 33856
rect 26200 33804 26206 33856
rect 26326 33804 26332 33856
rect 26384 33844 26390 33856
rect 26421 33847 26479 33853
rect 26421 33844 26433 33847
rect 26384 33816 26433 33844
rect 26384 33804 26390 33816
rect 26421 33813 26433 33816
rect 26467 33813 26479 33847
rect 26421 33807 26479 33813
rect 27522 33804 27528 33856
rect 27580 33804 27586 33856
rect 28442 33804 28448 33856
rect 28500 33844 28506 33856
rect 28997 33847 29055 33853
rect 28997 33844 29009 33847
rect 28500 33816 29009 33844
rect 28500 33804 28506 33816
rect 28997 33813 29009 33816
rect 29043 33813 29055 33847
rect 28997 33807 29055 33813
rect 552 33754 31648 33776
rect 552 33702 3662 33754
rect 3714 33702 3726 33754
rect 3778 33702 3790 33754
rect 3842 33702 3854 33754
rect 3906 33702 3918 33754
rect 3970 33702 11436 33754
rect 11488 33702 11500 33754
rect 11552 33702 11564 33754
rect 11616 33702 11628 33754
rect 11680 33702 11692 33754
rect 11744 33702 19210 33754
rect 19262 33702 19274 33754
rect 19326 33702 19338 33754
rect 19390 33702 19402 33754
rect 19454 33702 19466 33754
rect 19518 33702 26984 33754
rect 27036 33702 27048 33754
rect 27100 33702 27112 33754
rect 27164 33702 27176 33754
rect 27228 33702 27240 33754
rect 27292 33702 31648 33754
rect 552 33680 31648 33702
rect 13630 33600 13636 33652
rect 13688 33640 13694 33652
rect 13817 33643 13875 33649
rect 13817 33640 13829 33643
rect 13688 33612 13829 33640
rect 13688 33600 13694 33612
rect 13817 33609 13829 33612
rect 13863 33609 13875 33643
rect 13817 33603 13875 33609
rect 16117 33643 16175 33649
rect 16117 33609 16129 33643
rect 16163 33640 16175 33643
rect 17126 33640 17132 33652
rect 16163 33612 17132 33640
rect 16163 33609 16175 33612
rect 16117 33603 16175 33609
rect 17126 33600 17132 33612
rect 17184 33600 17190 33652
rect 18874 33600 18880 33652
rect 18932 33600 18938 33652
rect 21726 33600 21732 33652
rect 21784 33600 21790 33652
rect 23842 33600 23848 33652
rect 23900 33600 23906 33652
rect 26142 33640 26148 33652
rect 25976 33612 26148 33640
rect 10502 33532 10508 33584
rect 10560 33572 10566 33584
rect 12342 33572 12348 33584
rect 10560 33544 10824 33572
rect 10560 33532 10566 33544
rect 9858 33464 9864 33516
rect 9916 33504 9922 33516
rect 10410 33504 10416 33516
rect 9916 33476 10416 33504
rect 9916 33464 9922 33476
rect 10410 33464 10416 33476
rect 10468 33504 10474 33516
rect 10796 33504 10824 33544
rect 11532 33544 12348 33572
rect 11532 33504 11560 33544
rect 12342 33532 12348 33544
rect 12400 33572 12406 33584
rect 12802 33572 12808 33584
rect 12400 33544 12808 33572
rect 12400 33532 12406 33544
rect 12802 33532 12808 33544
rect 12860 33532 12866 33584
rect 15562 33532 15568 33584
rect 15620 33572 15626 33584
rect 16758 33572 16764 33584
rect 15620 33544 16764 33572
rect 15620 33532 15626 33544
rect 16758 33532 16764 33544
rect 16816 33532 16822 33584
rect 18785 33575 18843 33581
rect 18785 33541 18797 33575
rect 18831 33572 18843 33575
rect 19058 33572 19064 33584
rect 18831 33544 19064 33572
rect 18831 33541 18843 33544
rect 18785 33535 18843 33541
rect 19058 33532 19064 33544
rect 19116 33532 19122 33584
rect 21637 33575 21695 33581
rect 21637 33541 21649 33575
rect 21683 33572 21695 33575
rect 22370 33572 22376 33584
rect 21683 33544 22376 33572
rect 21683 33541 21695 33544
rect 21637 33535 21695 33541
rect 22370 33532 22376 33544
rect 22428 33532 22434 33584
rect 10468 33476 10640 33504
rect 10468 33464 10474 33476
rect 9217 33439 9275 33445
rect 9217 33405 9229 33439
rect 9263 33436 9275 33439
rect 10226 33436 10232 33448
rect 9263 33408 10232 33436
rect 9263 33405 9275 33408
rect 9217 33399 9275 33405
rect 10226 33396 10232 33408
rect 10284 33396 10290 33448
rect 10612 33445 10640 33476
rect 10796 33476 11560 33504
rect 10796 33445 10824 33476
rect 10597 33439 10655 33445
rect 10597 33405 10609 33439
rect 10643 33405 10655 33439
rect 10597 33399 10655 33405
rect 10689 33439 10747 33445
rect 10689 33405 10701 33439
rect 10735 33405 10747 33439
rect 10689 33399 10747 33405
rect 10781 33439 10839 33445
rect 10781 33405 10793 33439
rect 10827 33405 10839 33439
rect 10781 33399 10839 33405
rect 9401 33371 9459 33377
rect 9401 33337 9413 33371
rect 9447 33368 9459 33371
rect 9858 33368 9864 33380
rect 9447 33340 9864 33368
rect 9447 33337 9459 33340
rect 9401 33331 9459 33337
rect 9858 33328 9864 33340
rect 9916 33328 9922 33380
rect 10042 33328 10048 33380
rect 10100 33368 10106 33380
rect 10704 33368 10732 33399
rect 10962 33396 10968 33448
rect 11020 33396 11026 33448
rect 11330 33396 11336 33448
rect 11388 33396 11394 33448
rect 11532 33445 11560 33476
rect 11790 33464 11796 33516
rect 11848 33464 11854 33516
rect 15286 33464 15292 33516
rect 15344 33504 15350 33516
rect 15344 33476 16528 33504
rect 15344 33464 15350 33476
rect 11425 33439 11483 33445
rect 11425 33405 11437 33439
rect 11471 33405 11483 33439
rect 11425 33399 11483 33405
rect 11517 33439 11575 33445
rect 11517 33405 11529 33439
rect 11563 33405 11575 33439
rect 11517 33399 11575 33405
rect 11701 33439 11759 33445
rect 11701 33405 11713 33439
rect 11747 33436 11759 33439
rect 11808 33436 11836 33464
rect 11747 33408 11836 33436
rect 11977 33439 12035 33445
rect 11747 33405 11759 33408
rect 11701 33399 11759 33405
rect 11977 33405 11989 33439
rect 12023 33436 12035 33439
rect 12066 33436 12072 33448
rect 12023 33408 12072 33436
rect 12023 33405 12035 33408
rect 11977 33399 12035 33405
rect 11440 33368 11468 33399
rect 12066 33396 12072 33408
rect 12124 33396 12130 33448
rect 12161 33439 12219 33445
rect 12161 33405 12173 33439
rect 12207 33436 12219 33439
rect 12253 33439 12311 33445
rect 12253 33436 12265 33439
rect 12207 33408 12265 33436
rect 12207 33405 12219 33408
rect 12161 33399 12219 33405
rect 12253 33405 12265 33408
rect 12299 33405 12311 33439
rect 12253 33399 12311 33405
rect 12342 33396 12348 33448
rect 12400 33433 12406 33448
rect 12437 33436 12495 33442
rect 12437 33433 12449 33436
rect 12400 33405 12449 33433
rect 12400 33396 12406 33405
rect 12437 33402 12449 33405
rect 12483 33402 12495 33436
rect 12437 33396 12495 33402
rect 12526 33396 12532 33448
rect 12584 33396 12590 33448
rect 12618 33396 12624 33448
rect 12676 33396 12682 33448
rect 13998 33396 14004 33448
rect 14056 33396 14062 33448
rect 14182 33396 14188 33448
rect 14240 33396 14246 33448
rect 16500 33445 16528 33476
rect 16850 33464 16856 33516
rect 16908 33464 16914 33516
rect 18506 33464 18512 33516
rect 18564 33504 18570 33516
rect 19610 33504 19616 33516
rect 18564 33476 19616 33504
rect 18564 33464 18570 33476
rect 19610 33464 19616 33476
rect 19668 33464 19674 33516
rect 20073 33507 20131 33513
rect 20073 33473 20085 33507
rect 20119 33504 20131 33507
rect 20257 33507 20315 33513
rect 20257 33504 20269 33507
rect 20119 33476 20269 33504
rect 20119 33473 20131 33476
rect 20073 33467 20131 33473
rect 20257 33473 20269 33476
rect 20303 33473 20315 33507
rect 24762 33504 24768 33516
rect 20257 33467 20315 33473
rect 24136 33476 24768 33504
rect 16393 33439 16451 33445
rect 16393 33405 16405 33439
rect 16439 33405 16451 33439
rect 16393 33399 16451 33405
rect 16485 33439 16543 33445
rect 16485 33405 16497 33439
rect 16531 33405 16543 33439
rect 16485 33399 16543 33405
rect 16577 33439 16635 33445
rect 16577 33405 16589 33439
rect 16623 33436 16635 33439
rect 16666 33436 16672 33448
rect 16623 33408 16672 33436
rect 16623 33405 16635 33408
rect 16577 33399 16635 33405
rect 11606 33368 11612 33380
rect 10100 33340 11612 33368
rect 10100 33328 10106 33340
rect 11606 33328 11612 33340
rect 11664 33328 11670 33380
rect 11793 33371 11851 33377
rect 11793 33337 11805 33371
rect 11839 33337 11851 33371
rect 11793 33331 11851 33337
rect 9585 33303 9643 33309
rect 9585 33269 9597 33303
rect 9631 33300 9643 33303
rect 9950 33300 9956 33312
rect 9631 33272 9956 33300
rect 9631 33269 9643 33272
rect 9585 33263 9643 33269
rect 9950 33260 9956 33272
rect 10008 33260 10014 33312
rect 10321 33303 10379 33309
rect 10321 33269 10333 33303
rect 10367 33300 10379 33303
rect 10686 33300 10692 33312
rect 10367 33272 10692 33300
rect 10367 33269 10379 33272
rect 10321 33263 10379 33269
rect 10686 33260 10692 33272
rect 10744 33260 10750 33312
rect 11054 33260 11060 33312
rect 11112 33260 11118 33312
rect 11808 33300 11836 33331
rect 12434 33300 12440 33312
rect 11808 33272 12440 33300
rect 12434 33260 12440 33272
rect 12492 33260 12498 33312
rect 12897 33303 12955 33309
rect 12897 33269 12909 33303
rect 12943 33300 12955 33303
rect 13630 33300 13636 33312
rect 12943 33272 13636 33300
rect 12943 33269 12955 33272
rect 12897 33263 12955 33269
rect 13630 33260 13636 33272
rect 13688 33260 13694 33312
rect 16408 33300 16436 33399
rect 16666 33396 16672 33408
rect 16724 33396 16730 33448
rect 16761 33439 16819 33445
rect 16761 33405 16773 33439
rect 16807 33436 16819 33439
rect 18046 33436 18052 33448
rect 16807 33408 18052 33436
rect 16807 33405 16819 33408
rect 16761 33399 16819 33405
rect 18046 33396 18052 33408
rect 18104 33396 18110 33448
rect 18138 33396 18144 33448
rect 18196 33436 18202 33448
rect 18693 33439 18751 33445
rect 18693 33436 18705 33439
rect 18196 33408 18705 33436
rect 18196 33396 18202 33408
rect 18693 33405 18705 33408
rect 18739 33405 18751 33439
rect 18693 33399 18751 33405
rect 18966 33396 18972 33448
rect 19024 33436 19030 33448
rect 20165 33439 20223 33445
rect 19024 33408 19196 33436
rect 19024 33396 19030 33408
rect 17126 33377 17132 33380
rect 17120 33368 17132 33377
rect 17087 33340 17132 33368
rect 17120 33331 17132 33340
rect 17126 33328 17132 33331
rect 17184 33328 17190 33380
rect 19058 33328 19064 33380
rect 19116 33328 19122 33380
rect 18138 33300 18144 33312
rect 16408 33272 18144 33300
rect 18138 33260 18144 33272
rect 18196 33260 18202 33312
rect 18233 33303 18291 33309
rect 18233 33269 18245 33303
rect 18279 33300 18291 33303
rect 18506 33300 18512 33312
rect 18279 33272 18512 33300
rect 18279 33269 18291 33272
rect 18233 33263 18291 33269
rect 18506 33260 18512 33272
rect 18564 33260 18570 33312
rect 18966 33260 18972 33312
rect 19024 33260 19030 33312
rect 19168 33300 19196 33408
rect 20165 33405 20177 33439
rect 20211 33436 20223 33439
rect 21726 33436 21732 33448
rect 20211 33408 21732 33436
rect 20211 33405 20223 33408
rect 20165 33399 20223 33405
rect 21726 33396 21732 33408
rect 21784 33396 21790 33448
rect 22370 33396 22376 33448
rect 22428 33436 22434 33448
rect 22428 33408 23152 33436
rect 22428 33396 22434 33408
rect 20524 33371 20582 33377
rect 20524 33337 20536 33371
rect 20570 33368 20582 33371
rect 21266 33368 21272 33380
rect 20570 33340 21272 33368
rect 20570 33337 20582 33340
rect 20524 33331 20582 33337
rect 21266 33328 21272 33340
rect 21324 33328 21330 33380
rect 22094 33328 22100 33380
rect 22152 33368 22158 33380
rect 22649 33371 22707 33377
rect 22649 33368 22661 33371
rect 22152 33340 22661 33368
rect 22152 33328 22158 33340
rect 22649 33337 22661 33340
rect 22695 33337 22707 33371
rect 23124 33368 23152 33408
rect 23474 33396 23480 33448
rect 23532 33396 23538 33448
rect 24136 33445 24164 33476
rect 24762 33464 24768 33476
rect 24820 33504 24826 33516
rect 25130 33504 25136 33516
rect 24820 33476 25136 33504
rect 24820 33464 24826 33476
rect 25130 33464 25136 33476
rect 25188 33464 25194 33516
rect 25976 33513 26004 33612
rect 26142 33600 26148 33612
rect 26200 33600 26206 33652
rect 27338 33600 27344 33652
rect 27396 33600 27402 33652
rect 28350 33532 28356 33584
rect 28408 33532 28414 33584
rect 25961 33507 26019 33513
rect 25961 33473 25973 33507
rect 26007 33473 26019 33507
rect 25961 33467 26019 33473
rect 28442 33464 28448 33516
rect 28500 33464 28506 33516
rect 29546 33504 29552 33516
rect 28644 33476 29552 33504
rect 24121 33439 24179 33445
rect 24121 33405 24133 33439
rect 24167 33405 24179 33439
rect 24121 33399 24179 33405
rect 24210 33396 24216 33448
rect 24268 33396 24274 33448
rect 24302 33396 24308 33448
rect 24360 33396 24366 33448
rect 24394 33396 24400 33448
rect 24452 33396 24458 33448
rect 24486 33396 24492 33448
rect 24544 33436 24550 33448
rect 24581 33439 24639 33445
rect 24581 33436 24593 33439
rect 24544 33408 24593 33436
rect 24544 33396 24550 33408
rect 24581 33405 24593 33408
rect 24627 33405 24639 33439
rect 24581 33399 24639 33405
rect 25777 33439 25835 33445
rect 25777 33405 25789 33439
rect 25823 33436 25835 33439
rect 26050 33436 26056 33448
rect 25823 33408 26056 33436
rect 25823 33405 25835 33408
rect 25777 33399 25835 33405
rect 26050 33396 26056 33408
rect 26108 33396 26114 33448
rect 28074 33396 28080 33448
rect 28132 33436 28138 33448
rect 28644 33445 28672 33476
rect 29546 33464 29552 33476
rect 29604 33464 29610 33516
rect 28629 33439 28687 33445
rect 28629 33436 28641 33439
rect 28132 33408 28641 33436
rect 28132 33396 28138 33408
rect 28629 33405 28641 33408
rect 28675 33405 28687 33439
rect 28629 33399 28687 33405
rect 28721 33439 28779 33445
rect 28721 33405 28733 33439
rect 28767 33436 28779 33439
rect 28902 33436 28908 33448
rect 28767 33408 28908 33436
rect 28767 33405 28779 33408
rect 28721 33399 28779 33405
rect 28902 33396 28908 33408
rect 28960 33396 28966 33448
rect 24504 33368 24532 33396
rect 23124 33340 24532 33368
rect 26228 33371 26286 33377
rect 22649 33331 22707 33337
rect 26228 33337 26240 33371
rect 26274 33368 26286 33371
rect 26418 33368 26424 33380
rect 26274 33340 26424 33368
rect 26274 33337 26286 33340
rect 26228 33331 26286 33337
rect 26418 33328 26424 33340
rect 26476 33328 26482 33380
rect 28353 33371 28411 33377
rect 28353 33337 28365 33371
rect 28399 33368 28411 33371
rect 28445 33371 28503 33377
rect 28445 33368 28457 33371
rect 28399 33340 28457 33368
rect 28399 33337 28411 33340
rect 28353 33331 28411 33337
rect 28445 33337 28457 33340
rect 28491 33337 28503 33371
rect 28445 33331 28503 33337
rect 20806 33300 20812 33312
rect 19168 33272 20812 33300
rect 20806 33260 20812 33272
rect 20864 33260 20870 33312
rect 28169 33303 28227 33309
rect 28169 33269 28181 33303
rect 28215 33300 28227 33303
rect 29086 33300 29092 33312
rect 28215 33272 29092 33300
rect 28215 33269 28227 33272
rect 28169 33263 28227 33269
rect 29086 33260 29092 33272
rect 29144 33260 29150 33312
rect 552 33210 31648 33232
rect 552 33158 4322 33210
rect 4374 33158 4386 33210
rect 4438 33158 4450 33210
rect 4502 33158 4514 33210
rect 4566 33158 4578 33210
rect 4630 33158 12096 33210
rect 12148 33158 12160 33210
rect 12212 33158 12224 33210
rect 12276 33158 12288 33210
rect 12340 33158 12352 33210
rect 12404 33158 19870 33210
rect 19922 33158 19934 33210
rect 19986 33158 19998 33210
rect 20050 33158 20062 33210
rect 20114 33158 20126 33210
rect 20178 33158 27644 33210
rect 27696 33158 27708 33210
rect 27760 33158 27772 33210
rect 27824 33158 27836 33210
rect 27888 33158 27900 33210
rect 27952 33158 31648 33210
rect 552 33136 31648 33158
rect 10410 33056 10416 33108
rect 10468 33056 10474 33108
rect 13081 33099 13139 33105
rect 13081 33065 13093 33099
rect 13127 33065 13139 33099
rect 13081 33059 13139 33065
rect 9309 33031 9367 33037
rect 9309 33028 9321 33031
rect 9140 33000 9321 33028
rect 8846 32920 8852 32972
rect 8904 32920 8910 32972
rect 9140 32969 9168 33000
rect 9309 32997 9321 33000
rect 9355 32997 9367 33031
rect 10042 33028 10048 33040
rect 9309 32991 9367 32997
rect 9692 33000 10048 33028
rect 8941 32963 8999 32969
rect 8941 32929 8953 32963
rect 8987 32929 8999 32963
rect 8941 32923 8999 32929
rect 9125 32963 9183 32969
rect 9125 32929 9137 32963
rect 9171 32929 9183 32963
rect 9125 32923 9183 32929
rect 8956 32824 8984 32923
rect 9214 32920 9220 32972
rect 9272 32920 9278 32972
rect 9582 32920 9588 32972
rect 9640 32920 9646 32972
rect 9692 32969 9720 33000
rect 10042 32988 10048 33000
rect 10100 32988 10106 33040
rect 10134 32988 10140 33040
rect 10192 33028 10198 33040
rect 10505 33031 10563 33037
rect 10192 33000 10466 33028
rect 10192 32988 10198 33000
rect 9677 32963 9735 32969
rect 9677 32929 9689 32963
rect 9723 32929 9735 32963
rect 9677 32923 9735 32929
rect 9769 32963 9827 32969
rect 9769 32929 9781 32963
rect 9815 32929 9827 32963
rect 9769 32923 9827 32929
rect 9784 32892 9812 32923
rect 9950 32920 9956 32972
rect 10008 32920 10014 32972
rect 10438 32960 10466 33000
rect 10505 32997 10517 33031
rect 10551 33028 10563 33031
rect 10870 33028 10876 33040
rect 10551 33000 10876 33028
rect 10551 32997 10563 33000
rect 10505 32991 10563 32997
rect 10870 32988 10876 33000
rect 10928 33028 10934 33040
rect 12618 33028 12624 33040
rect 10928 33000 12624 33028
rect 10928 32988 10934 33000
rect 12618 32988 12624 33000
rect 12676 33028 12682 33040
rect 12713 33031 12771 33037
rect 12713 33028 12725 33031
rect 12676 33000 12725 33028
rect 12676 32988 12682 33000
rect 12713 32997 12725 33000
rect 12759 32997 12771 33031
rect 12713 32991 12771 32997
rect 10438 32932 10640 32960
rect 10502 32892 10508 32904
rect 9784 32864 10508 32892
rect 10502 32852 10508 32864
rect 10560 32852 10566 32904
rect 10612 32901 10640 32932
rect 10778 32920 10784 32972
rect 10836 32960 10842 32972
rect 11330 32960 11336 32972
rect 10836 32932 11336 32960
rect 10836 32920 10842 32932
rect 11330 32920 11336 32932
rect 11388 32960 11394 32972
rect 11517 32963 11575 32969
rect 11517 32960 11529 32963
rect 11388 32932 11529 32960
rect 11388 32920 11394 32932
rect 11517 32929 11529 32932
rect 11563 32929 11575 32963
rect 11517 32923 11575 32929
rect 11609 32963 11667 32969
rect 11609 32929 11621 32963
rect 11655 32960 11667 32963
rect 11790 32960 11796 32972
rect 11655 32932 11796 32960
rect 11655 32929 11667 32932
rect 11609 32923 11667 32929
rect 11790 32920 11796 32932
rect 11848 32920 11854 32972
rect 13096 32960 13124 33059
rect 16666 33056 16672 33108
rect 16724 33096 16730 33108
rect 16761 33099 16819 33105
rect 16761 33096 16773 33099
rect 16724 33068 16773 33096
rect 16724 33056 16730 33068
rect 16761 33065 16773 33068
rect 16807 33065 16819 33099
rect 16761 33059 16819 33065
rect 16850 33056 16856 33108
rect 16908 33096 16914 33108
rect 18877 33099 18935 33105
rect 16908 33068 18828 33096
rect 16908 33056 16914 33068
rect 14182 32988 14188 33040
rect 14240 32988 14246 33040
rect 15013 33031 15071 33037
rect 15013 32997 15025 33031
rect 15059 33028 15071 33031
rect 15194 33028 15200 33040
rect 15059 33000 15200 33028
rect 15059 32997 15071 33000
rect 15013 32991 15071 32997
rect 15194 32988 15200 33000
rect 15252 33028 15258 33040
rect 16482 33028 16488 33040
rect 15252 33000 16488 33028
rect 15252 32988 15258 33000
rect 16482 32988 16488 33000
rect 16540 32988 16546 33040
rect 16574 32988 16580 33040
rect 16632 32988 16638 33040
rect 18800 33028 18828 33068
rect 18877 33065 18889 33099
rect 18923 33096 18935 33099
rect 19058 33096 19064 33108
rect 18923 33068 19064 33096
rect 18923 33065 18935 33068
rect 18877 33059 18935 33065
rect 19058 33056 19064 33068
rect 19116 33096 19122 33108
rect 20073 33099 20131 33105
rect 19116 33068 19656 33096
rect 19116 33056 19122 33068
rect 19628 33037 19656 33068
rect 20073 33065 20085 33099
rect 20119 33096 20131 33099
rect 21818 33096 21824 33108
rect 20119 33068 21824 33096
rect 20119 33065 20131 33068
rect 20073 33059 20131 33065
rect 21818 33056 21824 33068
rect 21876 33056 21882 33108
rect 22554 33056 22560 33108
rect 22612 33056 22618 33108
rect 24210 33056 24216 33108
rect 24268 33056 24274 33108
rect 24765 33099 24823 33105
rect 24765 33065 24777 33099
rect 24811 33096 24823 33099
rect 24854 33096 24860 33108
rect 24811 33068 24860 33096
rect 24811 33065 24823 33068
rect 24765 33059 24823 33065
rect 24854 33056 24860 33068
rect 24912 33056 24918 33108
rect 26418 33056 26424 33108
rect 26476 33056 26482 33108
rect 26605 33099 26663 33105
rect 26605 33065 26617 33099
rect 26651 33096 26663 33099
rect 27522 33096 27528 33108
rect 26651 33068 27528 33096
rect 26651 33065 26663 33068
rect 26605 33059 26663 33065
rect 27522 33056 27528 33068
rect 27580 33056 27586 33108
rect 29086 33056 29092 33108
rect 29144 33056 29150 33108
rect 19613 33031 19671 33037
rect 18800 33000 19288 33028
rect 13357 32963 13415 32969
rect 13357 32960 13369 32963
rect 13096 32932 13369 32960
rect 13357 32929 13369 32932
rect 13403 32929 13415 32963
rect 13357 32923 13415 32929
rect 13446 32920 13452 32972
rect 13504 32920 13510 32972
rect 13630 32920 13636 32972
rect 13688 32920 13694 32972
rect 13725 32963 13783 32969
rect 13725 32929 13737 32963
rect 13771 32960 13783 32963
rect 13814 32960 13820 32972
rect 13771 32932 13820 32960
rect 13771 32929 13783 32932
rect 13725 32923 13783 32929
rect 13814 32920 13820 32932
rect 13872 32960 13878 32972
rect 14642 32960 14648 32972
rect 13872 32932 14648 32960
rect 13872 32920 13878 32932
rect 14642 32920 14648 32932
rect 14700 32920 14706 32972
rect 15378 32920 15384 32972
rect 15436 32920 15442 32972
rect 16022 32920 16028 32972
rect 16080 32960 16086 32972
rect 16592 32960 16620 32988
rect 16853 32963 16911 32969
rect 16853 32960 16865 32963
rect 16080 32932 16865 32960
rect 16080 32920 16086 32932
rect 16853 32929 16865 32932
rect 16899 32929 16911 32963
rect 16853 32923 16911 32929
rect 18414 32920 18420 32972
rect 18472 32960 18478 32972
rect 19260 32969 19288 33000
rect 19613 32997 19625 33031
rect 19659 32997 19671 33031
rect 26326 33028 26332 33040
rect 19613 32991 19671 32997
rect 25240 33000 26332 33028
rect 19091 32963 19149 32969
rect 19091 32960 19103 32963
rect 18472 32932 19103 32960
rect 18472 32920 18478 32932
rect 19091 32929 19103 32932
rect 19137 32929 19149 32963
rect 19091 32923 19149 32929
rect 19245 32963 19303 32969
rect 19245 32929 19257 32963
rect 19291 32929 19303 32963
rect 19245 32923 19303 32929
rect 19889 32963 19947 32969
rect 19889 32929 19901 32963
rect 19935 32960 19947 32963
rect 21450 32960 21456 32972
rect 19935 32932 21456 32960
rect 19935 32929 19947 32932
rect 19889 32923 19947 32929
rect 21450 32920 21456 32932
rect 21508 32920 21514 32972
rect 22002 32920 22008 32972
rect 22060 32960 22066 32972
rect 22189 32963 22247 32969
rect 22189 32960 22201 32963
rect 22060 32932 22201 32960
rect 22060 32920 22066 32932
rect 22189 32929 22201 32932
rect 22235 32929 22247 32963
rect 22189 32923 22247 32929
rect 22373 32963 22431 32969
rect 22373 32929 22385 32963
rect 22419 32960 22431 32963
rect 22462 32960 22468 32972
rect 22419 32932 22468 32960
rect 22419 32929 22431 32932
rect 22373 32923 22431 32929
rect 22462 32920 22468 32932
rect 22520 32920 22526 32972
rect 24118 32920 24124 32972
rect 24176 32960 24182 32972
rect 24213 32963 24271 32969
rect 24213 32960 24225 32963
rect 24176 32932 24225 32960
rect 24176 32920 24182 32932
rect 24213 32929 24225 32932
rect 24259 32929 24271 32963
rect 24213 32923 24271 32929
rect 24397 32963 24455 32969
rect 24397 32929 24409 32963
rect 24443 32929 24455 32963
rect 24397 32923 24455 32929
rect 10597 32895 10655 32901
rect 10597 32861 10609 32895
rect 10643 32892 10655 32895
rect 11701 32895 11759 32901
rect 11701 32892 11713 32895
rect 10643 32864 11713 32892
rect 10643 32861 10655 32864
rect 10597 32855 10655 32861
rect 11701 32861 11713 32864
rect 11747 32892 11759 32895
rect 12437 32895 12495 32901
rect 12437 32892 12449 32895
rect 11747 32864 12449 32892
rect 11747 32861 11759 32864
rect 11701 32855 11759 32861
rect 12437 32861 12449 32864
rect 12483 32861 12495 32895
rect 12437 32855 12495 32861
rect 12621 32895 12679 32901
rect 12621 32861 12633 32895
rect 12667 32892 12679 32895
rect 12710 32892 12716 32904
rect 12667 32864 12716 32892
rect 12667 32861 12679 32864
rect 12621 32855 12679 32861
rect 12710 32852 12716 32864
rect 12768 32852 12774 32904
rect 16298 32852 16304 32904
rect 16356 32852 16362 32904
rect 16393 32895 16451 32901
rect 16393 32861 16405 32895
rect 16439 32861 16451 32895
rect 16393 32855 16451 32861
rect 16485 32895 16543 32901
rect 16485 32861 16497 32895
rect 16531 32861 16543 32895
rect 16485 32855 16543 32861
rect 16577 32895 16635 32901
rect 16577 32861 16589 32895
rect 16623 32892 16635 32895
rect 16942 32892 16948 32904
rect 16623 32864 16948 32892
rect 16623 32861 16635 32864
rect 16577 32855 16635 32861
rect 8956 32796 10548 32824
rect 10520 32768 10548 32796
rect 15194 32784 15200 32836
rect 15252 32784 15258 32836
rect 8665 32759 8723 32765
rect 8665 32725 8677 32759
rect 8711 32756 8723 32759
rect 9398 32756 9404 32768
rect 8711 32728 9404 32756
rect 8711 32725 8723 32728
rect 8665 32719 8723 32725
rect 9398 32716 9404 32728
rect 9456 32716 9462 32768
rect 10045 32759 10103 32765
rect 10045 32725 10057 32759
rect 10091 32756 10103 32759
rect 10410 32756 10416 32768
rect 10091 32728 10416 32756
rect 10091 32725 10103 32728
rect 10045 32719 10103 32725
rect 10410 32716 10416 32728
rect 10468 32716 10474 32768
rect 10502 32716 10508 32768
rect 10560 32716 10566 32768
rect 11149 32759 11207 32765
rect 11149 32725 11161 32759
rect 11195 32756 11207 32759
rect 11330 32756 11336 32768
rect 11195 32728 11336 32756
rect 11195 32725 11207 32728
rect 11149 32719 11207 32725
rect 11330 32716 11336 32728
rect 11388 32716 11394 32768
rect 11422 32716 11428 32768
rect 11480 32756 11486 32768
rect 12342 32756 12348 32768
rect 11480 32728 12348 32756
rect 11480 32716 11486 32728
rect 12342 32716 12348 32728
rect 12400 32716 12406 32768
rect 12526 32716 12532 32768
rect 12584 32756 12590 32768
rect 13173 32759 13231 32765
rect 13173 32756 13185 32759
rect 12584 32728 13185 32756
rect 12584 32716 12590 32728
rect 13173 32725 13185 32728
rect 13219 32725 13231 32759
rect 16408 32756 16436 32855
rect 16500 32824 16528 32855
rect 16942 32852 16948 32864
rect 17000 32892 17006 32904
rect 17678 32892 17684 32904
rect 17000 32864 17684 32892
rect 17000 32852 17006 32864
rect 17678 32852 17684 32864
rect 17736 32852 17742 32904
rect 19702 32852 19708 32904
rect 19760 32852 19766 32904
rect 21174 32852 21180 32904
rect 21232 32892 21238 32904
rect 22020 32892 22048 32920
rect 21232 32864 22048 32892
rect 21232 32852 21238 32864
rect 16758 32824 16764 32836
rect 16500 32796 16764 32824
rect 16758 32784 16764 32796
rect 16816 32784 16822 32836
rect 24228 32824 24256 32923
rect 24412 32892 24440 32923
rect 24946 32920 24952 32972
rect 25004 32920 25010 32972
rect 25240 32969 25268 33000
rect 26326 32988 26332 33000
rect 26384 32988 26390 33040
rect 27985 33031 28043 33037
rect 27985 32997 27997 33031
rect 28031 33028 28043 33031
rect 28902 33028 28908 33040
rect 28031 33000 28908 33028
rect 28031 32997 28043 33000
rect 27985 32991 28043 32997
rect 28902 32988 28908 33000
rect 28960 33028 28966 33040
rect 28960 33000 29684 33028
rect 28960 32988 28966 33000
rect 25225 32963 25283 32969
rect 25225 32929 25237 32963
rect 25271 32929 25283 32963
rect 25225 32923 25283 32929
rect 25593 32963 25651 32969
rect 25593 32929 25605 32963
rect 25639 32960 25651 32963
rect 25682 32960 25688 32972
rect 25639 32932 25688 32960
rect 25639 32929 25651 32932
rect 25593 32923 25651 32929
rect 25682 32920 25688 32932
rect 25740 32920 25746 32972
rect 26145 32963 26203 32969
rect 26145 32929 26157 32963
rect 26191 32960 26203 32963
rect 26602 32960 26608 32972
rect 26191 32932 26608 32960
rect 26191 32929 26203 32932
rect 26145 32923 26203 32929
rect 26602 32920 26608 32932
rect 26660 32920 26666 32972
rect 26878 32920 26884 32972
rect 26936 32960 26942 32972
rect 26973 32963 27031 32969
rect 26973 32960 26985 32963
rect 26936 32932 26985 32960
rect 26936 32920 26942 32932
rect 26973 32929 26985 32932
rect 27019 32960 27031 32963
rect 27430 32960 27436 32972
rect 27019 32932 27436 32960
rect 27019 32929 27031 32932
rect 26973 32923 27031 32929
rect 27430 32920 27436 32932
rect 27488 32920 27494 32972
rect 28350 32920 28356 32972
rect 28408 32920 28414 32972
rect 29656 32969 29684 33000
rect 29641 32963 29699 32969
rect 29641 32929 29653 32963
rect 29687 32929 29699 32963
rect 29641 32923 29699 32929
rect 25038 32892 25044 32904
rect 24412 32864 25044 32892
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 25130 32852 25136 32904
rect 25188 32892 25194 32904
rect 25409 32895 25467 32901
rect 25409 32892 25421 32895
rect 25188 32864 25421 32892
rect 25188 32852 25194 32864
rect 25409 32861 25421 32864
rect 25455 32861 25467 32895
rect 25409 32855 25467 32861
rect 25869 32895 25927 32901
rect 25869 32861 25881 32895
rect 25915 32861 25927 32895
rect 27890 32892 27896 32904
rect 25869 32855 25927 32861
rect 26620 32864 27896 32892
rect 25884 32824 25912 32855
rect 25961 32827 26019 32833
rect 25961 32824 25973 32827
rect 24228 32796 25973 32824
rect 25961 32793 25973 32796
rect 26007 32793 26019 32827
rect 25961 32787 26019 32793
rect 17034 32756 17040 32768
rect 16408 32728 17040 32756
rect 13173 32719 13231 32725
rect 17034 32716 17040 32728
rect 17092 32716 17098 32768
rect 19794 32716 19800 32768
rect 19852 32716 19858 32768
rect 25498 32716 25504 32768
rect 25556 32756 25562 32768
rect 26620 32765 26648 32864
rect 27890 32852 27896 32864
rect 27948 32852 27954 32904
rect 27617 32827 27675 32833
rect 27617 32793 27629 32827
rect 27663 32824 27675 32827
rect 28442 32824 28448 32836
rect 27663 32796 28448 32824
rect 27663 32793 27675 32796
rect 27617 32787 27675 32793
rect 28442 32784 28448 32796
rect 28500 32784 28506 32836
rect 25777 32759 25835 32765
rect 25777 32756 25789 32759
rect 25556 32728 25789 32756
rect 25556 32716 25562 32728
rect 25777 32725 25789 32728
rect 25823 32725 25835 32759
rect 25777 32719 25835 32725
rect 26605 32759 26663 32765
rect 26605 32725 26617 32759
rect 26651 32725 26663 32759
rect 26605 32719 26663 32725
rect 27525 32759 27583 32765
rect 27525 32725 27537 32759
rect 27571 32756 27583 32759
rect 27706 32756 27712 32768
rect 27571 32728 27712 32756
rect 27571 32725 27583 32728
rect 27525 32719 27583 32725
rect 27706 32716 27712 32728
rect 27764 32716 27770 32768
rect 28994 32716 29000 32768
rect 29052 32716 29058 32768
rect 552 32666 31648 32688
rect 552 32614 3662 32666
rect 3714 32614 3726 32666
rect 3778 32614 3790 32666
rect 3842 32614 3854 32666
rect 3906 32614 3918 32666
rect 3970 32614 11436 32666
rect 11488 32614 11500 32666
rect 11552 32614 11564 32666
rect 11616 32614 11628 32666
rect 11680 32614 11692 32666
rect 11744 32614 19210 32666
rect 19262 32614 19274 32666
rect 19326 32614 19338 32666
rect 19390 32614 19402 32666
rect 19454 32614 19466 32666
rect 19518 32614 26984 32666
rect 27036 32614 27048 32666
rect 27100 32614 27112 32666
rect 27164 32614 27176 32666
rect 27228 32614 27240 32666
rect 27292 32614 31648 32666
rect 552 32592 31648 32614
rect 8846 32512 8852 32564
rect 8904 32552 8910 32564
rect 9401 32555 9459 32561
rect 9401 32552 9413 32555
rect 8904 32524 9413 32552
rect 8904 32512 8910 32524
rect 9401 32521 9413 32524
rect 9447 32521 9459 32555
rect 9401 32515 9459 32521
rect 9858 32512 9864 32564
rect 9916 32552 9922 32564
rect 10778 32552 10784 32564
rect 9916 32524 10784 32552
rect 9916 32512 9922 32524
rect 10778 32512 10784 32524
rect 10836 32512 10842 32564
rect 11238 32512 11244 32564
rect 11296 32552 11302 32564
rect 13446 32552 13452 32564
rect 11296 32524 13452 32552
rect 11296 32512 11302 32524
rect 13446 32512 13452 32524
rect 13504 32512 13510 32564
rect 15378 32512 15384 32564
rect 15436 32552 15442 32564
rect 15838 32552 15844 32564
rect 15436 32524 15844 32552
rect 15436 32512 15442 32524
rect 15838 32512 15844 32524
rect 15896 32512 15902 32564
rect 16114 32512 16120 32564
rect 16172 32552 16178 32564
rect 16172 32524 16620 32552
rect 16172 32512 16178 32524
rect 9214 32444 9220 32496
rect 9272 32484 9278 32496
rect 13814 32484 13820 32496
rect 9272 32456 13820 32484
rect 9272 32444 9278 32456
rect 10045 32419 10103 32425
rect 10045 32385 10057 32419
rect 10091 32416 10103 32419
rect 10134 32416 10140 32428
rect 10091 32388 10140 32416
rect 10091 32385 10103 32388
rect 10045 32379 10103 32385
rect 10134 32376 10140 32388
rect 10192 32376 10198 32428
rect 9674 32308 9680 32360
rect 9732 32348 9738 32360
rect 9769 32351 9827 32357
rect 9769 32348 9781 32351
rect 9732 32320 9781 32348
rect 9732 32308 9738 32320
rect 9769 32317 9781 32320
rect 9815 32348 9827 32351
rect 9815 32320 10088 32348
rect 9815 32317 9827 32320
rect 9769 32311 9827 32317
rect 10060 32292 10088 32320
rect 10410 32308 10416 32360
rect 10468 32308 10474 32360
rect 10502 32308 10508 32360
rect 10560 32308 10566 32360
rect 10686 32308 10692 32360
rect 10744 32308 10750 32360
rect 10980 32357 11008 32456
rect 13814 32444 13820 32456
rect 13872 32444 13878 32496
rect 16592 32484 16620 32524
rect 16666 32512 16672 32564
rect 16724 32552 16730 32564
rect 17129 32555 17187 32561
rect 17129 32552 17141 32555
rect 16724 32524 17141 32552
rect 16724 32512 16730 32524
rect 17129 32521 17141 32524
rect 17175 32521 17187 32555
rect 17129 32515 17187 32521
rect 17678 32512 17684 32564
rect 17736 32512 17742 32564
rect 18874 32512 18880 32564
rect 18932 32552 18938 32564
rect 18932 32524 21956 32552
rect 18932 32512 18938 32524
rect 16592 32456 17464 32484
rect 11790 32376 11796 32428
rect 11848 32416 11854 32428
rect 14277 32419 14335 32425
rect 11848 32388 12756 32416
rect 11848 32376 11854 32388
rect 10781 32351 10839 32357
rect 10781 32317 10793 32351
rect 10827 32348 10839 32351
rect 10965 32351 11023 32357
rect 10965 32348 10977 32351
rect 10827 32320 10977 32348
rect 10827 32317 10839 32320
rect 10781 32311 10839 32317
rect 10965 32317 10977 32320
rect 11011 32317 11023 32351
rect 10965 32311 11023 32317
rect 11054 32308 11060 32360
rect 11112 32308 11118 32360
rect 11238 32308 11244 32360
rect 11296 32308 11302 32360
rect 11330 32308 11336 32360
rect 11388 32308 11394 32360
rect 12342 32308 12348 32360
rect 12400 32308 12406 32360
rect 12526 32308 12532 32360
rect 12584 32308 12590 32360
rect 12728 32357 12756 32388
rect 14277 32385 14289 32419
rect 14323 32416 14335 32419
rect 14461 32419 14519 32425
rect 14461 32416 14473 32419
rect 14323 32388 14473 32416
rect 14323 32385 14335 32388
rect 14277 32379 14335 32385
rect 14461 32385 14473 32388
rect 14507 32385 14519 32419
rect 14461 32379 14519 32385
rect 16114 32376 16120 32428
rect 16172 32376 16178 32428
rect 16209 32419 16267 32425
rect 16209 32385 16221 32419
rect 16255 32385 16267 32419
rect 16209 32379 16267 32385
rect 12621 32351 12679 32357
rect 12621 32317 12633 32351
rect 12667 32317 12679 32351
rect 12621 32311 12679 32317
rect 12713 32351 12771 32357
rect 12713 32317 12725 32351
rect 12759 32348 12771 32351
rect 12802 32348 12808 32360
rect 12759 32320 12808 32348
rect 12759 32317 12771 32320
rect 12713 32311 12771 32317
rect 10042 32240 10048 32292
rect 10100 32240 10106 32292
rect 10520 32280 10548 32308
rect 11256 32280 11284 32308
rect 10520 32252 11284 32280
rect 9674 32172 9680 32224
rect 9732 32212 9738 32224
rect 9858 32212 9864 32224
rect 9732 32184 9864 32212
rect 9732 32172 9738 32184
rect 9858 32172 9864 32184
rect 9916 32172 9922 32224
rect 9950 32172 9956 32224
rect 10008 32212 10014 32224
rect 10229 32215 10287 32221
rect 10229 32212 10241 32215
rect 10008 32184 10241 32212
rect 10008 32172 10014 32184
rect 10229 32181 10241 32184
rect 10275 32181 10287 32215
rect 10229 32175 10287 32181
rect 11238 32172 11244 32224
rect 11296 32212 11302 32224
rect 11517 32215 11575 32221
rect 11517 32212 11529 32215
rect 11296 32184 11529 32212
rect 11296 32172 11302 32184
rect 11517 32181 11529 32184
rect 11563 32181 11575 32215
rect 11517 32175 11575 32181
rect 11882 32172 11888 32224
rect 11940 32212 11946 32224
rect 12360 32212 12388 32308
rect 12434 32240 12440 32292
rect 12492 32280 12498 32292
rect 12636 32280 12664 32311
rect 12802 32308 12808 32320
rect 12860 32308 12866 32360
rect 14369 32351 14427 32357
rect 14369 32317 14381 32351
rect 14415 32348 14427 32351
rect 16022 32348 16028 32360
rect 14415 32320 16028 32348
rect 14415 32317 14427 32320
rect 14369 32311 14427 32317
rect 16022 32308 16028 32320
rect 16080 32308 16086 32360
rect 14728 32283 14786 32289
rect 12492 32252 12664 32280
rect 12912 32252 13952 32280
rect 12492 32240 12498 32252
rect 12912 32212 12940 32252
rect 11940 32184 12940 32212
rect 12989 32215 13047 32221
rect 11940 32172 11946 32184
rect 12989 32181 13001 32215
rect 13035 32212 13047 32215
rect 13814 32212 13820 32224
rect 13035 32184 13820 32212
rect 13035 32181 13047 32184
rect 12989 32175 13047 32181
rect 13814 32172 13820 32184
rect 13872 32172 13878 32224
rect 13924 32212 13952 32252
rect 14728 32249 14740 32283
rect 14774 32280 14786 32283
rect 14918 32280 14924 32292
rect 14774 32252 14924 32280
rect 14774 32249 14786 32252
rect 14728 32243 14786 32249
rect 14918 32240 14924 32252
rect 14976 32240 14982 32292
rect 16224 32280 16252 32379
rect 16390 32376 16396 32428
rect 16448 32376 16454 32428
rect 16301 32351 16359 32357
rect 16301 32317 16313 32351
rect 16347 32348 16359 32351
rect 17310 32348 17316 32360
rect 16347 32320 17316 32348
rect 16347 32317 16359 32320
rect 16301 32311 16359 32317
rect 17310 32308 17316 32320
rect 17368 32308 17374 32360
rect 17436 32357 17464 32456
rect 19426 32444 19432 32496
rect 19484 32484 19490 32496
rect 20162 32484 20168 32496
rect 19484 32456 20168 32484
rect 19484 32444 19490 32456
rect 20162 32444 20168 32456
rect 20220 32484 20226 32496
rect 20220 32456 20484 32484
rect 20220 32444 20226 32456
rect 18966 32416 18972 32428
rect 17880 32388 18972 32416
rect 17405 32351 17464 32357
rect 17405 32317 17417 32351
rect 17451 32320 17464 32351
rect 17451 32317 17463 32320
rect 17405 32311 17463 32317
rect 17494 32308 17500 32360
rect 17552 32348 17558 32360
rect 17880 32357 17908 32388
rect 18966 32376 18972 32388
rect 19024 32376 19030 32428
rect 20456 32416 20484 32456
rect 20898 32444 20904 32496
rect 20956 32484 20962 32496
rect 21818 32484 21824 32496
rect 20956 32456 21824 32484
rect 20956 32444 20962 32456
rect 21818 32444 21824 32456
rect 21876 32444 21882 32496
rect 20625 32419 20683 32425
rect 20625 32416 20637 32419
rect 20456 32388 20637 32416
rect 20625 32385 20637 32388
rect 20671 32385 20683 32419
rect 21928 32416 21956 32524
rect 22462 32512 22468 32564
rect 22520 32512 22526 32564
rect 23474 32552 23480 32564
rect 22572 32524 23480 32552
rect 22002 32416 22008 32428
rect 21928 32388 22008 32416
rect 20625 32379 20683 32385
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22572 32416 22600 32524
rect 23474 32512 23480 32524
rect 23532 32512 23538 32564
rect 28813 32555 28871 32561
rect 28813 32521 28825 32555
rect 28859 32552 28871 32555
rect 28902 32552 28908 32564
rect 28859 32524 28908 32552
rect 28859 32521 28871 32524
rect 28813 32515 28871 32521
rect 28902 32512 28908 32524
rect 28960 32512 28966 32564
rect 24394 32484 24400 32496
rect 22112 32388 22600 32416
rect 22756 32456 24400 32484
rect 17589 32351 17647 32357
rect 17589 32348 17601 32351
rect 17552 32320 17601 32348
rect 17552 32308 17558 32320
rect 17589 32317 17601 32320
rect 17635 32317 17647 32351
rect 17589 32311 17647 32317
rect 17865 32351 17923 32357
rect 17865 32317 17877 32351
rect 17911 32317 17923 32351
rect 17865 32311 17923 32317
rect 16758 32280 16764 32292
rect 16224 32252 16764 32280
rect 16758 32240 16764 32252
rect 16816 32240 16822 32292
rect 16942 32240 16948 32292
rect 17000 32240 17006 32292
rect 17161 32283 17219 32289
rect 17161 32249 17173 32283
rect 17207 32280 17219 32283
rect 17880 32280 17908 32311
rect 17954 32308 17960 32360
rect 18012 32348 18018 32360
rect 19058 32348 19064 32360
rect 18012 32320 19064 32348
rect 18012 32308 18018 32320
rect 19058 32308 19064 32320
rect 19116 32348 19122 32360
rect 19613 32351 19671 32357
rect 19613 32348 19625 32351
rect 19116 32320 19625 32348
rect 19116 32308 19122 32320
rect 19613 32317 19625 32320
rect 19659 32317 19671 32351
rect 19613 32311 19671 32317
rect 20162 32308 20168 32360
rect 20220 32308 20226 32360
rect 20254 32308 20260 32360
rect 20312 32308 20318 32360
rect 20732 32357 20852 32358
rect 20705 32351 20852 32357
rect 20705 32317 20717 32351
rect 20751 32348 20852 32351
rect 21082 32348 21088 32360
rect 20751 32330 21088 32348
rect 20751 32317 20763 32330
rect 20824 32320 21088 32330
rect 20705 32311 20763 32317
rect 21082 32308 21088 32320
rect 21140 32308 21146 32360
rect 21174 32308 21180 32360
rect 21232 32308 21238 32360
rect 21266 32308 21272 32360
rect 21324 32308 21330 32360
rect 21726 32308 21732 32360
rect 21784 32348 21790 32360
rect 22112 32348 22140 32388
rect 21784 32320 22140 32348
rect 21784 32308 21790 32320
rect 22186 32308 22192 32360
rect 22244 32308 22250 32360
rect 22554 32308 22560 32360
rect 22612 32348 22618 32360
rect 22756 32357 22784 32456
rect 24394 32444 24400 32456
rect 24452 32484 24458 32496
rect 24452 32456 25268 32484
rect 24452 32444 24458 32456
rect 22649 32351 22707 32357
rect 22649 32348 22661 32351
rect 22612 32320 22661 32348
rect 22612 32308 22618 32320
rect 22649 32317 22661 32320
rect 22695 32317 22707 32351
rect 22649 32311 22707 32317
rect 22741 32351 22799 32357
rect 22741 32317 22753 32351
rect 22787 32317 22799 32351
rect 22741 32311 22799 32317
rect 22830 32308 22836 32360
rect 22888 32308 22894 32360
rect 23014 32357 23020 32360
rect 22971 32351 23020 32357
rect 22971 32317 22983 32351
rect 23017 32317 23020 32351
rect 22971 32311 23020 32317
rect 23014 32308 23020 32311
rect 23072 32308 23078 32360
rect 23106 32308 23112 32360
rect 23164 32308 23170 32360
rect 23385 32351 23443 32357
rect 23385 32317 23397 32351
rect 23431 32348 23443 32351
rect 23474 32348 23480 32360
rect 23431 32320 23480 32348
rect 23431 32317 23443 32320
rect 23385 32311 23443 32317
rect 23474 32308 23480 32320
rect 23532 32308 23538 32360
rect 25240 32357 25268 32456
rect 25225 32351 25283 32357
rect 25225 32317 25237 32351
rect 25271 32317 25283 32351
rect 25225 32311 25283 32317
rect 26234 32308 26240 32360
rect 26292 32348 26298 32360
rect 27157 32351 27215 32357
rect 27157 32348 27169 32351
rect 26292 32320 27169 32348
rect 26292 32308 26298 32320
rect 27157 32317 27169 32320
rect 27203 32317 27215 32351
rect 27157 32311 27215 32317
rect 27249 32351 27307 32357
rect 27249 32317 27261 32351
rect 27295 32348 27307 32351
rect 27433 32351 27491 32357
rect 27433 32348 27445 32351
rect 27295 32320 27445 32348
rect 27295 32317 27307 32320
rect 27249 32311 27307 32317
rect 27433 32317 27445 32320
rect 27479 32317 27491 32351
rect 28997 32351 29055 32357
rect 28997 32348 29009 32351
rect 27433 32311 27491 32317
rect 27540 32320 29009 32348
rect 17207 32252 17908 32280
rect 17207 32249 17219 32252
rect 17161 32243 17219 32249
rect 19150 32240 19156 32292
rect 19208 32280 19214 32292
rect 19981 32283 20039 32289
rect 19981 32280 19993 32283
rect 19208 32252 19993 32280
rect 19208 32240 19214 32252
rect 19981 32249 19993 32252
rect 20027 32249 20039 32283
rect 19981 32243 20039 32249
rect 20070 32240 20076 32292
rect 20128 32280 20134 32292
rect 20349 32283 20407 32289
rect 20349 32280 20361 32283
rect 20128 32252 20361 32280
rect 20128 32240 20134 32252
rect 20349 32249 20361 32252
rect 20395 32249 20407 32283
rect 20349 32243 20407 32249
rect 20487 32283 20545 32289
rect 20487 32249 20499 32283
rect 20533 32280 20545 32283
rect 20990 32280 20996 32292
rect 20533 32252 20996 32280
rect 20533 32249 20545 32252
rect 20487 32243 20545 32249
rect 20990 32240 20996 32252
rect 21048 32240 21054 32292
rect 27172 32280 27200 32311
rect 27338 32280 27344 32292
rect 27172 32252 27344 32280
rect 27338 32240 27344 32252
rect 27396 32280 27402 32292
rect 27540 32280 27568 32320
rect 28997 32317 29009 32320
rect 29043 32317 29055 32351
rect 28997 32311 29055 32317
rect 27706 32289 27712 32292
rect 27700 32280 27712 32289
rect 27396 32252 27568 32280
rect 27667 32252 27712 32280
rect 27396 32240 27402 32252
rect 27700 32243 27712 32252
rect 27706 32240 27712 32243
rect 27764 32240 27770 32292
rect 15654 32212 15660 32224
rect 13924 32184 15660 32212
rect 15654 32172 15660 32184
rect 15712 32172 15718 32224
rect 15930 32172 15936 32224
rect 15988 32172 15994 32224
rect 17310 32172 17316 32224
rect 17368 32172 17374 32224
rect 17402 32172 17408 32224
rect 17460 32212 17466 32224
rect 17497 32215 17555 32221
rect 17497 32212 17509 32215
rect 17460 32184 17509 32212
rect 17460 32172 17466 32184
rect 17497 32181 17509 32184
rect 17543 32181 17555 32215
rect 17497 32175 17555 32181
rect 19518 32172 19524 32224
rect 19576 32212 19582 32224
rect 19705 32215 19763 32221
rect 19705 32212 19717 32215
rect 19576 32184 19717 32212
rect 19576 32172 19582 32184
rect 19705 32181 19717 32184
rect 19751 32181 19763 32215
rect 19705 32175 19763 32181
rect 21453 32215 21511 32221
rect 21453 32181 21465 32215
rect 21499 32212 21511 32215
rect 21542 32212 21548 32224
rect 21499 32184 21548 32212
rect 21499 32181 21511 32184
rect 21453 32175 21511 32181
rect 21542 32172 21548 32184
rect 21600 32172 21606 32224
rect 21634 32172 21640 32224
rect 21692 32172 21698 32224
rect 22370 32172 22376 32224
rect 22428 32172 22434 32224
rect 23290 32172 23296 32224
rect 23348 32172 23354 32224
rect 25314 32172 25320 32224
rect 25372 32172 25378 32224
rect 29089 32215 29147 32221
rect 29089 32181 29101 32215
rect 29135 32212 29147 32215
rect 29362 32212 29368 32224
rect 29135 32184 29368 32212
rect 29135 32181 29147 32184
rect 29089 32175 29147 32181
rect 29362 32172 29368 32184
rect 29420 32172 29426 32224
rect 552 32122 31648 32144
rect 552 32070 4322 32122
rect 4374 32070 4386 32122
rect 4438 32070 4450 32122
rect 4502 32070 4514 32122
rect 4566 32070 4578 32122
rect 4630 32070 12096 32122
rect 12148 32070 12160 32122
rect 12212 32070 12224 32122
rect 12276 32070 12288 32122
rect 12340 32070 12352 32122
rect 12404 32070 19870 32122
rect 19922 32070 19934 32122
rect 19986 32070 19998 32122
rect 20050 32070 20062 32122
rect 20114 32070 20126 32122
rect 20178 32070 27644 32122
rect 27696 32070 27708 32122
rect 27760 32070 27772 32122
rect 27824 32070 27836 32122
rect 27888 32070 27900 32122
rect 27952 32070 31648 32122
rect 552 32048 31648 32070
rect 10781 32011 10839 32017
rect 10781 31977 10793 32011
rect 10827 32008 10839 32011
rect 10962 32008 10968 32020
rect 10827 31980 10968 32008
rect 10827 31977 10839 31980
rect 10781 31971 10839 31977
rect 10962 31968 10968 31980
rect 11020 31968 11026 32020
rect 14918 31968 14924 32020
rect 14976 31968 14982 32020
rect 15657 32011 15715 32017
rect 15657 32008 15669 32011
rect 15120 31980 15669 32008
rect 10226 31900 10232 31952
rect 10284 31940 10290 31952
rect 10413 31943 10471 31949
rect 10413 31940 10425 31943
rect 10284 31912 10425 31940
rect 10284 31900 10290 31912
rect 10413 31909 10425 31912
rect 10459 31909 10471 31943
rect 10413 31903 10471 31909
rect 10597 31943 10655 31949
rect 10597 31909 10609 31943
rect 10643 31940 10655 31943
rect 10870 31940 10876 31952
rect 10643 31912 10876 31940
rect 10643 31909 10655 31912
rect 10597 31903 10655 31909
rect 10870 31900 10876 31912
rect 10928 31940 10934 31952
rect 11330 31940 11336 31952
rect 10928 31912 11336 31940
rect 10928 31900 10934 31912
rect 11330 31900 11336 31912
rect 11388 31900 11394 31952
rect 14458 31900 14464 31952
rect 14516 31940 14522 31952
rect 15120 31940 15148 31980
rect 15657 31977 15669 31980
rect 15703 31977 15715 32011
rect 15657 31971 15715 31977
rect 16485 32011 16543 32017
rect 16485 31977 16497 32011
rect 16531 32008 16543 32011
rect 16758 32008 16764 32020
rect 16531 31980 16764 32008
rect 16531 31977 16543 31980
rect 16485 31971 16543 31977
rect 16758 31968 16764 31980
rect 16816 31968 16822 32020
rect 17310 31968 17316 32020
rect 17368 32008 17374 32020
rect 20901 32011 20959 32017
rect 17368 31980 18000 32008
rect 17368 31968 17374 31980
rect 15930 31940 15936 31952
rect 14516 31912 15148 31940
rect 15396 31912 15936 31940
rect 14516 31900 14522 31912
rect 9122 31832 9128 31884
rect 9180 31832 9186 31884
rect 12621 31875 12679 31881
rect 12621 31841 12633 31875
rect 12667 31872 12679 31875
rect 12710 31872 12716 31884
rect 12667 31844 12716 31872
rect 12667 31841 12679 31844
rect 12621 31835 12679 31841
rect 12710 31832 12716 31844
rect 12768 31832 12774 31884
rect 13538 31832 13544 31884
rect 13596 31832 13602 31884
rect 13722 31881 13728 31884
rect 13679 31875 13728 31881
rect 13679 31841 13691 31875
rect 13725 31841 13728 31875
rect 13679 31835 13728 31841
rect 13722 31832 13728 31835
rect 13780 31832 13786 31884
rect 15194 31832 15200 31884
rect 15252 31832 15258 31884
rect 15286 31832 15292 31884
rect 15344 31832 15350 31884
rect 15396 31881 15424 31912
rect 15930 31900 15936 31912
rect 15988 31900 15994 31952
rect 16666 31949 16672 31952
rect 16653 31943 16672 31949
rect 16653 31909 16665 31943
rect 16653 31903 16672 31909
rect 16666 31900 16672 31903
rect 16724 31900 16730 31952
rect 16853 31943 16911 31949
rect 16853 31909 16865 31943
rect 16899 31940 16911 31943
rect 16945 31943 17003 31949
rect 16945 31940 16957 31943
rect 16899 31912 16957 31940
rect 16899 31909 16911 31912
rect 16853 31903 16911 31909
rect 16945 31909 16957 31912
rect 16991 31940 17003 31943
rect 16991 31912 17540 31940
rect 16991 31909 17003 31912
rect 16945 31903 17003 31909
rect 15381 31875 15439 31881
rect 15381 31841 15393 31875
rect 15427 31841 15439 31875
rect 15381 31835 15439 31841
rect 15565 31875 15623 31881
rect 15565 31841 15577 31875
rect 15611 31872 15623 31875
rect 15654 31872 15660 31884
rect 15611 31844 15660 31872
rect 15611 31841 15623 31844
rect 15565 31835 15623 31841
rect 15654 31832 15660 31844
rect 15712 31832 15718 31884
rect 15746 31832 15752 31884
rect 15804 31872 15810 31884
rect 17512 31881 17540 31912
rect 17972 31881 18000 31980
rect 20901 31977 20913 32011
rect 20947 32008 20959 32011
rect 21358 32008 21364 32020
rect 20947 31980 21364 32008
rect 20947 31977 20959 31980
rect 20901 31971 20959 31977
rect 21358 31968 21364 31980
rect 21416 32008 21422 32020
rect 24213 32011 24271 32017
rect 21416 31980 23704 32008
rect 21416 31968 21422 31980
rect 19061 31943 19119 31949
rect 19061 31909 19073 31943
rect 19107 31940 19119 31943
rect 19766 31943 19824 31949
rect 19766 31940 19778 31943
rect 19107 31912 19778 31940
rect 19107 31909 19119 31912
rect 19061 31903 19119 31909
rect 19766 31909 19778 31912
rect 19812 31909 19824 31943
rect 21634 31940 21640 31952
rect 19766 31903 19824 31909
rect 21284 31912 21640 31940
rect 15841 31875 15899 31881
rect 15841 31872 15853 31875
rect 15804 31844 15853 31872
rect 15804 31832 15810 31844
rect 15841 31841 15853 31844
rect 15887 31841 15899 31875
rect 17129 31875 17187 31881
rect 17129 31872 17141 31875
rect 15841 31835 15899 31841
rect 16868 31844 17141 31872
rect 16868 31816 16896 31844
rect 17129 31841 17141 31844
rect 17175 31841 17187 31875
rect 17129 31835 17187 31841
rect 17497 31875 17555 31881
rect 17497 31841 17509 31875
rect 17543 31841 17555 31875
rect 17497 31835 17555 31841
rect 17865 31875 17923 31881
rect 17865 31841 17877 31875
rect 17911 31841 17923 31875
rect 17865 31835 17923 31841
rect 17957 31875 18015 31881
rect 17957 31841 17969 31875
rect 18003 31841 18015 31875
rect 17957 31835 18015 31841
rect 12802 31764 12808 31816
rect 12860 31764 12866 31816
rect 13265 31807 13323 31813
rect 13265 31773 13277 31807
rect 13311 31773 13323 31807
rect 13265 31767 13323 31773
rect 13817 31807 13875 31813
rect 13817 31773 13829 31807
rect 13863 31804 13875 31807
rect 14550 31804 14556 31816
rect 13863 31776 14556 31804
rect 13863 31773 13875 31776
rect 13817 31767 13875 31773
rect 12710 31696 12716 31748
rect 12768 31736 12774 31748
rect 13280 31736 13308 31767
rect 14550 31764 14556 31776
rect 14608 31764 14614 31816
rect 16850 31764 16856 31816
rect 16908 31764 16914 31816
rect 17313 31807 17371 31813
rect 17313 31804 17325 31807
rect 17144 31776 17325 31804
rect 17144 31748 17172 31776
rect 17313 31773 17325 31776
rect 17359 31773 17371 31807
rect 17880 31804 17908 31835
rect 18046 31832 18052 31884
rect 18104 31872 18110 31884
rect 18874 31872 18880 31884
rect 18104 31844 18880 31872
rect 18104 31832 18110 31844
rect 18874 31832 18880 31844
rect 18932 31872 18938 31884
rect 18969 31875 19027 31881
rect 18969 31872 18981 31875
rect 18932 31844 18981 31872
rect 18932 31832 18938 31844
rect 18969 31841 18981 31844
rect 19015 31841 19027 31875
rect 18969 31835 19027 31841
rect 19150 31832 19156 31884
rect 19208 31832 19214 31884
rect 19518 31832 19524 31884
rect 19576 31832 19582 31884
rect 21284 31881 21312 31912
rect 21634 31900 21640 31912
rect 21692 31900 21698 31952
rect 23290 31940 23296 31952
rect 22756 31912 23296 31940
rect 21542 31881 21548 31884
rect 21269 31875 21327 31881
rect 21269 31841 21281 31875
rect 21315 31841 21327 31875
rect 21536 31872 21548 31881
rect 21503 31844 21548 31872
rect 21269 31835 21327 31841
rect 21536 31835 21548 31844
rect 21542 31832 21548 31835
rect 21600 31832 21606 31884
rect 22756 31881 22784 31912
rect 23290 31900 23296 31912
rect 23348 31900 23354 31952
rect 22741 31875 22799 31881
rect 22741 31841 22753 31875
rect 22787 31841 22799 31875
rect 22997 31875 23055 31881
rect 22997 31872 23009 31875
rect 22741 31835 22799 31841
rect 22848 31844 23009 31872
rect 19426 31804 19432 31816
rect 17880 31776 19432 31804
rect 17313 31767 17371 31773
rect 19426 31764 19432 31776
rect 19484 31764 19490 31816
rect 22370 31764 22376 31816
rect 22428 31804 22434 31816
rect 22848 31804 22876 31844
rect 22997 31841 23009 31844
rect 23043 31841 23055 31875
rect 23676 31872 23704 31980
rect 24213 31977 24225 32011
rect 24259 32008 24271 32011
rect 24302 32008 24308 32020
rect 24259 31980 24308 32008
rect 24259 31977 24271 31980
rect 24213 31971 24271 31977
rect 24302 31968 24308 31980
rect 24360 31968 24366 32020
rect 27985 32011 28043 32017
rect 27985 31977 27997 32011
rect 28031 32008 28043 32011
rect 28074 32008 28080 32020
rect 28031 31980 28080 32008
rect 28031 31977 28043 31980
rect 27985 31971 28043 31977
rect 28074 31968 28080 31980
rect 28132 31968 28138 32020
rect 24486 31900 24492 31952
rect 24544 31940 24550 31952
rect 24673 31943 24731 31949
rect 24673 31940 24685 31943
rect 24544 31912 24685 31940
rect 24544 31900 24550 31912
rect 24673 31909 24685 31912
rect 24719 31909 24731 31943
rect 24673 31903 24731 31909
rect 28994 31900 29000 31952
rect 29052 31940 29058 31952
rect 29098 31943 29156 31949
rect 29098 31940 29110 31943
rect 29052 31912 29110 31940
rect 29052 31900 29058 31912
rect 29098 31909 29110 31912
rect 29144 31909 29156 31943
rect 29098 31903 29156 31909
rect 24397 31875 24455 31881
rect 24397 31872 24409 31875
rect 23676 31844 24409 31872
rect 22997 31835 23055 31841
rect 24397 31841 24409 31844
rect 24443 31872 24455 31875
rect 24443 31844 24624 31872
rect 24443 31841 24455 31844
rect 24397 31835 24455 31841
rect 22428 31776 22876 31804
rect 24489 31807 24547 31813
rect 22428 31764 22434 31776
rect 24489 31773 24501 31807
rect 24535 31773 24547 31807
rect 24489 31767 24547 31773
rect 12768 31708 13308 31736
rect 12768 31696 12774 31708
rect 17126 31696 17132 31748
rect 17184 31696 17190 31748
rect 24026 31696 24032 31748
rect 24084 31736 24090 31748
rect 24121 31739 24179 31745
rect 24121 31736 24133 31739
rect 24084 31708 24133 31736
rect 24084 31696 24090 31708
rect 24121 31705 24133 31708
rect 24167 31736 24179 31739
rect 24504 31736 24532 31767
rect 24167 31708 24532 31736
rect 24596 31736 24624 31844
rect 26326 31832 26332 31884
rect 26384 31872 26390 31884
rect 26421 31875 26479 31881
rect 26421 31872 26433 31875
rect 26384 31844 26433 31872
rect 26384 31832 26390 31844
rect 26421 31841 26433 31844
rect 26467 31841 26479 31875
rect 26421 31835 26479 31841
rect 26605 31875 26663 31881
rect 26605 31841 26617 31875
rect 26651 31872 26663 31875
rect 26694 31872 26700 31884
rect 26651 31844 26700 31872
rect 26651 31841 26663 31844
rect 26605 31835 26663 31841
rect 26694 31832 26700 31844
rect 26752 31832 26758 31884
rect 29362 31832 29368 31884
rect 29420 31832 29426 31884
rect 26878 31736 26884 31748
rect 24596 31708 26884 31736
rect 24167 31705 24179 31708
rect 24121 31699 24179 31705
rect 26878 31696 26884 31708
rect 26936 31696 26942 31748
rect 8846 31628 8852 31680
rect 8904 31668 8910 31680
rect 9033 31671 9091 31677
rect 9033 31668 9045 31671
rect 8904 31640 9045 31668
rect 8904 31628 8910 31640
rect 9033 31637 9045 31640
rect 9079 31637 9091 31671
rect 9033 31631 9091 31637
rect 9306 31628 9312 31680
rect 9364 31668 9370 31680
rect 11054 31668 11060 31680
rect 9364 31640 11060 31668
rect 9364 31628 9370 31640
rect 11054 31628 11060 31640
rect 11112 31668 11118 31680
rect 12342 31668 12348 31680
rect 11112 31640 12348 31668
rect 11112 31628 11118 31640
rect 12342 31628 12348 31640
rect 12400 31628 12406 31680
rect 14458 31628 14464 31680
rect 14516 31628 14522 31680
rect 16669 31671 16727 31677
rect 16669 31637 16681 31671
rect 16715 31668 16727 31671
rect 16942 31668 16948 31680
rect 16715 31640 16948 31668
rect 16715 31637 16727 31640
rect 16669 31631 16727 31637
rect 16942 31628 16948 31640
rect 17000 31628 17006 31680
rect 17681 31671 17739 31677
rect 17681 31637 17693 31671
rect 17727 31668 17739 31671
rect 17770 31668 17776 31680
rect 17727 31640 17776 31668
rect 17727 31637 17739 31640
rect 17681 31631 17739 31637
rect 17770 31628 17776 31640
rect 17828 31628 17834 31680
rect 22370 31628 22376 31680
rect 22428 31668 22434 31680
rect 22649 31671 22707 31677
rect 22649 31668 22661 31671
rect 22428 31640 22661 31668
rect 22428 31628 22434 31640
rect 22649 31637 22661 31640
rect 22695 31668 22707 31671
rect 24673 31671 24731 31677
rect 24673 31668 24685 31671
rect 22695 31640 24685 31668
rect 22695 31637 22707 31640
rect 22649 31631 22707 31637
rect 24673 31637 24685 31640
rect 24719 31668 24731 31671
rect 25130 31668 25136 31680
rect 24719 31640 25136 31668
rect 24719 31637 24731 31640
rect 24673 31631 24731 31637
rect 25130 31628 25136 31640
rect 25188 31628 25194 31680
rect 26510 31628 26516 31680
rect 26568 31628 26574 31680
rect 552 31578 31648 31600
rect 552 31526 3662 31578
rect 3714 31526 3726 31578
rect 3778 31526 3790 31578
rect 3842 31526 3854 31578
rect 3906 31526 3918 31578
rect 3970 31526 11436 31578
rect 11488 31526 11500 31578
rect 11552 31526 11564 31578
rect 11616 31526 11628 31578
rect 11680 31526 11692 31578
rect 11744 31526 19210 31578
rect 19262 31526 19274 31578
rect 19326 31526 19338 31578
rect 19390 31526 19402 31578
rect 19454 31526 19466 31578
rect 19518 31526 26984 31578
rect 27036 31526 27048 31578
rect 27100 31526 27112 31578
rect 27164 31526 27176 31578
rect 27228 31526 27240 31578
rect 27292 31526 31648 31578
rect 552 31504 31648 31526
rect 11146 31424 11152 31476
rect 11204 31464 11210 31476
rect 11701 31467 11759 31473
rect 11701 31464 11713 31467
rect 11204 31436 11713 31464
rect 11204 31424 11210 31436
rect 11701 31433 11713 31436
rect 11747 31433 11759 31467
rect 11701 31427 11759 31433
rect 12802 31424 12808 31476
rect 12860 31464 12866 31476
rect 14921 31467 14979 31473
rect 14921 31464 14933 31467
rect 12860 31436 14933 31464
rect 12860 31424 12866 31436
rect 14921 31433 14933 31436
rect 14967 31433 14979 31467
rect 14921 31427 14979 31433
rect 20254 31424 20260 31476
rect 20312 31464 20318 31476
rect 21269 31467 21327 31473
rect 21269 31464 21281 31467
rect 20312 31436 21281 31464
rect 20312 31424 20318 31436
rect 21269 31433 21281 31436
rect 21315 31433 21327 31467
rect 21269 31427 21327 31433
rect 22186 31424 22192 31476
rect 22244 31464 22250 31476
rect 22373 31467 22431 31473
rect 22373 31464 22385 31467
rect 22244 31436 22385 31464
rect 22244 31424 22250 31436
rect 22373 31433 22385 31436
rect 22419 31433 22431 31467
rect 22373 31427 22431 31433
rect 22646 31424 22652 31476
rect 22704 31464 22710 31476
rect 24026 31464 24032 31476
rect 22704 31436 24032 31464
rect 22704 31424 22710 31436
rect 24026 31424 24032 31436
rect 24084 31464 24090 31476
rect 24084 31436 26004 31464
rect 24084 31424 24090 31436
rect 9306 31396 9312 31408
rect 9048 31368 9312 31396
rect 8938 31220 8944 31272
rect 8996 31220 9002 31272
rect 9048 31269 9076 31368
rect 9306 31356 9312 31368
rect 9364 31356 9370 31408
rect 11882 31396 11888 31408
rect 9600 31368 10088 31396
rect 9398 31328 9404 31340
rect 9140 31300 9404 31328
rect 9140 31269 9168 31300
rect 9398 31288 9404 31300
rect 9456 31288 9462 31340
rect 9033 31263 9091 31269
rect 9033 31229 9045 31263
rect 9079 31229 9091 31263
rect 9033 31223 9091 31229
rect 9125 31263 9183 31269
rect 9125 31229 9137 31263
rect 9171 31229 9183 31263
rect 9125 31223 9183 31229
rect 9309 31263 9367 31269
rect 9309 31229 9321 31263
rect 9355 31260 9367 31263
rect 9600 31260 9628 31368
rect 9355 31232 9628 31260
rect 9355 31229 9367 31232
rect 9309 31223 9367 31229
rect 9674 31220 9680 31272
rect 9732 31220 9738 31272
rect 9769 31263 9827 31269
rect 9769 31229 9781 31263
rect 9815 31229 9827 31263
rect 9769 31223 9827 31229
rect 9861 31263 9919 31269
rect 9861 31229 9873 31263
rect 9907 31260 9919 31263
rect 9950 31260 9956 31272
rect 9907 31232 9956 31260
rect 9907 31229 9919 31232
rect 9861 31223 9919 31229
rect 8662 31084 8668 31136
rect 8720 31084 8726 31136
rect 9401 31127 9459 31133
rect 9401 31093 9413 31127
rect 9447 31124 9459 31127
rect 9582 31124 9588 31136
rect 9447 31096 9588 31124
rect 9447 31093 9459 31096
rect 9401 31087 9459 31093
rect 9582 31084 9588 31096
rect 9640 31084 9646 31136
rect 9784 31124 9812 31223
rect 9950 31220 9956 31232
rect 10008 31220 10014 31272
rect 10060 31269 10088 31368
rect 10796 31368 11888 31396
rect 10796 31269 10824 31368
rect 11882 31356 11888 31368
rect 11940 31396 11946 31408
rect 12342 31396 12348 31408
rect 11940 31368 12348 31396
rect 11940 31356 11946 31368
rect 12342 31356 12348 31368
rect 12400 31356 12406 31408
rect 16850 31396 16856 31408
rect 15304 31368 16856 31396
rect 11238 31328 11244 31340
rect 10980 31300 11244 31328
rect 10980 31269 11008 31300
rect 11238 31288 11244 31300
rect 11296 31288 11302 31340
rect 13446 31328 13452 31340
rect 12176 31300 13452 31328
rect 10045 31263 10103 31269
rect 10045 31229 10057 31263
rect 10091 31260 10103 31263
rect 10781 31263 10839 31269
rect 10781 31260 10793 31263
rect 10091 31232 10793 31260
rect 10091 31229 10103 31232
rect 10045 31223 10103 31229
rect 10781 31229 10793 31232
rect 10827 31229 10839 31263
rect 10781 31223 10839 31229
rect 10965 31263 11023 31269
rect 10965 31229 10977 31263
rect 11011 31229 11023 31263
rect 10965 31223 11023 31229
rect 11054 31220 11060 31272
rect 11112 31220 11118 31272
rect 11149 31263 11207 31269
rect 11149 31229 11161 31263
rect 11195 31260 11207 31263
rect 11330 31260 11336 31272
rect 11195 31232 11336 31260
rect 11195 31229 11207 31232
rect 11149 31223 11207 31229
rect 11330 31220 11336 31232
rect 11388 31260 11394 31272
rect 11882 31260 11888 31272
rect 11388 31232 11888 31260
rect 11388 31220 11394 31232
rect 11882 31220 11888 31232
rect 11940 31220 11946 31272
rect 12176 31269 12204 31300
rect 13446 31288 13452 31300
rect 13504 31288 13510 31340
rect 15304 31337 15332 31368
rect 16850 31356 16856 31368
rect 16908 31356 16914 31408
rect 17037 31399 17095 31405
rect 17037 31365 17049 31399
rect 17083 31396 17095 31399
rect 18506 31396 18512 31408
rect 17083 31368 18512 31396
rect 17083 31365 17095 31368
rect 17037 31359 17095 31365
rect 18506 31356 18512 31368
rect 18564 31356 18570 31408
rect 20990 31356 20996 31408
rect 21048 31396 21054 31408
rect 21048 31368 21772 31396
rect 21048 31356 21054 31368
rect 15289 31331 15347 31337
rect 15289 31297 15301 31331
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 15473 31331 15531 31337
rect 15473 31297 15485 31331
rect 15519 31328 15531 31331
rect 16301 31331 16359 31337
rect 15519 31300 16252 31328
rect 15519 31297 15531 31300
rect 15473 31291 15531 31297
rect 11977 31263 12035 31269
rect 11977 31229 11989 31263
rect 12023 31229 12035 31263
rect 11977 31223 12035 31229
rect 12069 31263 12127 31269
rect 12069 31229 12081 31263
rect 12115 31229 12127 31263
rect 12069 31223 12127 31229
rect 12161 31263 12219 31269
rect 12161 31229 12173 31263
rect 12207 31229 12219 31263
rect 12161 31223 12219 31229
rect 11072 31124 11100 31220
rect 9784 31096 11100 31124
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 11425 31127 11483 31133
rect 11425 31124 11437 31127
rect 11388 31096 11437 31124
rect 11388 31084 11394 31096
rect 11425 31093 11437 31096
rect 11471 31093 11483 31127
rect 11992 31124 12020 31223
rect 12084 31192 12112 31223
rect 12342 31220 12348 31272
rect 12400 31220 12406 31272
rect 12434 31220 12440 31272
rect 12492 31260 12498 31272
rect 13814 31269 13820 31272
rect 13173 31263 13231 31269
rect 13173 31260 13185 31263
rect 12492 31232 13185 31260
rect 12492 31220 12498 31232
rect 13173 31229 13185 31232
rect 13219 31229 13231 31263
rect 13173 31223 13231 31229
rect 13265 31263 13323 31269
rect 13265 31229 13277 31263
rect 13311 31260 13323 31263
rect 13541 31263 13599 31269
rect 13541 31260 13553 31263
rect 13311 31232 13553 31260
rect 13311 31229 13323 31232
rect 13265 31223 13323 31229
rect 13541 31229 13553 31232
rect 13587 31229 13599 31263
rect 13541 31223 13599 31229
rect 13808 31223 13820 31269
rect 12802 31192 12808 31204
rect 12084 31164 12808 31192
rect 12802 31152 12808 31164
rect 12860 31152 12866 31204
rect 13188 31192 13216 31223
rect 13814 31220 13820 31223
rect 13872 31220 13878 31272
rect 15194 31220 15200 31272
rect 15252 31260 15258 31272
rect 15378 31260 15384 31272
rect 15252 31232 15384 31260
rect 15252 31220 15258 31232
rect 15378 31220 15384 31232
rect 15436 31220 15442 31272
rect 15749 31263 15807 31269
rect 15749 31229 15761 31263
rect 15795 31229 15807 31263
rect 15749 31223 15807 31229
rect 14182 31192 14188 31204
rect 13188 31164 14188 31192
rect 14182 31152 14188 31164
rect 14240 31152 14246 31204
rect 15764 31192 15792 31223
rect 15838 31220 15844 31272
rect 15896 31220 15902 31272
rect 15930 31220 15936 31272
rect 15988 31260 15994 31272
rect 16025 31263 16083 31269
rect 16025 31260 16037 31263
rect 15988 31232 16037 31260
rect 15988 31220 15994 31232
rect 16025 31229 16037 31232
rect 16071 31229 16083 31263
rect 16025 31223 16083 31229
rect 16114 31220 16120 31272
rect 16172 31220 16178 31272
rect 16224 31260 16252 31300
rect 16301 31297 16313 31331
rect 16347 31328 16359 31331
rect 17865 31331 17923 31337
rect 17865 31328 17877 31331
rect 16347 31300 17877 31328
rect 16347 31297 16359 31300
rect 16301 31291 16359 31297
rect 17865 31297 17877 31300
rect 17911 31297 17923 31331
rect 17865 31291 17923 31297
rect 21266 31288 21272 31340
rect 21324 31328 21330 31340
rect 21453 31331 21511 31337
rect 21453 31328 21465 31331
rect 21324 31300 21465 31328
rect 21324 31288 21330 31300
rect 21453 31297 21465 31300
rect 21499 31297 21511 31331
rect 21744 31328 21772 31368
rect 21818 31356 21824 31408
rect 21876 31396 21882 31408
rect 23658 31396 23664 31408
rect 21876 31368 23664 31396
rect 21876 31356 21882 31368
rect 21910 31328 21916 31340
rect 21744 31300 21916 31328
rect 21453 31291 21511 31297
rect 21910 31288 21916 31300
rect 21968 31288 21974 31340
rect 22097 31331 22155 31337
rect 22097 31297 22109 31331
rect 22143 31328 22155 31331
rect 22278 31328 22284 31340
rect 22143 31300 22284 31328
rect 22143 31297 22155 31300
rect 22097 31291 22155 31297
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 22848 31328 22876 31368
rect 23658 31356 23664 31368
rect 23716 31396 23722 31408
rect 24118 31396 24124 31408
rect 23716 31368 24124 31396
rect 23716 31356 23722 31368
rect 24118 31356 24124 31368
rect 24176 31356 24182 31408
rect 25976 31337 26004 31436
rect 22756 31300 22876 31328
rect 23569 31331 23627 31337
rect 16574 31260 16580 31272
rect 16224 31232 16580 31260
rect 16574 31220 16580 31232
rect 16632 31220 16638 31272
rect 16850 31220 16856 31272
rect 16908 31260 16914 31272
rect 17494 31260 17500 31272
rect 16908 31232 17500 31260
rect 16908 31220 16914 31232
rect 17494 31220 17500 31232
rect 17552 31220 17558 31272
rect 17589 31263 17647 31269
rect 17589 31229 17601 31263
rect 17635 31229 17647 31263
rect 17589 31223 17647 31229
rect 17034 31192 17040 31204
rect 15764 31164 17040 31192
rect 17034 31152 17040 31164
rect 17092 31152 17098 31204
rect 17313 31195 17371 31201
rect 17313 31161 17325 31195
rect 17359 31161 17371 31195
rect 17604 31192 17632 31223
rect 17770 31220 17776 31272
rect 17828 31220 17834 31272
rect 17954 31220 17960 31272
rect 18012 31220 18018 31272
rect 18141 31263 18199 31269
rect 18141 31229 18153 31263
rect 18187 31229 18199 31263
rect 18141 31223 18199 31229
rect 18046 31192 18052 31204
rect 17604 31164 18052 31192
rect 17313 31155 17371 31161
rect 13078 31124 13084 31136
rect 11992 31096 13084 31124
rect 11425 31087 11483 31093
rect 13078 31084 13084 31096
rect 13136 31084 13142 31136
rect 15657 31127 15715 31133
rect 15657 31093 15669 31127
rect 15703 31124 15715 31127
rect 15746 31124 15752 31136
rect 15703 31096 15752 31124
rect 15703 31093 15715 31096
rect 15657 31087 15715 31093
rect 15746 31084 15752 31096
rect 15804 31124 15810 31136
rect 16482 31124 16488 31136
rect 15804 31096 16488 31124
rect 15804 31084 15810 31096
rect 16482 31084 16488 31096
rect 16540 31084 16546 31136
rect 16850 31084 16856 31136
rect 16908 31084 16914 31136
rect 17328 31124 17356 31155
rect 18046 31152 18052 31164
rect 18104 31152 18110 31204
rect 18156 31124 18184 31223
rect 18690 31220 18696 31272
rect 18748 31220 18754 31272
rect 20806 31220 20812 31272
rect 20864 31220 20870 31272
rect 20990 31220 20996 31272
rect 21048 31220 21054 31272
rect 21358 31220 21364 31272
rect 21416 31220 21422 31272
rect 21637 31263 21695 31269
rect 21637 31229 21649 31263
rect 21683 31229 21695 31263
rect 21637 31223 21695 31229
rect 21729 31263 21787 31269
rect 21729 31229 21741 31263
rect 21775 31260 21787 31263
rect 22370 31260 22376 31272
rect 21775 31232 22376 31260
rect 21775 31229 21787 31232
rect 21729 31223 21787 31229
rect 18325 31195 18383 31201
rect 18325 31161 18337 31195
rect 18371 31192 18383 31195
rect 18938 31195 18996 31201
rect 18938 31192 18950 31195
rect 18371 31164 18950 31192
rect 18371 31161 18383 31164
rect 18325 31155 18383 31161
rect 18938 31161 18950 31164
rect 18984 31161 18996 31195
rect 18938 31155 18996 31161
rect 21085 31195 21143 31201
rect 21085 31161 21097 31195
rect 21131 31192 21143 31195
rect 21652 31192 21680 31223
rect 22370 31220 22376 31232
rect 22428 31220 22434 31272
rect 22554 31220 22560 31272
rect 22612 31220 22618 31272
rect 22756 31269 22784 31300
rect 23569 31297 23581 31331
rect 23615 31328 23627 31331
rect 24213 31331 24271 31337
rect 24213 31328 24225 31331
rect 23615 31300 24225 31328
rect 23615 31297 23627 31300
rect 23569 31291 23627 31297
rect 24213 31297 24225 31300
rect 24259 31297 24271 31331
rect 24213 31291 24271 31297
rect 25961 31331 26019 31337
rect 25961 31297 25973 31331
rect 26007 31297 26019 31331
rect 25961 31291 26019 31297
rect 26418 31288 26424 31340
rect 26476 31288 26482 31340
rect 22741 31263 22799 31269
rect 22741 31229 22753 31263
rect 22787 31229 22799 31263
rect 22741 31223 22799 31229
rect 23014 31220 23020 31272
rect 23072 31220 23078 31272
rect 23474 31220 23480 31272
rect 23532 31260 23538 31272
rect 23937 31263 23995 31269
rect 23937 31260 23949 31263
rect 23532 31232 23949 31260
rect 23532 31220 23538 31232
rect 23937 31229 23949 31232
rect 23983 31229 23995 31263
rect 23937 31223 23995 31229
rect 26050 31220 26056 31272
rect 26108 31220 26114 31272
rect 26878 31220 26884 31272
rect 26936 31260 26942 31272
rect 27341 31263 27399 31269
rect 27341 31260 27353 31263
rect 26936 31232 27353 31260
rect 26936 31220 26942 31232
rect 27341 31229 27353 31232
rect 27387 31260 27399 31263
rect 27433 31263 27491 31269
rect 27433 31260 27445 31263
rect 27387 31232 27445 31260
rect 27387 31229 27399 31232
rect 27341 31223 27399 31229
rect 27433 31229 27445 31232
rect 27479 31229 27491 31263
rect 27433 31223 27491 31229
rect 27617 31263 27675 31269
rect 27617 31229 27629 31263
rect 27663 31260 27675 31263
rect 27982 31260 27988 31272
rect 27663 31232 27988 31260
rect 27663 31229 27675 31232
rect 27617 31223 27675 31229
rect 21131 31164 21680 31192
rect 21131 31161 21143 31164
rect 21085 31155 21143 31161
rect 18414 31124 18420 31136
rect 17328 31096 18420 31124
rect 18414 31084 18420 31096
rect 18472 31124 18478 31136
rect 20073 31127 20131 31133
rect 20073 31124 20085 31127
rect 18472 31096 20085 31124
rect 18472 31084 18478 31096
rect 20073 31093 20085 31096
rect 20119 31093 20131 31127
rect 21652 31124 21680 31164
rect 21818 31152 21824 31204
rect 21876 31152 21882 31204
rect 21910 31152 21916 31204
rect 21968 31201 21974 31204
rect 21968 31195 21997 31201
rect 21985 31192 21997 31195
rect 21985 31164 22600 31192
rect 21985 31161 21997 31164
rect 21968 31155 21997 31161
rect 21968 31152 21974 31155
rect 22462 31124 22468 31136
rect 21652 31096 22468 31124
rect 20073 31087 20131 31093
rect 22462 31084 22468 31096
rect 22520 31084 22526 31136
rect 22572 31124 22600 31164
rect 22646 31152 22652 31204
rect 22704 31152 22710 31204
rect 22879 31195 22937 31201
rect 22879 31192 22891 31195
rect 22756 31164 22891 31192
rect 22756 31124 22784 31164
rect 22879 31161 22891 31164
rect 22925 31161 22937 31195
rect 22879 31155 22937 31161
rect 23658 31152 23664 31204
rect 23716 31192 23722 31204
rect 24458 31195 24516 31201
rect 24458 31192 24470 31195
rect 23716 31164 24470 31192
rect 23716 31152 23722 31164
rect 24458 31161 24470 31164
rect 24504 31161 24516 31195
rect 24458 31155 24516 31161
rect 26513 31195 26571 31201
rect 26513 31161 26525 31195
rect 26559 31161 26571 31195
rect 26513 31155 26571 31161
rect 23106 31124 23112 31136
rect 22572 31096 23112 31124
rect 23106 31084 23112 31096
rect 23164 31084 23170 31136
rect 24029 31127 24087 31133
rect 24029 31093 24041 31127
rect 24075 31124 24087 31127
rect 24210 31124 24216 31136
rect 24075 31096 24216 31124
rect 24075 31093 24087 31096
rect 24029 31087 24087 31093
rect 24210 31084 24216 31096
rect 24268 31084 24274 31136
rect 24946 31084 24952 31136
rect 25004 31124 25010 31136
rect 25593 31127 25651 31133
rect 25593 31124 25605 31127
rect 25004 31096 25605 31124
rect 25004 31084 25010 31096
rect 25593 31093 25605 31096
rect 25639 31124 25651 31127
rect 26326 31124 26332 31136
rect 25639 31096 26332 31124
rect 25639 31093 25651 31096
rect 25593 31087 25651 31093
rect 26326 31084 26332 31096
rect 26384 31124 26390 31136
rect 26528 31124 26556 31155
rect 26694 31152 26700 31204
rect 26752 31152 26758 31204
rect 27157 31195 27215 31201
rect 27157 31161 27169 31195
rect 27203 31192 27215 31195
rect 27632 31192 27660 31223
rect 27982 31220 27988 31232
rect 28040 31220 28046 31272
rect 27203 31164 27660 31192
rect 27203 31161 27215 31164
rect 27157 31155 27215 31161
rect 26384 31096 26556 31124
rect 26384 31084 26390 31096
rect 26878 31084 26884 31136
rect 26936 31084 26942 31136
rect 26970 31084 26976 31136
rect 27028 31084 27034 31136
rect 27522 31084 27528 31136
rect 27580 31084 27586 31136
rect 552 31034 31648 31056
rect 552 30982 4322 31034
rect 4374 30982 4386 31034
rect 4438 30982 4450 31034
rect 4502 30982 4514 31034
rect 4566 30982 4578 31034
rect 4630 30982 12096 31034
rect 12148 30982 12160 31034
rect 12212 30982 12224 31034
rect 12276 30982 12288 31034
rect 12340 30982 12352 31034
rect 12404 30982 19870 31034
rect 19922 30982 19934 31034
rect 19986 30982 19998 31034
rect 20050 30982 20062 31034
rect 20114 30982 20126 31034
rect 20178 30982 27644 31034
rect 27696 30982 27708 31034
rect 27760 30982 27772 31034
rect 27824 30982 27836 31034
rect 27888 30982 27900 31034
rect 27952 30982 31648 31034
rect 552 30960 31648 30982
rect 8938 30880 8944 30932
rect 8996 30920 9002 30932
rect 10229 30923 10287 30929
rect 10229 30920 10241 30923
rect 8996 30892 10241 30920
rect 8996 30880 9002 30892
rect 10229 30889 10241 30892
rect 10275 30920 10287 30923
rect 10318 30920 10324 30932
rect 10275 30892 10324 30920
rect 10275 30889 10287 30892
rect 10229 30883 10287 30889
rect 10318 30880 10324 30892
rect 10376 30880 10382 30932
rect 11606 30880 11612 30932
rect 11664 30920 11670 30932
rect 12710 30920 12716 30932
rect 11664 30892 12716 30920
rect 11664 30880 11670 30892
rect 12710 30880 12716 30892
rect 12768 30880 12774 30932
rect 12802 30880 12808 30932
rect 12860 30880 12866 30932
rect 13446 30880 13452 30932
rect 13504 30920 13510 30932
rect 13541 30923 13599 30929
rect 13541 30920 13553 30923
rect 13504 30892 13553 30920
rect 13504 30880 13510 30892
rect 13541 30889 13553 30892
rect 13587 30889 13599 30923
rect 13541 30883 13599 30889
rect 15838 30880 15844 30932
rect 15896 30880 15902 30932
rect 16209 30923 16267 30929
rect 16209 30889 16221 30923
rect 16255 30920 16267 30923
rect 16298 30920 16304 30932
rect 16255 30892 16304 30920
rect 16255 30889 16267 30892
rect 16209 30883 16267 30889
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 17862 30920 17868 30932
rect 16500 30892 17868 30920
rect 8662 30812 8668 30864
rect 8720 30852 8726 30864
rect 9094 30855 9152 30861
rect 9094 30852 9106 30855
rect 8720 30824 9106 30852
rect 8720 30812 8726 30824
rect 9094 30821 9106 30824
rect 9140 30821 9152 30855
rect 13909 30855 13967 30861
rect 9094 30815 9152 30821
rect 13280 30824 13860 30852
rect 13280 30796 13308 30824
rect 8846 30744 8852 30796
rect 8904 30744 8910 30796
rect 10042 30744 10048 30796
rect 10100 30784 10106 30796
rect 11149 30787 11207 30793
rect 11149 30784 11161 30787
rect 10100 30756 11161 30784
rect 10100 30744 10106 30756
rect 11149 30753 11161 30756
rect 11195 30753 11207 30787
rect 11149 30747 11207 30753
rect 11882 30744 11888 30796
rect 11940 30744 11946 30796
rect 13078 30744 13084 30796
rect 13136 30784 13142 30796
rect 13262 30784 13268 30796
rect 13136 30756 13268 30784
rect 13136 30744 13142 30756
rect 13262 30744 13268 30756
rect 13320 30744 13326 30796
rect 13357 30787 13415 30793
rect 13357 30753 13369 30787
rect 13403 30784 13415 30787
rect 13725 30787 13783 30793
rect 13725 30784 13737 30787
rect 13403 30756 13737 30784
rect 13403 30753 13415 30756
rect 13357 30747 13415 30753
rect 13725 30753 13737 30756
rect 13771 30753 13783 30787
rect 13832 30784 13860 30824
rect 13909 30821 13921 30855
rect 13955 30852 13967 30855
rect 14458 30852 14464 30864
rect 13955 30824 14464 30852
rect 13955 30821 13967 30824
rect 13909 30815 13967 30821
rect 14458 30812 14464 30824
rect 14516 30812 14522 30864
rect 15286 30812 15292 30864
rect 15344 30852 15350 30864
rect 15381 30855 15439 30861
rect 15381 30852 15393 30855
rect 15344 30824 15393 30852
rect 15344 30812 15350 30824
rect 15381 30821 15393 30824
rect 15427 30852 15439 30855
rect 16500 30852 16528 30892
rect 17862 30880 17868 30892
rect 17920 30880 17926 30932
rect 18138 30880 18144 30932
rect 18196 30920 18202 30932
rect 18233 30923 18291 30929
rect 18233 30920 18245 30923
rect 18196 30892 18245 30920
rect 18196 30880 18202 30892
rect 18233 30889 18245 30892
rect 18279 30889 18291 30923
rect 18233 30883 18291 30889
rect 18690 30880 18696 30932
rect 18748 30920 18754 30932
rect 19061 30923 19119 30929
rect 19061 30920 19073 30923
rect 18748 30892 19073 30920
rect 18748 30880 18754 30892
rect 19061 30889 19073 30892
rect 19107 30889 19119 30923
rect 19061 30883 19119 30889
rect 23658 30880 23664 30932
rect 23716 30880 23722 30932
rect 26050 30880 26056 30932
rect 26108 30920 26114 30932
rect 26326 30920 26332 30932
rect 26108 30892 26332 30920
rect 26108 30880 26114 30892
rect 26326 30880 26332 30892
rect 26384 30880 26390 30932
rect 26878 30920 26884 30932
rect 26712 30892 26884 30920
rect 15427 30824 16528 30852
rect 15427 30821 15439 30824
rect 15381 30815 15439 30821
rect 16574 30812 16580 30864
rect 16632 30852 16638 30864
rect 26712 30861 26740 30892
rect 26878 30880 26884 30892
rect 26936 30880 26942 30932
rect 26970 30880 26976 30932
rect 27028 30880 27034 30932
rect 24121 30855 24179 30861
rect 16632 30824 17172 30852
rect 16632 30812 16638 30824
rect 14185 30787 14243 30793
rect 14185 30784 14197 30787
rect 13832 30756 14197 30784
rect 13725 30747 13783 30753
rect 14185 30753 14197 30756
rect 14231 30753 14243 30787
rect 14185 30747 14243 30753
rect 14550 30744 14556 30796
rect 14608 30744 14614 30796
rect 14921 30787 14979 30793
rect 14921 30784 14933 30787
rect 14660 30756 14933 30784
rect 10318 30676 10324 30728
rect 10376 30716 10382 30728
rect 10965 30719 11023 30725
rect 10965 30716 10977 30719
rect 10376 30688 10977 30716
rect 10376 30676 10382 30688
rect 10965 30685 10977 30688
rect 11011 30685 11023 30719
rect 10965 30679 11023 30685
rect 11606 30676 11612 30728
rect 11664 30676 11670 30728
rect 12066 30725 12072 30728
rect 12023 30719 12072 30725
rect 12023 30685 12035 30719
rect 12069 30685 12072 30719
rect 12023 30679 12072 30685
rect 12066 30676 12072 30679
rect 12124 30676 12130 30728
rect 12158 30676 12164 30728
rect 12216 30716 12222 30728
rect 14568 30716 14596 30744
rect 12216 30688 14596 30716
rect 12216 30676 12222 30688
rect 12710 30608 12716 30660
rect 12768 30648 12774 30660
rect 14182 30648 14188 30660
rect 12768 30620 14188 30648
rect 12768 30608 12774 30620
rect 14182 30608 14188 30620
rect 14240 30648 14246 30660
rect 14660 30648 14688 30756
rect 14921 30753 14933 30756
rect 14967 30753 14979 30787
rect 14921 30747 14979 30753
rect 15562 30744 15568 30796
rect 15620 30784 15626 30796
rect 15749 30787 15807 30793
rect 15749 30784 15761 30787
rect 15620 30756 15761 30784
rect 15620 30744 15626 30756
rect 15749 30753 15761 30756
rect 15795 30753 15807 30787
rect 15749 30747 15807 30753
rect 16482 30744 16488 30796
rect 16540 30744 16546 30796
rect 16761 30787 16819 30793
rect 16761 30753 16773 30787
rect 16807 30753 16819 30787
rect 16761 30747 16819 30753
rect 16776 30716 16804 30747
rect 16850 30744 16856 30796
rect 16908 30784 16914 30796
rect 16945 30787 17003 30793
rect 16945 30784 16957 30787
rect 16908 30756 16957 30784
rect 16908 30744 16914 30756
rect 16945 30753 16957 30756
rect 16991 30753 17003 30787
rect 17144 30784 17172 30824
rect 23308 30824 23796 30852
rect 17144 30756 17264 30784
rect 16945 30747 17003 30753
rect 17126 30716 17132 30728
rect 16776 30688 17132 30716
rect 17126 30676 17132 30688
rect 17184 30676 17190 30728
rect 14240 30620 14688 30648
rect 14240 30608 14246 30620
rect 16298 30608 16304 30660
rect 16356 30648 16362 30660
rect 17236 30657 17264 30756
rect 18506 30744 18512 30796
rect 18564 30784 18570 30796
rect 18785 30787 18843 30793
rect 18785 30784 18797 30787
rect 18564 30756 18797 30784
rect 18564 30744 18570 30756
rect 18785 30753 18797 30756
rect 18831 30753 18843 30787
rect 18785 30747 18843 30753
rect 19058 30744 19064 30796
rect 19116 30784 19122 30796
rect 19153 30787 19211 30793
rect 19153 30784 19165 30787
rect 19116 30756 19165 30784
rect 19116 30744 19122 30756
rect 19153 30753 19165 30756
rect 19199 30753 19211 30787
rect 19153 30747 19211 30753
rect 22002 30744 22008 30796
rect 22060 30784 22066 30796
rect 22370 30784 22376 30796
rect 22060 30756 22376 30784
rect 22060 30744 22066 30756
rect 22370 30744 22376 30756
rect 22428 30784 22434 30796
rect 23308 30793 23336 30824
rect 23768 30793 23796 30824
rect 24121 30821 24133 30855
rect 24167 30852 24179 30855
rect 24458 30855 24516 30861
rect 24458 30852 24470 30855
rect 24167 30824 24470 30852
rect 24167 30821 24179 30824
rect 24121 30815 24179 30821
rect 24458 30821 24470 30824
rect 24504 30821 24516 30855
rect 24458 30815 24516 30821
rect 26697 30855 26755 30861
rect 26697 30821 26709 30855
rect 26743 30821 26755 30855
rect 26697 30815 26755 30821
rect 26789 30855 26847 30861
rect 26789 30821 26801 30855
rect 26835 30852 26847 30855
rect 26988 30852 27016 30880
rect 26835 30824 27016 30852
rect 26835 30821 26847 30824
rect 26789 30815 26847 30821
rect 27430 30812 27436 30864
rect 27488 30852 27494 30864
rect 28077 30855 28135 30861
rect 28077 30852 28089 30855
rect 27488 30824 28089 30852
rect 27488 30812 27494 30824
rect 28077 30821 28089 30824
rect 28123 30852 28135 30855
rect 28442 30852 28448 30864
rect 28123 30824 28448 30852
rect 28123 30821 28135 30824
rect 28077 30815 28135 30821
rect 28442 30812 28448 30824
rect 28500 30812 28506 30864
rect 23293 30787 23351 30793
rect 23293 30784 23305 30787
rect 22428 30756 23305 30784
rect 22428 30744 22434 30756
rect 23293 30753 23305 30756
rect 23339 30753 23351 30787
rect 23293 30747 23351 30753
rect 23477 30787 23535 30793
rect 23477 30753 23489 30787
rect 23523 30753 23535 30787
rect 23477 30747 23535 30753
rect 23753 30787 23811 30793
rect 23753 30753 23765 30787
rect 23799 30753 23811 30787
rect 23753 30747 23811 30753
rect 17589 30719 17647 30725
rect 17589 30716 17601 30719
rect 17328 30688 17601 30716
rect 17221 30651 17279 30657
rect 16356 30620 17080 30648
rect 16356 30608 16362 30620
rect 11882 30540 11888 30592
rect 11940 30580 11946 30592
rect 12526 30580 12532 30592
rect 11940 30552 12532 30580
rect 11940 30540 11946 30552
rect 12526 30540 12532 30552
rect 12584 30540 12590 30592
rect 16390 30540 16396 30592
rect 16448 30580 16454 30592
rect 16577 30583 16635 30589
rect 16577 30580 16589 30583
rect 16448 30552 16589 30580
rect 16448 30540 16454 30552
rect 16577 30549 16589 30552
rect 16623 30549 16635 30583
rect 16577 30543 16635 30549
rect 16666 30540 16672 30592
rect 16724 30540 16730 30592
rect 17052 30580 17080 30620
rect 17221 30617 17233 30651
rect 17267 30617 17279 30651
rect 17221 30611 17279 30617
rect 17328 30580 17356 30688
rect 17589 30685 17601 30688
rect 17635 30685 17647 30719
rect 17589 30679 17647 30685
rect 17052 30552 17356 30580
rect 23492 30580 23520 30747
rect 23934 30744 23940 30796
rect 23992 30744 23998 30796
rect 24210 30744 24216 30796
rect 24268 30744 24274 30796
rect 26418 30744 26424 30796
rect 26476 30744 26482 30796
rect 26510 30744 26516 30796
rect 26568 30784 26574 30796
rect 26927 30787 26985 30793
rect 26568 30756 26613 30784
rect 26568 30744 26574 30756
rect 26927 30753 26939 30787
rect 26973 30784 26985 30787
rect 27522 30784 27528 30796
rect 26973 30756 27528 30784
rect 26973 30753 26985 30756
rect 26927 30747 26985 30753
rect 27522 30744 27528 30756
rect 27580 30744 27586 30796
rect 27893 30787 27951 30793
rect 27893 30753 27905 30787
rect 27939 30784 27951 30787
rect 27982 30784 27988 30796
rect 27939 30756 27988 30784
rect 27939 30753 27951 30756
rect 27893 30747 27951 30753
rect 27982 30744 27988 30756
rect 28040 30784 28046 30796
rect 28902 30784 28908 30796
rect 28040 30756 28908 30784
rect 28040 30744 28046 30756
rect 28902 30744 28908 30756
rect 28960 30744 28966 30796
rect 25222 30580 25228 30592
rect 23492 30552 25228 30580
rect 25222 30540 25228 30552
rect 25280 30540 25286 30592
rect 25590 30540 25596 30592
rect 25648 30540 25654 30592
rect 26694 30540 26700 30592
rect 26752 30580 26758 30592
rect 27065 30583 27123 30589
rect 27065 30580 27077 30583
rect 26752 30552 27077 30580
rect 26752 30540 26758 30552
rect 27065 30549 27077 30552
rect 27111 30549 27123 30583
rect 27065 30543 27123 30549
rect 27709 30583 27767 30589
rect 27709 30549 27721 30583
rect 27755 30580 27767 30583
rect 27982 30580 27988 30592
rect 27755 30552 27988 30580
rect 27755 30549 27767 30552
rect 27709 30543 27767 30549
rect 27982 30540 27988 30552
rect 28040 30540 28046 30592
rect 552 30490 31648 30512
rect 552 30438 3662 30490
rect 3714 30438 3726 30490
rect 3778 30438 3790 30490
rect 3842 30438 3854 30490
rect 3906 30438 3918 30490
rect 3970 30438 11436 30490
rect 11488 30438 11500 30490
rect 11552 30438 11564 30490
rect 11616 30438 11628 30490
rect 11680 30438 11692 30490
rect 11744 30438 19210 30490
rect 19262 30438 19274 30490
rect 19326 30438 19338 30490
rect 19390 30438 19402 30490
rect 19454 30438 19466 30490
rect 19518 30438 26984 30490
rect 27036 30438 27048 30490
rect 27100 30438 27112 30490
rect 27164 30438 27176 30490
rect 27228 30438 27240 30490
rect 27292 30438 31648 30490
rect 552 30416 31648 30438
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 10689 30379 10747 30385
rect 10689 30376 10701 30379
rect 9732 30348 10701 30376
rect 9732 30336 9738 30348
rect 10689 30345 10701 30348
rect 10735 30376 10747 30379
rect 12066 30376 12072 30388
rect 10735 30348 12072 30376
rect 10735 30345 10747 30348
rect 10689 30339 10747 30345
rect 12066 30336 12072 30348
rect 12124 30336 12130 30388
rect 15562 30336 15568 30388
rect 15620 30336 15626 30388
rect 15933 30379 15991 30385
rect 15933 30345 15945 30379
rect 15979 30376 15991 30379
rect 15979 30348 16344 30376
rect 15979 30345 15991 30348
rect 15933 30339 15991 30345
rect 12437 30311 12495 30317
rect 12437 30277 12449 30311
rect 12483 30308 12495 30311
rect 12526 30308 12532 30320
rect 12483 30280 12532 30308
rect 12483 30277 12495 30280
rect 12437 30271 12495 30277
rect 12526 30268 12532 30280
rect 12584 30268 12590 30320
rect 16206 30268 16212 30320
rect 16264 30268 16270 30320
rect 15378 30200 15384 30252
rect 15436 30240 15442 30252
rect 15841 30243 15899 30249
rect 15841 30240 15853 30243
rect 15436 30212 15853 30240
rect 15436 30200 15442 30212
rect 15841 30209 15853 30212
rect 15887 30240 15899 30243
rect 16316 30240 16344 30348
rect 16666 30336 16672 30388
rect 16724 30336 16730 30388
rect 23014 30336 23020 30388
rect 23072 30376 23078 30388
rect 23845 30379 23903 30385
rect 23072 30348 23520 30376
rect 23072 30336 23078 30348
rect 16482 30268 16488 30320
rect 16540 30308 16546 30320
rect 16577 30311 16635 30317
rect 16577 30308 16589 30311
rect 16540 30280 16589 30308
rect 16540 30268 16546 30280
rect 16577 30277 16589 30280
rect 16623 30277 16635 30311
rect 16577 30271 16635 30277
rect 16684 30240 16712 30336
rect 17034 30268 17040 30320
rect 17092 30268 17098 30320
rect 23492 30308 23520 30348
rect 23845 30345 23857 30379
rect 23891 30376 23903 30379
rect 23934 30376 23940 30388
rect 23891 30348 23940 30376
rect 23891 30345 23903 30348
rect 23845 30339 23903 30345
rect 23934 30336 23940 30348
rect 23992 30336 23998 30388
rect 24118 30336 24124 30388
rect 24176 30376 24182 30388
rect 24854 30376 24860 30388
rect 24176 30348 24860 30376
rect 24176 30336 24182 30348
rect 24854 30336 24860 30348
rect 24912 30336 24918 30388
rect 23492 30280 24624 30308
rect 17773 30243 17831 30249
rect 17773 30240 17785 30243
rect 15887 30212 16252 30240
rect 16316 30212 16620 30240
rect 16684 30212 17785 30240
rect 15887 30209 15899 30212
rect 15841 30203 15899 30209
rect 16224 30184 16252 30212
rect 16592 30184 16620 30212
rect 9030 30132 9036 30184
rect 9088 30132 9094 30184
rect 11330 30181 11336 30184
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30172 9183 30175
rect 9309 30175 9367 30181
rect 9309 30172 9321 30175
rect 9171 30144 9321 30172
rect 9171 30141 9183 30144
rect 9125 30135 9183 30141
rect 9309 30141 9321 30144
rect 9355 30141 9367 30175
rect 10781 30175 10839 30181
rect 10781 30172 10793 30175
rect 9309 30135 9367 30141
rect 9508 30144 10793 30172
rect 9048 30104 9076 30132
rect 9398 30104 9404 30116
rect 9048 30076 9404 30104
rect 9398 30064 9404 30076
rect 9456 30104 9462 30116
rect 9508 30104 9536 30144
rect 10781 30141 10793 30144
rect 10827 30141 10839 30175
rect 10781 30135 10839 30141
rect 10873 30175 10931 30181
rect 10873 30141 10885 30175
rect 10919 30172 10931 30175
rect 11057 30175 11115 30181
rect 11057 30172 11069 30175
rect 10919 30144 11069 30172
rect 10919 30141 10931 30144
rect 10873 30135 10931 30141
rect 11057 30141 11069 30144
rect 11103 30141 11115 30175
rect 11324 30172 11336 30181
rect 11291 30144 11336 30172
rect 11057 30135 11115 30141
rect 11324 30135 11336 30144
rect 11330 30132 11336 30135
rect 11388 30132 11394 30184
rect 14274 30132 14280 30184
rect 14332 30172 14338 30184
rect 14369 30175 14427 30181
rect 14369 30172 14381 30175
rect 14332 30144 14381 30172
rect 14332 30132 14338 30144
rect 14369 30141 14381 30144
rect 14415 30141 14427 30175
rect 14369 30135 14427 30141
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30141 15991 30175
rect 15933 30135 15991 30141
rect 9582 30113 9588 30116
rect 9456 30076 9536 30104
rect 9456 30064 9462 30076
rect 9576 30067 9588 30113
rect 9640 30104 9646 30116
rect 15948 30104 15976 30135
rect 16206 30132 16212 30184
rect 16264 30132 16270 30184
rect 16390 30132 16396 30184
rect 16448 30172 16454 30184
rect 16485 30175 16543 30181
rect 16485 30172 16497 30175
rect 16448 30144 16497 30172
rect 16448 30132 16454 30144
rect 16485 30141 16497 30144
rect 16531 30141 16543 30175
rect 16485 30135 16543 30141
rect 16574 30132 16580 30184
rect 16632 30132 16638 30184
rect 16666 30132 16672 30184
rect 16724 30172 16730 30184
rect 16761 30175 16819 30181
rect 16761 30172 16773 30175
rect 16724 30144 16773 30172
rect 16724 30132 16730 30144
rect 16761 30141 16773 30144
rect 16807 30141 16819 30175
rect 16761 30135 16819 30141
rect 16945 30175 17003 30181
rect 16945 30141 16957 30175
rect 16991 30141 17003 30175
rect 16945 30135 17003 30141
rect 16850 30104 16856 30116
rect 9640 30076 9676 30104
rect 15948 30076 16856 30104
rect 9582 30064 9588 30067
rect 9640 30064 9646 30076
rect 16850 30064 16856 30076
rect 16908 30064 16914 30116
rect 14090 29996 14096 30048
rect 14148 30036 14154 30048
rect 14277 30039 14335 30045
rect 14277 30036 14289 30039
rect 14148 30008 14289 30036
rect 14148 29996 14154 30008
rect 14277 30005 14289 30008
rect 14323 30005 14335 30039
rect 14277 29999 14335 30005
rect 16114 29996 16120 30048
rect 16172 30036 16178 30048
rect 16298 30036 16304 30048
rect 16172 30008 16304 30036
rect 16172 29996 16178 30008
rect 16298 29996 16304 30008
rect 16356 30036 16362 30048
rect 16960 30036 16988 30135
rect 17218 30132 17224 30184
rect 17276 30132 17282 30184
rect 17512 30181 17540 30212
rect 17773 30209 17785 30212
rect 17819 30209 17831 30243
rect 17773 30203 17831 30209
rect 23198 30200 23204 30252
rect 23256 30240 23262 30252
rect 23842 30240 23848 30252
rect 23256 30212 23848 30240
rect 23256 30200 23262 30212
rect 23842 30200 23848 30212
rect 23900 30240 23906 30252
rect 24596 30249 24624 30280
rect 25222 30268 25228 30320
rect 25280 30268 25286 30320
rect 24489 30243 24547 30249
rect 24489 30240 24501 30243
rect 23900 30212 24501 30240
rect 23900 30200 23906 30212
rect 24489 30209 24501 30212
rect 24535 30209 24547 30243
rect 24489 30203 24547 30209
rect 24581 30243 24639 30249
rect 24581 30209 24593 30243
rect 24627 30209 24639 30243
rect 24581 30203 24639 30209
rect 24780 30212 25084 30240
rect 17313 30175 17371 30181
rect 17313 30141 17325 30175
rect 17359 30141 17371 30175
rect 17313 30135 17371 30141
rect 17497 30175 17555 30181
rect 17497 30141 17509 30175
rect 17543 30141 17555 30175
rect 17497 30135 17555 30141
rect 17328 30104 17356 30135
rect 17586 30132 17592 30184
rect 17644 30132 17650 30184
rect 17862 30132 17868 30184
rect 17920 30132 17926 30184
rect 19058 30132 19064 30184
rect 19116 30172 19122 30184
rect 19245 30175 19303 30181
rect 19245 30172 19257 30175
rect 19116 30144 19257 30172
rect 19116 30132 19122 30144
rect 19245 30141 19257 30144
rect 19291 30141 19303 30175
rect 19245 30135 19303 30141
rect 22002 30132 22008 30184
rect 22060 30172 22066 30184
rect 23934 30172 23940 30184
rect 22060 30144 23940 30172
rect 22060 30132 22066 30144
rect 23934 30132 23940 30144
rect 23992 30172 23998 30184
rect 24029 30175 24087 30181
rect 24029 30172 24041 30175
rect 23992 30144 24041 30172
rect 23992 30132 23998 30144
rect 24029 30141 24041 30144
rect 24075 30172 24087 30175
rect 24780 30172 24808 30212
rect 24075 30144 24808 30172
rect 24075 30141 24087 30144
rect 24029 30135 24087 30141
rect 24854 30132 24860 30184
rect 24912 30132 24918 30184
rect 25056 30181 25084 30212
rect 25041 30175 25099 30181
rect 25041 30141 25053 30175
rect 25087 30141 25099 30175
rect 25041 30135 25099 30141
rect 27157 30175 27215 30181
rect 27157 30141 27169 30175
rect 27203 30141 27215 30175
rect 27157 30135 27215 30141
rect 27249 30175 27307 30181
rect 27249 30141 27261 30175
rect 27295 30172 27307 30175
rect 27433 30175 27491 30181
rect 27433 30172 27445 30175
rect 27295 30144 27445 30172
rect 27295 30141 27307 30144
rect 27249 30135 27307 30141
rect 27433 30141 27445 30144
rect 27479 30141 27491 30175
rect 27433 30135 27491 30141
rect 18506 30104 18512 30116
rect 17328 30076 18512 30104
rect 18506 30064 18512 30076
rect 18564 30064 18570 30116
rect 24121 30107 24179 30113
rect 24121 30073 24133 30107
rect 24167 30073 24179 30107
rect 24121 30067 24179 30073
rect 16356 30008 16988 30036
rect 16356 29996 16362 30008
rect 18966 29996 18972 30048
rect 19024 30036 19030 30048
rect 19153 30039 19211 30045
rect 19153 30036 19165 30039
rect 19024 30008 19165 30036
rect 19024 29996 19030 30008
rect 19153 30005 19165 30008
rect 19199 30005 19211 30039
rect 24136 30036 24164 30067
rect 24210 30064 24216 30116
rect 24268 30064 24274 30116
rect 24302 30064 24308 30116
rect 24360 30113 24366 30116
rect 24360 30107 24389 30113
rect 24377 30104 24389 30107
rect 24719 30107 24777 30113
rect 24719 30104 24731 30107
rect 24377 30076 24731 30104
rect 24377 30073 24389 30076
rect 24360 30067 24389 30073
rect 24719 30073 24731 30076
rect 24765 30073 24777 30107
rect 24719 30067 24777 30073
rect 24360 30064 24366 30067
rect 24946 30064 24952 30116
rect 25004 30064 25010 30116
rect 27172 30104 27200 30135
rect 27338 30104 27344 30116
rect 27172 30076 27344 30104
rect 27338 30064 27344 30076
rect 27396 30064 27402 30116
rect 27522 30064 27528 30116
rect 27580 30104 27586 30116
rect 27678 30107 27736 30113
rect 27678 30104 27690 30107
rect 27580 30076 27690 30104
rect 27580 30064 27586 30076
rect 27678 30073 27690 30076
rect 27724 30073 27736 30107
rect 27678 30067 27736 30073
rect 25590 30036 25596 30048
rect 24136 30008 25596 30036
rect 19153 29999 19211 30005
rect 25590 29996 25596 30008
rect 25648 29996 25654 30048
rect 28813 30039 28871 30045
rect 28813 30005 28825 30039
rect 28859 30036 28871 30039
rect 28902 30036 28908 30048
rect 28859 30008 28908 30036
rect 28859 30005 28871 30008
rect 28813 29999 28871 30005
rect 28902 29996 28908 30008
rect 28960 29996 28966 30048
rect 552 29946 31648 29968
rect 552 29894 4322 29946
rect 4374 29894 4386 29946
rect 4438 29894 4450 29946
rect 4502 29894 4514 29946
rect 4566 29894 4578 29946
rect 4630 29894 12096 29946
rect 12148 29894 12160 29946
rect 12212 29894 12224 29946
rect 12276 29894 12288 29946
rect 12340 29894 12352 29946
rect 12404 29894 19870 29946
rect 19922 29894 19934 29946
rect 19986 29894 19998 29946
rect 20050 29894 20062 29946
rect 20114 29894 20126 29946
rect 20178 29894 27644 29946
rect 27696 29894 27708 29946
rect 27760 29894 27772 29946
rect 27824 29894 27836 29946
rect 27888 29894 27900 29946
rect 27952 29894 31648 29946
rect 552 29872 31648 29894
rect 16758 29792 16764 29844
rect 16816 29792 16822 29844
rect 17586 29792 17592 29844
rect 17644 29792 17650 29844
rect 18601 29835 18659 29841
rect 18601 29801 18613 29835
rect 18647 29832 18659 29835
rect 18647 29804 19334 29832
rect 18647 29801 18659 29804
rect 18601 29795 18659 29801
rect 11882 29724 11888 29776
rect 11940 29764 11946 29776
rect 14642 29764 14648 29776
rect 11940 29736 14648 29764
rect 11940 29724 11946 29736
rect 14642 29724 14648 29736
rect 14700 29724 14706 29776
rect 16666 29724 16672 29776
rect 16724 29764 16730 29776
rect 17221 29767 17279 29773
rect 17221 29764 17233 29767
rect 16724 29736 17233 29764
rect 16724 29724 16730 29736
rect 17221 29733 17233 29736
rect 17267 29733 17279 29767
rect 17221 29727 17279 29733
rect 17402 29724 17408 29776
rect 17460 29773 17466 29776
rect 17460 29767 17479 29773
rect 17467 29733 17479 29767
rect 17460 29727 17479 29733
rect 17773 29767 17831 29773
rect 17773 29733 17785 29767
rect 17819 29764 17831 29767
rect 18138 29764 18144 29776
rect 17819 29736 18144 29764
rect 17819 29733 17831 29736
rect 17773 29727 17831 29733
rect 17460 29724 17466 29727
rect 18138 29724 18144 29736
rect 18196 29764 18202 29776
rect 19306 29764 19334 29804
rect 19610 29792 19616 29844
rect 19668 29832 19674 29844
rect 20349 29835 20407 29841
rect 20349 29832 20361 29835
rect 19668 29804 20361 29832
rect 19668 29792 19674 29804
rect 20272 29776 20300 29804
rect 20349 29801 20361 29804
rect 20395 29801 20407 29835
rect 20349 29795 20407 29801
rect 21726 29792 21732 29844
rect 21784 29832 21790 29844
rect 24302 29832 24308 29844
rect 21784 29804 24308 29832
rect 21784 29792 21790 29804
rect 24302 29792 24308 29804
rect 24360 29792 24366 29844
rect 26510 29792 26516 29844
rect 26568 29832 26574 29844
rect 26786 29832 26792 29844
rect 26568 29804 26792 29832
rect 26568 29792 26574 29804
rect 26786 29792 26792 29804
rect 26844 29792 26850 29844
rect 27614 29792 27620 29844
rect 27672 29792 27678 29844
rect 27801 29835 27859 29841
rect 27801 29801 27813 29835
rect 27847 29832 27859 29835
rect 28074 29832 28080 29844
rect 27847 29804 28080 29832
rect 27847 29801 27859 29804
rect 27801 29795 27859 29801
rect 28074 29792 28080 29804
rect 28132 29792 28138 29844
rect 19886 29764 19892 29776
rect 18196 29736 18644 29764
rect 19306 29736 19892 29764
rect 18196 29724 18202 29736
rect 14090 29656 14096 29708
rect 14148 29656 14154 29708
rect 14360 29699 14418 29705
rect 14360 29665 14372 29699
rect 14406 29696 14418 29699
rect 14734 29696 14740 29708
rect 14406 29668 14740 29696
rect 14406 29665 14418 29668
rect 14360 29659 14418 29665
rect 14734 29656 14740 29668
rect 14792 29656 14798 29708
rect 15930 29656 15936 29708
rect 15988 29696 15994 29708
rect 16393 29699 16451 29705
rect 16393 29696 16405 29699
rect 15988 29668 16405 29696
rect 15988 29656 15994 29668
rect 16393 29665 16405 29668
rect 16439 29696 16451 29699
rect 16482 29696 16488 29708
rect 16439 29668 16488 29696
rect 16439 29665 16451 29668
rect 16393 29659 16451 29665
rect 16482 29656 16488 29668
rect 16540 29656 16546 29708
rect 16853 29699 16911 29705
rect 16853 29665 16865 29699
rect 16899 29696 16911 29699
rect 17310 29696 17316 29708
rect 16899 29668 17316 29696
rect 16899 29665 16911 29668
rect 16853 29659 16911 29665
rect 17310 29656 17316 29668
rect 17368 29656 17374 29708
rect 17681 29699 17739 29705
rect 17681 29665 17693 29699
rect 17727 29665 17739 29699
rect 17681 29659 17739 29665
rect 16577 29631 16635 29637
rect 16577 29597 16589 29631
rect 16623 29628 16635 29631
rect 17034 29628 17040 29640
rect 16623 29600 17040 29628
rect 16623 29597 16635 29600
rect 16577 29591 16635 29597
rect 17034 29588 17040 29600
rect 17092 29588 17098 29640
rect 17218 29588 17224 29640
rect 17276 29628 17282 29640
rect 17696 29628 17724 29659
rect 17954 29656 17960 29708
rect 18012 29696 18018 29708
rect 18616 29705 18644 29736
rect 19886 29724 19892 29736
rect 19944 29764 19950 29776
rect 19944 29736 20208 29764
rect 19944 29724 19950 29736
rect 18233 29699 18291 29705
rect 18233 29696 18245 29699
rect 18012 29668 18245 29696
rect 18012 29656 18018 29668
rect 18233 29665 18245 29668
rect 18279 29665 18291 29699
rect 18233 29659 18291 29665
rect 18601 29699 18659 29705
rect 18601 29665 18613 29699
rect 18647 29665 18659 29699
rect 18601 29659 18659 29665
rect 18966 29656 18972 29708
rect 19024 29656 19030 29708
rect 19236 29699 19294 29705
rect 19236 29665 19248 29699
rect 19282 29696 19294 29699
rect 19610 29696 19616 29708
rect 19282 29668 19616 29696
rect 19282 29665 19294 29668
rect 19236 29659 19294 29665
rect 19610 29656 19616 29668
rect 19668 29656 19674 29708
rect 20180 29696 20208 29736
rect 20254 29724 20260 29776
rect 20312 29724 20318 29776
rect 23474 29764 23480 29776
rect 20732 29736 23480 29764
rect 20438 29696 20444 29708
rect 20180 29668 20444 29696
rect 20438 29656 20444 29668
rect 20496 29656 20502 29708
rect 20732 29705 20760 29736
rect 20717 29699 20775 29705
rect 20717 29665 20729 29699
rect 20763 29665 20775 29699
rect 20717 29659 20775 29665
rect 21726 29656 21732 29708
rect 21784 29656 21790 29708
rect 21818 29656 21824 29708
rect 21876 29656 21882 29708
rect 22002 29656 22008 29708
rect 22060 29656 22066 29708
rect 22278 29656 22284 29708
rect 22336 29656 22342 29708
rect 22370 29656 22376 29708
rect 22428 29656 22434 29708
rect 22756 29705 22784 29736
rect 23474 29724 23480 29736
rect 23532 29764 23538 29776
rect 26421 29767 26479 29773
rect 23532 29736 23888 29764
rect 23532 29724 23538 29736
rect 22741 29699 22799 29705
rect 22741 29665 22753 29699
rect 22787 29665 22799 29699
rect 22741 29659 22799 29665
rect 23566 29656 23572 29708
rect 23624 29656 23630 29708
rect 23860 29705 23888 29736
rect 26421 29733 26433 29767
rect 26467 29764 26479 29767
rect 26602 29764 26608 29776
rect 26467 29736 26608 29764
rect 26467 29733 26479 29736
rect 26421 29727 26479 29733
rect 26602 29724 26608 29736
rect 26660 29724 26666 29776
rect 23845 29699 23903 29705
rect 23845 29665 23857 29699
rect 23891 29665 23903 29699
rect 23845 29659 23903 29665
rect 25222 29656 25228 29708
rect 25280 29656 25286 29708
rect 25318 29699 25376 29705
rect 25318 29665 25330 29699
rect 25364 29665 25376 29699
rect 25318 29659 25376 29665
rect 18785 29631 18843 29637
rect 18785 29628 18797 29631
rect 17276 29600 18797 29628
rect 17276 29588 17282 29600
rect 18785 29597 18797 29600
rect 18831 29597 18843 29631
rect 18785 29591 18843 29597
rect 20806 29588 20812 29640
rect 20864 29628 20870 29640
rect 21836 29628 21864 29656
rect 20864 29600 21864 29628
rect 20864 29588 20870 29600
rect 15473 29563 15531 29569
rect 15473 29529 15485 29563
rect 15519 29560 15531 29563
rect 15519 29532 16620 29560
rect 15519 29529 15531 29532
rect 15473 29523 15531 29529
rect 16592 29504 16620 29532
rect 21174 29520 21180 29572
rect 21232 29560 21238 29572
rect 22388 29560 22416 29656
rect 25130 29588 25136 29640
rect 25188 29628 25194 29640
rect 25332 29628 25360 29659
rect 26694 29656 26700 29708
rect 26752 29656 26758 29708
rect 28442 29656 28448 29708
rect 28500 29656 28506 29708
rect 25188 29600 25360 29628
rect 25188 29588 25194 29600
rect 26602 29588 26608 29640
rect 26660 29588 26666 29640
rect 26786 29588 26792 29640
rect 26844 29588 26850 29640
rect 26881 29631 26939 29637
rect 26881 29597 26893 29631
rect 26927 29628 26939 29631
rect 27430 29628 27436 29640
rect 26927 29600 27436 29628
rect 26927 29597 26939 29600
rect 26881 29591 26939 29597
rect 27430 29588 27436 29600
rect 27488 29588 27494 29640
rect 28629 29631 28687 29637
rect 28629 29597 28641 29631
rect 28675 29628 28687 29631
rect 28902 29628 28908 29640
rect 28675 29600 28908 29628
rect 28675 29597 28687 29600
rect 28629 29591 28687 29597
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 21232 29532 22416 29560
rect 21232 29520 21238 29532
rect 23106 29520 23112 29572
rect 23164 29560 23170 29572
rect 23753 29563 23811 29569
rect 23753 29560 23765 29563
rect 23164 29532 23765 29560
rect 23164 29520 23170 29532
rect 23753 29529 23765 29532
rect 23799 29529 23811 29563
rect 23753 29523 23811 29529
rect 25593 29563 25651 29569
rect 25593 29529 25605 29563
rect 25639 29560 25651 29563
rect 25774 29560 25780 29572
rect 25639 29532 25780 29560
rect 25639 29529 25651 29532
rect 25593 29523 25651 29529
rect 25774 29520 25780 29532
rect 25832 29520 25838 29572
rect 28166 29520 28172 29572
rect 28224 29560 28230 29572
rect 28261 29563 28319 29569
rect 28261 29560 28273 29563
rect 28224 29532 28273 29560
rect 28224 29520 28230 29532
rect 28261 29529 28273 29532
rect 28307 29529 28319 29563
rect 28261 29523 28319 29529
rect 16114 29452 16120 29504
rect 16172 29452 16178 29504
rect 16482 29452 16488 29504
rect 16540 29452 16546 29504
rect 16574 29452 16580 29504
rect 16632 29452 16638 29504
rect 17405 29495 17463 29501
rect 17405 29461 17417 29495
rect 17451 29492 17463 29495
rect 18046 29492 18052 29504
rect 17451 29464 18052 29492
rect 17451 29461 17463 29464
rect 17405 29455 17463 29461
rect 18046 29452 18052 29464
rect 18104 29452 18110 29504
rect 18141 29495 18199 29501
rect 18141 29461 18153 29495
rect 18187 29492 18199 29495
rect 20346 29492 20352 29504
rect 18187 29464 20352 29492
rect 18187 29461 18199 29464
rect 18141 29455 18199 29461
rect 20346 29452 20352 29464
rect 20404 29452 20410 29504
rect 20438 29452 20444 29504
rect 20496 29492 20502 29504
rect 20625 29495 20683 29501
rect 20625 29492 20637 29495
rect 20496 29464 20637 29492
rect 20496 29452 20502 29464
rect 20625 29461 20637 29464
rect 20671 29461 20683 29495
rect 20625 29455 20683 29461
rect 22097 29495 22155 29501
rect 22097 29461 22109 29495
rect 22143 29492 22155 29495
rect 22186 29492 22192 29504
rect 22143 29464 22192 29492
rect 22143 29461 22155 29464
rect 22097 29455 22155 29461
rect 22186 29452 22192 29464
rect 22244 29452 22250 29504
rect 22646 29452 22652 29504
rect 22704 29452 22710 29504
rect 23198 29452 23204 29504
rect 23256 29492 23262 29504
rect 23385 29495 23443 29501
rect 23385 29492 23397 29495
rect 23256 29464 23397 29492
rect 23256 29452 23262 29464
rect 23385 29461 23397 29464
rect 23431 29461 23443 29495
rect 23385 29455 23443 29461
rect 27801 29495 27859 29501
rect 27801 29461 27813 29495
rect 27847 29492 27859 29495
rect 27982 29492 27988 29504
rect 27847 29464 27988 29492
rect 27847 29461 27859 29464
rect 27801 29455 27859 29461
rect 27982 29452 27988 29464
rect 28040 29452 28046 29504
rect 552 29402 31648 29424
rect 552 29350 3662 29402
rect 3714 29350 3726 29402
rect 3778 29350 3790 29402
rect 3842 29350 3854 29402
rect 3906 29350 3918 29402
rect 3970 29350 11436 29402
rect 11488 29350 11500 29402
rect 11552 29350 11564 29402
rect 11616 29350 11628 29402
rect 11680 29350 11692 29402
rect 11744 29350 19210 29402
rect 19262 29350 19274 29402
rect 19326 29350 19338 29402
rect 19390 29350 19402 29402
rect 19454 29350 19466 29402
rect 19518 29350 26984 29402
rect 27036 29350 27048 29402
rect 27100 29350 27112 29402
rect 27164 29350 27176 29402
rect 27228 29350 27240 29402
rect 27292 29350 31648 29402
rect 552 29328 31648 29350
rect 11514 29248 11520 29300
rect 11572 29288 11578 29300
rect 11882 29288 11888 29300
rect 11572 29260 11888 29288
rect 11572 29248 11578 29260
rect 11882 29248 11888 29260
rect 11940 29248 11946 29300
rect 13078 29248 13084 29300
rect 13136 29288 13142 29300
rect 14366 29288 14372 29300
rect 13136 29260 14372 29288
rect 13136 29248 13142 29260
rect 14366 29248 14372 29260
rect 14424 29248 14430 29300
rect 14734 29248 14740 29300
rect 14792 29248 14798 29300
rect 16666 29248 16672 29300
rect 16724 29288 16730 29300
rect 17497 29291 17555 29297
rect 17497 29288 17509 29291
rect 16724 29260 17509 29288
rect 16724 29248 16730 29260
rect 17497 29257 17509 29260
rect 17543 29288 17555 29291
rect 17954 29288 17960 29300
rect 17543 29260 17960 29288
rect 17543 29257 17555 29260
rect 17497 29251 17555 29257
rect 17954 29248 17960 29260
rect 18012 29248 18018 29300
rect 18138 29248 18144 29300
rect 18196 29248 18202 29300
rect 19610 29248 19616 29300
rect 19668 29248 19674 29300
rect 25590 29248 25596 29300
rect 25648 29288 25654 29300
rect 26053 29291 26111 29297
rect 26053 29288 26065 29291
rect 25648 29260 26065 29288
rect 25648 29248 25654 29260
rect 26053 29257 26065 29260
rect 26099 29257 26111 29291
rect 26053 29251 26111 29257
rect 11330 29180 11336 29232
rect 11388 29220 11394 29232
rect 11425 29223 11483 29229
rect 11425 29220 11437 29223
rect 11388 29192 11437 29220
rect 11388 29180 11394 29192
rect 11425 29189 11437 29192
rect 11471 29189 11483 29223
rect 11425 29183 11483 29189
rect 11698 29180 11704 29232
rect 11756 29220 11762 29232
rect 15286 29220 15292 29232
rect 11756 29192 14044 29220
rect 11756 29180 11762 29192
rect 14016 29152 14044 29192
rect 15120 29192 15292 29220
rect 14645 29155 14703 29161
rect 14645 29152 14657 29155
rect 11256 29124 12388 29152
rect 9398 29044 9404 29096
rect 9456 29084 9462 29096
rect 11256 29093 11284 29124
rect 11241 29087 11299 29093
rect 11241 29084 11253 29087
rect 9456 29056 11253 29084
rect 9456 29044 9462 29056
rect 11241 29053 11253 29056
rect 11287 29053 11299 29087
rect 11241 29047 11299 29053
rect 11425 29087 11483 29093
rect 11425 29053 11437 29087
rect 11471 29084 11483 29087
rect 11514 29084 11520 29096
rect 11471 29056 11520 29084
rect 11471 29053 11483 29056
rect 11425 29047 11483 29053
rect 11514 29044 11520 29056
rect 11572 29044 11578 29096
rect 11698 29044 11704 29096
rect 11756 29044 11762 29096
rect 12360 29093 12388 29124
rect 14016 29124 14657 29152
rect 12345 29087 12403 29093
rect 12345 29053 12357 29087
rect 12391 29084 12403 29087
rect 12434 29084 12440 29096
rect 12391 29056 12440 29084
rect 12391 29053 12403 29056
rect 12345 29047 12403 29053
rect 12434 29044 12440 29056
rect 12492 29044 12498 29096
rect 12805 29087 12863 29093
rect 12805 29053 12817 29087
rect 12851 29084 12863 29087
rect 12851 29056 12940 29084
rect 12851 29053 12863 29056
rect 12805 29047 12863 29053
rect 11609 29019 11667 29025
rect 11609 28985 11621 29019
rect 11655 29016 11667 29019
rect 11974 29016 11980 29028
rect 11655 28988 11980 29016
rect 11655 28985 11667 28988
rect 11609 28979 11667 28985
rect 11974 28976 11980 28988
rect 12032 28976 12038 29028
rect 11054 28908 11060 28960
rect 11112 28948 11118 28960
rect 11149 28951 11207 28957
rect 11149 28948 11161 28951
rect 11112 28920 11161 28948
rect 11112 28908 11118 28920
rect 11149 28917 11161 28920
rect 11195 28917 11207 28951
rect 11149 28911 11207 28917
rect 12434 28908 12440 28960
rect 12492 28908 12498 28960
rect 12618 28908 12624 28960
rect 12676 28908 12682 28960
rect 12912 28948 12940 29056
rect 13078 29044 13084 29096
rect 13136 29044 13142 29096
rect 13170 29044 13176 29096
rect 13228 29044 13234 29096
rect 13357 29087 13415 29093
rect 13357 29053 13369 29087
rect 13403 29084 13415 29087
rect 14016 29084 14044 29124
rect 14645 29121 14657 29124
rect 14691 29121 14703 29155
rect 14645 29115 14703 29121
rect 13403 29056 14044 29084
rect 13403 29053 13415 29056
rect 13357 29047 13415 29053
rect 14182 29044 14188 29096
rect 14240 29044 14246 29096
rect 14277 29087 14335 29093
rect 14277 29053 14289 29087
rect 14323 29084 14335 29087
rect 14366 29084 14372 29096
rect 14323 29056 14372 29084
rect 14323 29053 14335 29056
rect 14277 29047 14335 29053
rect 14366 29044 14372 29056
rect 14424 29044 14430 29096
rect 15120 29093 15148 29192
rect 15286 29180 15292 29192
rect 15344 29180 15350 29232
rect 16206 29180 16212 29232
rect 16264 29220 16270 29232
rect 17313 29223 17371 29229
rect 17313 29220 17325 29223
rect 16264 29192 17325 29220
rect 16264 29180 16270 29192
rect 17313 29189 17325 29192
rect 17359 29189 17371 29223
rect 19886 29220 19892 29232
rect 17313 29183 17371 29189
rect 19536 29192 19892 29220
rect 16114 29152 16120 29164
rect 15212 29124 16120 29152
rect 15212 29093 15240 29124
rect 16114 29112 16120 29124
rect 16172 29112 16178 29164
rect 18506 29152 18512 29164
rect 18340 29124 18512 29152
rect 15013 29087 15071 29093
rect 15013 29053 15025 29087
rect 15059 29053 15071 29087
rect 15013 29047 15071 29053
rect 15105 29087 15163 29093
rect 15105 29053 15117 29087
rect 15151 29053 15163 29087
rect 15105 29047 15163 29053
rect 15197 29087 15255 29093
rect 15197 29053 15209 29087
rect 15243 29053 15255 29087
rect 15197 29047 15255 29053
rect 15381 29087 15439 29093
rect 15381 29053 15393 29087
rect 15427 29084 15439 29087
rect 15654 29084 15660 29096
rect 15427 29056 15660 29084
rect 15427 29053 15439 29056
rect 15381 29047 15439 29053
rect 12989 29019 13047 29025
rect 12989 28985 13001 29019
rect 13035 29016 13047 29019
rect 13541 29019 13599 29025
rect 13541 29016 13553 29019
rect 13035 28988 13553 29016
rect 13035 28985 13047 28988
rect 12989 28979 13047 28985
rect 13541 28985 13553 28988
rect 13587 28985 13599 29019
rect 14200 29016 14228 29044
rect 14461 29019 14519 29025
rect 14461 29016 14473 29019
rect 14200 28988 14473 29016
rect 13541 28979 13599 28985
rect 14461 28985 14473 28988
rect 14507 28985 14519 29019
rect 15028 29016 15056 29047
rect 15654 29044 15660 29056
rect 15712 29044 15718 29096
rect 18340 29093 18368 29124
rect 18506 29112 18512 29124
rect 18564 29112 18570 29164
rect 18325 29087 18383 29093
rect 18325 29053 18337 29087
rect 18371 29053 18383 29087
rect 18325 29047 18383 29053
rect 19337 29087 19395 29093
rect 19337 29053 19349 29087
rect 19383 29084 19395 29087
rect 19426 29084 19432 29096
rect 19383 29056 19432 29084
rect 19383 29053 19395 29056
rect 19337 29047 19395 29053
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 19536 29093 19564 29192
rect 19886 29180 19892 29192
rect 19944 29180 19950 29232
rect 25869 29223 25927 29229
rect 25869 29189 25881 29223
rect 25915 29220 25927 29223
rect 26878 29220 26884 29232
rect 25915 29192 26884 29220
rect 25915 29189 25927 29192
rect 25869 29183 25927 29189
rect 26878 29180 26884 29192
rect 26936 29180 26942 29232
rect 20346 29152 20352 29164
rect 20088 29124 20352 29152
rect 19521 29087 19579 29093
rect 19521 29053 19533 29087
rect 19567 29053 19579 29087
rect 19521 29047 19579 29053
rect 19889 29087 19947 29093
rect 19889 29053 19901 29087
rect 19935 29084 19947 29087
rect 20088 29084 20116 29124
rect 20346 29112 20352 29124
rect 20404 29112 20410 29164
rect 20438 29112 20444 29164
rect 20496 29112 20502 29164
rect 23658 29112 23664 29164
rect 23716 29152 23722 29164
rect 24213 29155 24271 29161
rect 24213 29152 24225 29155
rect 23716 29124 24225 29152
rect 23716 29112 23722 29124
rect 24213 29121 24225 29124
rect 24259 29121 24271 29155
rect 24213 29115 24271 29121
rect 25774 29112 25780 29164
rect 25832 29112 25838 29164
rect 27801 29155 27859 29161
rect 27801 29121 27813 29155
rect 27847 29152 27859 29155
rect 28350 29152 28356 29164
rect 27847 29124 28356 29152
rect 27847 29121 27859 29124
rect 27801 29115 27859 29121
rect 28350 29112 28356 29124
rect 28408 29112 28414 29164
rect 19935 29056 20116 29084
rect 20165 29087 20223 29093
rect 19935 29053 19947 29056
rect 19889 29047 19947 29053
rect 20165 29053 20177 29087
rect 20211 29053 20223 29087
rect 20165 29047 20223 29053
rect 21913 29087 21971 29093
rect 21913 29053 21925 29087
rect 21959 29084 21971 29087
rect 22646 29084 22652 29096
rect 21959 29056 22652 29084
rect 21959 29053 21971 29056
rect 21913 29047 21971 29053
rect 16666 29016 16672 29028
rect 15028 28988 16672 29016
rect 14461 28979 14519 28985
rect 16666 28976 16672 28988
rect 16724 29016 16730 29028
rect 17037 29019 17095 29025
rect 17037 29016 17049 29019
rect 16724 28988 17049 29016
rect 16724 28976 16730 28988
rect 17037 28985 17049 28988
rect 17083 28985 17095 29019
rect 17037 28979 17095 28985
rect 18414 28976 18420 29028
rect 18472 29016 18478 29028
rect 18509 29019 18567 29025
rect 18509 29016 18521 29019
rect 18472 28988 18521 29016
rect 18472 28976 18478 28988
rect 18509 28985 18521 28988
rect 18555 28985 18567 29019
rect 18509 28979 18567 28985
rect 19794 28976 19800 29028
rect 19852 29016 19858 29028
rect 20073 29019 20131 29025
rect 20073 29016 20085 29019
rect 19852 28988 20085 29016
rect 19852 28976 19858 28988
rect 20073 28985 20085 28988
rect 20119 28985 20131 29019
rect 20180 29016 20208 29047
rect 22646 29044 22652 29056
rect 22704 29044 22710 29096
rect 23382 29044 23388 29096
rect 23440 29084 23446 29096
rect 23845 29087 23903 29093
rect 23845 29084 23857 29087
rect 23440 29056 23857 29084
rect 23440 29044 23446 29056
rect 23845 29053 23857 29056
rect 23891 29053 23903 29087
rect 23845 29047 23903 29053
rect 24026 29044 24032 29096
rect 24084 29044 24090 29096
rect 25130 29044 25136 29096
rect 25188 29044 25194 29096
rect 25222 29044 25228 29096
rect 25280 29084 25286 29096
rect 25501 29087 25559 29093
rect 25280 29056 25452 29084
rect 25280 29044 25286 29056
rect 20438 29016 20444 29028
rect 20180 28988 20444 29016
rect 20073 28979 20131 28985
rect 20438 28976 20444 28988
rect 20496 28976 20502 29028
rect 20530 28976 20536 29028
rect 20588 29016 20594 29028
rect 22186 29025 22192 29028
rect 20686 29019 20744 29025
rect 20686 29016 20698 29019
rect 20588 28988 20698 29016
rect 20588 28976 20594 28988
rect 20686 28985 20698 28988
rect 20732 28985 20744 29019
rect 22180 29016 22192 29025
rect 20686 28979 20744 28985
rect 21652 28988 21956 29016
rect 22147 28988 22192 29016
rect 13173 28951 13231 28957
rect 13173 28948 13185 28951
rect 12912 28920 13185 28948
rect 13173 28917 13185 28920
rect 13219 28917 13231 28951
rect 13173 28911 13231 28917
rect 19334 28908 19340 28960
rect 19392 28948 19398 28960
rect 21652 28948 21680 28988
rect 21928 28960 21956 28988
rect 22180 28979 22192 28988
rect 22186 28976 22192 28979
rect 22244 28976 22250 29028
rect 23198 28976 23204 29028
rect 23256 29016 23262 29028
rect 23477 29019 23535 29025
rect 23477 29016 23489 29019
rect 23256 28988 23489 29016
rect 23256 28976 23262 28988
rect 23477 28985 23489 28988
rect 23523 28985 23535 29019
rect 25424 29016 25452 29056
rect 25501 29053 25513 29087
rect 25547 29084 25559 29087
rect 25685 29087 25743 29093
rect 25685 29084 25697 29087
rect 25547 29056 25697 29084
rect 25547 29053 25559 29056
rect 25501 29047 25559 29053
rect 25685 29053 25697 29056
rect 25731 29053 25743 29087
rect 25685 29047 25743 29053
rect 25866 29044 25872 29096
rect 25924 29044 25930 29096
rect 25958 29044 25964 29096
rect 26016 29084 26022 29096
rect 26145 29087 26203 29093
rect 26145 29084 26157 29087
rect 26016 29056 26157 29084
rect 26016 29044 26022 29056
rect 26145 29053 26157 29056
rect 26191 29053 26203 29087
rect 26145 29047 26203 29053
rect 27338 29044 27344 29096
rect 27396 29084 27402 29096
rect 28445 29087 28503 29093
rect 28445 29084 28457 29087
rect 27396 29056 28457 29084
rect 27396 29044 27402 29056
rect 28445 29053 28457 29056
rect 28491 29053 28503 29087
rect 28445 29047 28503 29053
rect 27985 29019 28043 29025
rect 27985 29016 27997 29019
rect 25424 28988 27997 29016
rect 23477 28979 23535 28985
rect 27985 28985 27997 28988
rect 28031 29016 28043 29019
rect 28031 28988 28120 29016
rect 28031 28985 28043 28988
rect 27985 28979 28043 28985
rect 28092 28960 28120 28988
rect 28166 28976 28172 29028
rect 28224 28976 28230 29028
rect 28353 29019 28411 29025
rect 28353 28985 28365 29019
rect 28399 29016 28411 29019
rect 29086 29016 29092 29028
rect 28399 28988 29092 29016
rect 28399 28985 28411 28988
rect 28353 28979 28411 28985
rect 29086 28976 29092 28988
rect 29144 28976 29150 29028
rect 19392 28920 21680 28948
rect 19392 28908 19398 28920
rect 21726 28908 21732 28960
rect 21784 28948 21790 28960
rect 21821 28951 21879 28957
rect 21821 28948 21833 28951
rect 21784 28920 21833 28948
rect 21784 28908 21790 28920
rect 21821 28917 21833 28920
rect 21867 28917 21879 28951
rect 21821 28911 21879 28917
rect 21910 28908 21916 28960
rect 21968 28908 21974 28960
rect 22462 28908 22468 28960
rect 22520 28948 22526 28960
rect 23290 28948 23296 28960
rect 22520 28920 23296 28948
rect 22520 28908 22526 28920
rect 23290 28908 23296 28920
rect 23348 28908 23354 28960
rect 28074 28908 28080 28960
rect 28132 28908 28138 28960
rect 552 28858 31648 28880
rect 552 28806 4322 28858
rect 4374 28806 4386 28858
rect 4438 28806 4450 28858
rect 4502 28806 4514 28858
rect 4566 28806 4578 28858
rect 4630 28806 12096 28858
rect 12148 28806 12160 28858
rect 12212 28806 12224 28858
rect 12276 28806 12288 28858
rect 12340 28806 12352 28858
rect 12404 28806 19870 28858
rect 19922 28806 19934 28858
rect 19986 28806 19998 28858
rect 20050 28806 20062 28858
rect 20114 28806 20126 28858
rect 20178 28806 27644 28858
rect 27696 28806 27708 28858
rect 27760 28806 27772 28858
rect 27824 28806 27836 28858
rect 27888 28806 27900 28858
rect 27952 28806 31648 28858
rect 552 28784 31648 28806
rect 11974 28704 11980 28756
rect 12032 28744 12038 28756
rect 12345 28747 12403 28753
rect 12345 28744 12357 28747
rect 12032 28716 12357 28744
rect 12032 28704 12038 28716
rect 12345 28713 12357 28716
rect 12391 28713 12403 28747
rect 12345 28707 12403 28713
rect 14274 28704 14280 28756
rect 14332 28704 14338 28756
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 14921 28747 14979 28753
rect 14921 28744 14933 28747
rect 14884 28716 14933 28744
rect 14884 28704 14890 28716
rect 14921 28713 14933 28716
rect 14967 28713 14979 28747
rect 15565 28747 15623 28753
rect 15565 28744 15577 28747
rect 14921 28707 14979 28713
rect 15120 28716 15577 28744
rect 14182 28636 14188 28688
rect 14240 28636 14246 28688
rect 10965 28611 11023 28617
rect 10965 28577 10977 28611
rect 11011 28608 11023 28611
rect 11054 28608 11060 28620
rect 11011 28580 11060 28608
rect 11011 28577 11023 28580
rect 10965 28571 11023 28577
rect 11054 28568 11060 28580
rect 11112 28568 11118 28620
rect 11238 28617 11244 28620
rect 11232 28608 11244 28617
rect 11199 28580 11244 28608
rect 11232 28571 11244 28580
rect 11238 28568 11244 28571
rect 11296 28568 11302 28620
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 12529 28611 12587 28617
rect 12529 28608 12541 28611
rect 12492 28580 12541 28608
rect 12492 28568 12498 28580
rect 12529 28577 12541 28580
rect 12575 28577 12587 28611
rect 12529 28571 12587 28577
rect 12618 28568 12624 28620
rect 12676 28608 12682 28620
rect 12805 28611 12863 28617
rect 12805 28608 12817 28611
rect 12676 28580 12817 28608
rect 12676 28568 12682 28580
rect 12805 28577 12817 28580
rect 12851 28577 12863 28611
rect 12805 28571 12863 28577
rect 14645 28611 14703 28617
rect 14645 28577 14657 28611
rect 14691 28608 14703 28611
rect 14844 28608 14872 28704
rect 15120 28688 15148 28716
rect 15565 28713 15577 28716
rect 15611 28713 15623 28747
rect 15565 28707 15623 28713
rect 15733 28747 15791 28753
rect 15733 28713 15745 28747
rect 15779 28744 15791 28747
rect 16298 28744 16304 28756
rect 15779 28716 16304 28744
rect 15779 28713 15791 28716
rect 15733 28707 15791 28713
rect 16298 28704 16304 28716
rect 16356 28744 16362 28756
rect 16853 28747 16911 28753
rect 16853 28744 16865 28747
rect 16356 28716 16865 28744
rect 16356 28704 16362 28716
rect 16853 28713 16865 28716
rect 16899 28713 16911 28747
rect 16853 28707 16911 28713
rect 17402 28704 17408 28756
rect 17460 28704 17466 28756
rect 20530 28704 20536 28756
rect 20588 28704 20594 28756
rect 20898 28704 20904 28756
rect 20956 28744 20962 28756
rect 20956 28716 21864 28744
rect 20956 28704 20962 28716
rect 15102 28636 15108 28688
rect 15160 28636 15166 28688
rect 15933 28679 15991 28685
rect 15933 28645 15945 28679
rect 15979 28645 15991 28679
rect 18506 28676 18512 28688
rect 15933 28639 15991 28645
rect 16776 28648 18512 28676
rect 14691 28580 14872 28608
rect 15289 28611 15347 28617
rect 14691 28577 14703 28580
rect 14645 28571 14703 28577
rect 15289 28577 15301 28611
rect 15335 28577 15347 28611
rect 15948 28608 15976 28639
rect 16298 28608 16304 28620
rect 15948 28580 16304 28608
rect 15289 28571 15347 28577
rect 13170 28500 13176 28552
rect 13228 28540 13234 28552
rect 13228 28512 13492 28540
rect 13228 28500 13234 28512
rect 13464 28472 13492 28512
rect 14458 28500 14464 28552
rect 14516 28500 14522 28552
rect 14550 28500 14556 28552
rect 14608 28500 14614 28552
rect 14734 28500 14740 28552
rect 14792 28500 14798 28552
rect 15304 28540 15332 28571
rect 16298 28568 16304 28580
rect 16356 28568 16362 28620
rect 16776 28617 16804 28648
rect 16761 28611 16819 28617
rect 16761 28577 16773 28611
rect 16807 28608 16819 28611
rect 16850 28608 16856 28620
rect 16807 28580 16856 28608
rect 16807 28577 16819 28580
rect 16761 28571 16819 28577
rect 16850 28568 16856 28580
rect 16908 28568 16914 28620
rect 17512 28617 17540 28648
rect 18506 28636 18512 28648
rect 18564 28636 18570 28688
rect 21634 28636 21640 28688
rect 21692 28636 21698 28688
rect 21836 28676 21864 28716
rect 21910 28704 21916 28756
rect 21968 28744 21974 28756
rect 21968 28716 22232 28744
rect 21968 28704 21974 28716
rect 22204 28676 22232 28716
rect 22278 28704 22284 28756
rect 22336 28744 22342 28756
rect 22741 28747 22799 28753
rect 22741 28744 22753 28747
rect 22336 28716 22753 28744
rect 22336 28704 22342 28716
rect 22741 28713 22753 28716
rect 22787 28713 22799 28747
rect 22741 28707 22799 28713
rect 26786 28704 26792 28756
rect 26844 28744 26850 28756
rect 27157 28747 27215 28753
rect 27157 28744 27169 28747
rect 26844 28716 27169 28744
rect 26844 28704 26850 28716
rect 27157 28713 27169 28716
rect 27203 28713 27215 28747
rect 27157 28707 27215 28713
rect 23198 28676 23204 28688
rect 21836 28648 22140 28676
rect 22204 28648 23204 28676
rect 16945 28611 17003 28617
rect 16945 28577 16957 28611
rect 16991 28608 17003 28611
rect 17313 28611 17371 28617
rect 17313 28608 17325 28611
rect 16991 28580 17325 28608
rect 16991 28577 17003 28580
rect 16945 28571 17003 28577
rect 17313 28577 17325 28580
rect 17359 28577 17371 28611
rect 17313 28571 17371 28577
rect 17497 28611 17555 28617
rect 17497 28577 17509 28611
rect 17543 28577 17555 28611
rect 17497 28571 17555 28577
rect 15930 28540 15936 28552
rect 15304 28512 15936 28540
rect 15930 28500 15936 28512
rect 15988 28500 15994 28552
rect 17328 28540 17356 28571
rect 17862 28568 17868 28620
rect 17920 28568 17926 28620
rect 18049 28611 18107 28617
rect 18049 28577 18061 28611
rect 18095 28608 18107 28611
rect 19334 28608 19340 28620
rect 18095 28580 19340 28608
rect 18095 28577 18107 28580
rect 18049 28571 18107 28577
rect 18414 28540 18420 28552
rect 17328 28512 18420 28540
rect 18414 28500 18420 28512
rect 18472 28500 18478 28552
rect 16206 28472 16212 28484
rect 13464 28444 16212 28472
rect 16206 28432 16212 28444
rect 16264 28472 16270 28484
rect 18524 28472 18552 28580
rect 19334 28568 19340 28580
rect 19392 28568 19398 28620
rect 20165 28611 20223 28617
rect 20165 28577 20177 28611
rect 20211 28608 20223 28611
rect 20254 28608 20260 28620
rect 20211 28580 20260 28608
rect 20211 28577 20223 28580
rect 20165 28571 20223 28577
rect 20254 28568 20260 28580
rect 20312 28568 20318 28620
rect 20717 28611 20775 28617
rect 20717 28577 20729 28611
rect 20763 28608 20775 28611
rect 21269 28611 21327 28617
rect 21269 28608 21281 28611
rect 20763 28580 21281 28608
rect 20763 28577 20775 28580
rect 20717 28571 20775 28577
rect 21269 28577 21281 28580
rect 21315 28577 21327 28611
rect 21269 28571 21327 28577
rect 21450 28568 21456 28620
rect 21508 28568 21514 28620
rect 21545 28611 21603 28617
rect 21545 28577 21557 28611
rect 21591 28577 21603 28611
rect 21545 28571 21603 28577
rect 21755 28611 21813 28617
rect 21755 28577 21767 28611
rect 21801 28577 21813 28611
rect 21755 28571 21813 28577
rect 20349 28543 20407 28549
rect 20349 28509 20361 28543
rect 20395 28540 20407 28543
rect 20530 28540 20536 28552
rect 20395 28512 20536 28540
rect 20395 28509 20407 28512
rect 20349 28503 20407 28509
rect 20530 28500 20536 28512
rect 20588 28500 20594 28552
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28540 20959 28543
rect 21174 28540 21180 28552
rect 20947 28512 21180 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 21174 28500 21180 28512
rect 21232 28500 21238 28552
rect 16264 28444 18552 28472
rect 16264 28432 16270 28444
rect 15749 28407 15807 28413
rect 15749 28373 15761 28407
rect 15795 28404 15807 28407
rect 16666 28404 16672 28416
rect 15795 28376 16672 28404
rect 15795 28373 15807 28376
rect 15749 28367 15807 28373
rect 16666 28364 16672 28376
rect 16724 28364 16730 28416
rect 17954 28364 17960 28416
rect 18012 28364 18018 28416
rect 19978 28364 19984 28416
rect 20036 28364 20042 28416
rect 21560 28404 21588 28571
rect 21770 28540 21798 28571
rect 21910 28568 21916 28620
rect 21968 28568 21974 28620
rect 22112 28617 22140 28648
rect 23198 28636 23204 28648
rect 23256 28636 23262 28688
rect 23382 28685 23388 28688
rect 23376 28676 23388 28685
rect 23343 28648 23388 28676
rect 23376 28639 23388 28648
rect 23382 28636 23388 28639
rect 23440 28636 23446 28688
rect 25590 28636 25596 28688
rect 25648 28636 25654 28688
rect 22097 28611 22155 28617
rect 22097 28577 22109 28611
rect 22143 28577 22155 28611
rect 22097 28571 22155 28577
rect 22235 28611 22293 28617
rect 22235 28577 22247 28611
rect 22281 28577 22293 28611
rect 22235 28571 22293 28577
rect 22373 28611 22431 28617
rect 22373 28577 22385 28611
rect 22419 28577 22431 28611
rect 22373 28571 22431 28577
rect 22002 28540 22008 28552
rect 21770 28512 22008 28540
rect 22002 28500 22008 28512
rect 22060 28540 22066 28552
rect 22250 28540 22278 28571
rect 22060 28512 22278 28540
rect 22060 28500 22066 28512
rect 21634 28432 21640 28484
rect 21692 28472 21698 28484
rect 22388 28472 22416 28571
rect 22462 28568 22468 28620
rect 22520 28568 22526 28620
rect 22554 28568 22560 28620
rect 22612 28568 22618 28620
rect 23106 28568 23112 28620
rect 23164 28568 23170 28620
rect 24578 28608 24584 28620
rect 24136 28580 24584 28608
rect 21692 28444 22416 28472
rect 21692 28432 21698 28444
rect 21726 28404 21732 28416
rect 21560 28376 21732 28404
rect 21726 28364 21732 28376
rect 21784 28404 21790 28416
rect 24136 28404 24164 28580
rect 24578 28568 24584 28580
rect 24636 28608 24642 28620
rect 25317 28611 25375 28617
rect 25317 28608 25329 28611
rect 24636 28580 25329 28608
rect 24636 28568 24642 28580
rect 25317 28577 25329 28580
rect 25363 28577 25375 28611
rect 25317 28571 25375 28577
rect 25409 28611 25467 28617
rect 25409 28577 25421 28611
rect 25455 28608 25467 28611
rect 25961 28611 26019 28617
rect 25961 28608 25973 28611
rect 25455 28580 25973 28608
rect 25455 28577 25467 28580
rect 25409 28571 25467 28577
rect 25961 28577 25973 28580
rect 26007 28608 26019 28611
rect 26421 28611 26479 28617
rect 26421 28608 26433 28611
rect 26007 28580 26433 28608
rect 26007 28577 26019 28580
rect 25961 28571 26019 28577
rect 26421 28577 26433 28580
rect 26467 28577 26479 28611
rect 26421 28571 26479 28577
rect 26605 28611 26663 28617
rect 26605 28577 26617 28611
rect 26651 28577 26663 28611
rect 26605 28571 26663 28577
rect 25685 28543 25743 28549
rect 25685 28509 25697 28543
rect 25731 28509 25743 28543
rect 25685 28503 25743 28509
rect 26053 28543 26111 28549
rect 26053 28509 26065 28543
rect 26099 28540 26111 28543
rect 26620 28540 26648 28571
rect 26878 28568 26884 28620
rect 26936 28568 26942 28620
rect 28258 28568 28264 28620
rect 28316 28608 28322 28620
rect 28822 28611 28880 28617
rect 28822 28608 28834 28611
rect 28316 28580 28834 28608
rect 28316 28568 28322 28580
rect 28822 28577 28834 28580
rect 28868 28577 28880 28611
rect 28822 28571 28880 28577
rect 29086 28568 29092 28620
rect 29144 28568 29150 28620
rect 27338 28540 27344 28552
rect 26099 28512 27344 28540
rect 26099 28509 26111 28512
rect 26053 28503 26111 28509
rect 25700 28472 25728 28503
rect 27338 28500 27344 28512
rect 27396 28500 27402 28552
rect 25958 28472 25964 28484
rect 25700 28444 25964 28472
rect 25958 28432 25964 28444
rect 26016 28432 26022 28484
rect 21784 28376 24164 28404
rect 24489 28407 24547 28413
rect 21784 28364 21790 28376
rect 24489 28373 24501 28407
rect 24535 28404 24547 28407
rect 24946 28404 24952 28416
rect 24535 28376 24952 28404
rect 24535 28373 24547 28376
rect 24489 28367 24547 28373
rect 24946 28364 24952 28376
rect 25004 28364 25010 28416
rect 26237 28407 26295 28413
rect 26237 28373 26249 28407
rect 26283 28404 26295 28407
rect 26697 28407 26755 28413
rect 26697 28404 26709 28407
rect 26283 28376 26709 28404
rect 26283 28373 26295 28376
rect 26237 28367 26295 28373
rect 26697 28373 26709 28376
rect 26743 28373 26755 28407
rect 26697 28367 26755 28373
rect 26786 28364 26792 28416
rect 26844 28364 26850 28416
rect 27709 28407 27767 28413
rect 27709 28373 27721 28407
rect 27755 28404 27767 28407
rect 28074 28404 28080 28416
rect 27755 28376 28080 28404
rect 27755 28373 27767 28376
rect 27709 28367 27767 28373
rect 28074 28364 28080 28376
rect 28132 28404 28138 28416
rect 28442 28404 28448 28416
rect 28132 28376 28448 28404
rect 28132 28364 28138 28376
rect 28442 28364 28448 28376
rect 28500 28364 28506 28416
rect 552 28314 31648 28336
rect 552 28262 3662 28314
rect 3714 28262 3726 28314
rect 3778 28262 3790 28314
rect 3842 28262 3854 28314
rect 3906 28262 3918 28314
rect 3970 28262 11436 28314
rect 11488 28262 11500 28314
rect 11552 28262 11564 28314
rect 11616 28262 11628 28314
rect 11680 28262 11692 28314
rect 11744 28262 19210 28314
rect 19262 28262 19274 28314
rect 19326 28262 19338 28314
rect 19390 28262 19402 28314
rect 19454 28262 19466 28314
rect 19518 28262 26984 28314
rect 27036 28262 27048 28314
rect 27100 28262 27112 28314
rect 27164 28262 27176 28314
rect 27228 28262 27240 28314
rect 27292 28262 31648 28314
rect 552 28240 31648 28262
rect 11238 28160 11244 28212
rect 11296 28200 11302 28212
rect 11425 28203 11483 28209
rect 11425 28200 11437 28203
rect 11296 28172 11437 28200
rect 11296 28160 11302 28172
rect 11425 28169 11437 28172
rect 11471 28169 11483 28203
rect 11425 28163 11483 28169
rect 13725 28203 13783 28209
rect 13725 28169 13737 28203
rect 13771 28200 13783 28203
rect 14550 28200 14556 28212
rect 13771 28172 14556 28200
rect 13771 28169 13783 28172
rect 13725 28163 13783 28169
rect 14550 28160 14556 28172
rect 14608 28160 14614 28212
rect 15841 28203 15899 28209
rect 15841 28169 15853 28203
rect 15887 28200 15899 28203
rect 16390 28200 16396 28212
rect 15887 28172 16396 28200
rect 15887 28169 15899 28172
rect 15841 28163 15899 28169
rect 16390 28160 16396 28172
rect 16448 28160 16454 28212
rect 17494 28200 17500 28212
rect 16500 28172 17500 28200
rect 15930 28092 15936 28144
rect 15988 28092 15994 28144
rect 16114 28092 16120 28144
rect 16172 28132 16178 28144
rect 16500 28132 16528 28172
rect 17494 28160 17500 28172
rect 17552 28160 17558 28212
rect 18138 28200 18144 28212
rect 17604 28172 18144 28200
rect 16172 28104 16528 28132
rect 17313 28135 17371 28141
rect 16172 28092 16178 28104
rect 17313 28101 17325 28135
rect 17359 28132 17371 28135
rect 17604 28132 17632 28172
rect 18138 28160 18144 28172
rect 18196 28160 18202 28212
rect 19613 28203 19671 28209
rect 19613 28169 19625 28203
rect 19659 28200 19671 28203
rect 22094 28200 22100 28212
rect 19659 28172 22100 28200
rect 19659 28169 19671 28172
rect 19613 28163 19671 28169
rect 22094 28160 22100 28172
rect 22152 28160 22158 28212
rect 23845 28203 23903 28209
rect 23845 28169 23857 28203
rect 23891 28200 23903 28203
rect 24026 28200 24032 28212
rect 23891 28172 24032 28200
rect 23891 28169 23903 28172
rect 23845 28163 23903 28169
rect 24026 28160 24032 28172
rect 24084 28160 24090 28212
rect 24765 28203 24823 28209
rect 24765 28169 24777 28203
rect 24811 28200 24823 28203
rect 24946 28200 24952 28212
rect 24811 28172 24952 28200
rect 24811 28169 24823 28172
rect 24765 28163 24823 28169
rect 17359 28104 17632 28132
rect 17681 28135 17739 28141
rect 17359 28101 17371 28104
rect 17313 28095 17371 28101
rect 17681 28101 17693 28135
rect 17727 28132 17739 28135
rect 18414 28132 18420 28144
rect 17727 28104 18420 28132
rect 17727 28101 17739 28104
rect 17681 28095 17739 28101
rect 16758 28064 16764 28076
rect 15672 28036 16764 28064
rect 11330 27956 11336 28008
rect 11388 27956 11394 28008
rect 11517 27999 11575 28005
rect 11517 27965 11529 27999
rect 11563 27996 11575 27999
rect 11698 27996 11704 28008
rect 11563 27968 11704 27996
rect 11563 27965 11575 27968
rect 11517 27959 11575 27965
rect 11698 27956 11704 27968
rect 11756 27956 11762 28008
rect 11790 27956 11796 28008
rect 11848 27996 11854 28008
rect 12069 27999 12127 28005
rect 12069 27996 12081 27999
rect 11848 27968 12081 27996
rect 11848 27956 11854 27968
rect 12069 27965 12081 27968
rect 12115 27965 12127 27999
rect 12069 27959 12127 27965
rect 13262 27956 13268 28008
rect 13320 27996 13326 28008
rect 13541 27999 13599 28005
rect 13541 27996 13553 27999
rect 13320 27968 13553 27996
rect 13320 27956 13326 27968
rect 13541 27965 13553 27968
rect 13587 27965 13599 27999
rect 13541 27959 13599 27965
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27996 13691 27999
rect 15102 27996 15108 28008
rect 13679 27968 15108 27996
rect 13679 27965 13691 27968
rect 13633 27959 13691 27965
rect 15102 27956 15108 27968
rect 15160 27996 15166 28008
rect 15672 28005 15700 28036
rect 16758 28024 16764 28036
rect 16816 28024 16822 28076
rect 16850 28024 16856 28076
rect 16908 28064 16914 28076
rect 17957 28067 18015 28073
rect 17957 28064 17969 28067
rect 16908 28036 17969 28064
rect 16908 28024 16914 28036
rect 17957 28033 17969 28036
rect 18003 28033 18015 28067
rect 17957 28027 18015 28033
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 15160 27968 15301 27996
rect 15160 27956 15166 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 15289 27959 15347 27965
rect 15657 27999 15715 28005
rect 15657 27965 15669 27999
rect 15703 27965 15715 27999
rect 15657 27959 15715 27965
rect 16114 27956 16120 28008
rect 16172 27956 16178 28008
rect 16209 27999 16267 28005
rect 16209 27965 16221 27999
rect 16255 27965 16267 27999
rect 16209 27959 16267 27965
rect 11885 27931 11943 27937
rect 11885 27897 11897 27931
rect 11931 27928 11943 27931
rect 11974 27928 11980 27940
rect 11931 27900 11980 27928
rect 11931 27897 11943 27900
rect 11885 27891 11943 27897
rect 11974 27888 11980 27900
rect 12032 27888 12038 27940
rect 13814 27888 13820 27940
rect 13872 27888 13878 27940
rect 15378 27888 15384 27940
rect 15436 27928 15442 27940
rect 15473 27931 15531 27937
rect 15473 27928 15485 27931
rect 15436 27900 15485 27928
rect 15436 27888 15442 27900
rect 15473 27897 15485 27900
rect 15519 27897 15531 27931
rect 15473 27891 15531 27897
rect 15565 27931 15623 27937
rect 15565 27897 15577 27931
rect 15611 27897 15623 27931
rect 16224 27928 16252 27959
rect 16298 27956 16304 28008
rect 16356 27956 16362 28008
rect 16393 27999 16451 28005
rect 16393 27965 16405 27999
rect 16439 27996 16451 27999
rect 16577 27999 16635 28005
rect 16577 27996 16589 27999
rect 16439 27968 16589 27996
rect 16439 27965 16451 27968
rect 16393 27959 16451 27965
rect 16577 27965 16589 27968
rect 16623 27965 16635 27999
rect 16577 27959 16635 27965
rect 16666 27928 16672 27940
rect 16224 27900 16672 27928
rect 15565 27891 15623 27897
rect 15580 27860 15608 27891
rect 16666 27888 16672 27900
rect 16724 27928 16730 27940
rect 17310 27928 17316 27940
rect 16724 27900 17316 27928
rect 16724 27888 16730 27900
rect 17310 27888 17316 27900
rect 17368 27888 17374 27940
rect 16298 27860 16304 27872
rect 15580 27832 16304 27860
rect 16298 27820 16304 27832
rect 16356 27820 16362 27872
rect 16761 27863 16819 27869
rect 16761 27829 16773 27863
rect 16807 27860 16819 27863
rect 18064 27860 18092 28104
rect 18414 28092 18420 28104
rect 18472 28092 18478 28144
rect 21450 28092 21456 28144
rect 21508 28132 21514 28144
rect 22370 28132 22376 28144
rect 21508 28104 22376 28132
rect 21508 28092 21514 28104
rect 22370 28092 22376 28104
rect 22428 28132 22434 28144
rect 22554 28132 22560 28144
rect 22428 28104 22560 28132
rect 22428 28092 22434 28104
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 24780 28132 24808 28163
rect 24946 28160 24952 28172
rect 25004 28160 25010 28212
rect 25777 28203 25835 28209
rect 25777 28169 25789 28203
rect 25823 28200 25835 28203
rect 25866 28200 25872 28212
rect 25823 28172 25872 28200
rect 25823 28169 25835 28172
rect 25777 28163 25835 28169
rect 25866 28160 25872 28172
rect 25924 28160 25930 28212
rect 28077 28203 28135 28209
rect 28077 28169 28089 28203
rect 28123 28169 28135 28203
rect 28077 28163 28135 28169
rect 24136 28104 24808 28132
rect 19978 28024 19984 28076
rect 20036 28064 20042 28076
rect 20438 28064 20444 28076
rect 20036 28036 20444 28064
rect 20036 28024 20042 28036
rect 20438 28024 20444 28036
rect 20496 28064 20502 28076
rect 21726 28064 21732 28076
rect 20496 28036 21732 28064
rect 20496 28024 20502 28036
rect 21726 28024 21732 28036
rect 21784 28024 21790 28076
rect 18969 27999 19027 28005
rect 18969 27965 18981 27999
rect 19015 27996 19027 27999
rect 19058 27996 19064 28008
rect 19015 27968 19064 27996
rect 19015 27965 19027 27968
rect 18969 27959 19027 27965
rect 19058 27956 19064 27968
rect 19116 27956 19122 28008
rect 20898 27956 20904 28008
rect 20956 27956 20962 28008
rect 22278 27956 22284 28008
rect 22336 27956 22342 28008
rect 23750 27956 23756 28008
rect 23808 27996 23814 28008
rect 23934 27996 23940 28008
rect 23808 27968 23940 27996
rect 23808 27956 23814 27968
rect 23934 27956 23940 27968
rect 23992 27996 23998 28008
rect 24136 28005 24164 28104
rect 24854 28092 24860 28144
rect 24912 28092 24918 28144
rect 28092 28132 28120 28163
rect 28258 28160 28264 28212
rect 28316 28160 28322 28212
rect 28350 28132 28356 28144
rect 28092 28104 28356 28132
rect 28350 28092 28356 28104
rect 28408 28092 28414 28144
rect 24765 28067 24823 28073
rect 24765 28033 24777 28067
rect 24811 28064 24823 28067
rect 24872 28064 24900 28092
rect 24811 28036 24900 28064
rect 24811 28033 24823 28036
rect 24765 28027 24823 28033
rect 24029 27999 24087 28005
rect 24029 27996 24041 27999
rect 23992 27968 24041 27996
rect 23992 27956 23998 27968
rect 24029 27965 24041 27968
rect 24075 27965 24087 27999
rect 24029 27959 24087 27965
rect 24121 27999 24179 28005
rect 24121 27965 24133 27999
rect 24167 27965 24179 27999
rect 24121 27959 24179 27965
rect 24210 27956 24216 28008
rect 24268 27956 24274 28008
rect 24486 27956 24492 28008
rect 24544 27956 24550 28008
rect 24857 27999 24915 28005
rect 24857 27965 24869 27999
rect 24903 27996 24915 27999
rect 25498 27996 25504 28008
rect 24903 27968 25504 27996
rect 24903 27965 24915 27968
rect 24857 27959 24915 27965
rect 25498 27956 25504 27968
rect 25556 27956 25562 28008
rect 25774 28005 25780 28008
rect 25593 27999 25651 28005
rect 25593 27965 25605 27999
rect 25639 27965 25651 27999
rect 25593 27959 25651 27965
rect 25747 27999 25780 28005
rect 25747 27965 25759 27999
rect 25747 27959 25780 27965
rect 22830 27888 22836 27940
rect 22888 27928 22894 27940
rect 24302 27928 24308 27940
rect 24360 27937 24366 27940
rect 24360 27931 24389 27937
rect 22888 27900 24308 27928
rect 22888 27888 22894 27900
rect 24302 27888 24308 27900
rect 24377 27897 24389 27931
rect 24360 27891 24389 27897
rect 24360 27888 24366 27891
rect 16807 27832 18092 27860
rect 16807 27829 16819 27832
rect 16761 27823 16819 27829
rect 18690 27820 18696 27872
rect 18748 27860 18754 27872
rect 18877 27863 18935 27869
rect 18877 27860 18889 27863
rect 18748 27832 18889 27860
rect 18748 27820 18754 27832
rect 18877 27829 18889 27832
rect 18923 27829 18935 27863
rect 18877 27823 18935 27829
rect 22186 27820 22192 27872
rect 22244 27820 22250 27872
rect 23934 27820 23940 27872
rect 23992 27860 23998 27872
rect 24504 27860 24532 27956
rect 24581 27931 24639 27937
rect 24581 27897 24593 27931
rect 24627 27928 24639 27931
rect 24670 27928 24676 27940
rect 24627 27900 24676 27928
rect 24627 27897 24639 27900
rect 24581 27891 24639 27897
rect 24670 27888 24676 27900
rect 24728 27888 24734 27940
rect 25608 27928 25636 27959
rect 25774 27956 25780 27959
rect 25832 27956 25838 28008
rect 27614 27956 27620 28008
rect 27672 27996 27678 28008
rect 27709 27999 27767 28005
rect 27709 27996 27721 27999
rect 27672 27968 27721 27996
rect 27672 27956 27678 27968
rect 27709 27965 27721 27968
rect 27755 27965 27767 27999
rect 27709 27959 27767 27965
rect 26050 27928 26056 27940
rect 25608 27900 26056 27928
rect 26050 27888 26056 27900
rect 26108 27888 26114 27940
rect 27982 27888 27988 27940
rect 28040 27928 28046 27940
rect 28077 27931 28135 27937
rect 28077 27928 28089 27931
rect 28040 27900 28089 27928
rect 28040 27888 28046 27900
rect 28077 27897 28089 27900
rect 28123 27928 28135 27931
rect 28258 27928 28264 27940
rect 28123 27900 28264 27928
rect 28123 27897 28135 27900
rect 28077 27891 28135 27897
rect 28258 27888 28264 27900
rect 28316 27888 28322 27940
rect 23992 27832 24532 27860
rect 25041 27863 25099 27869
rect 23992 27820 23998 27832
rect 25041 27829 25053 27863
rect 25087 27860 25099 27863
rect 25130 27860 25136 27872
rect 25087 27832 25136 27860
rect 25087 27829 25099 27832
rect 25041 27823 25099 27829
rect 25130 27820 25136 27832
rect 25188 27820 25194 27872
rect 552 27770 31648 27792
rect 552 27718 4322 27770
rect 4374 27718 4386 27770
rect 4438 27718 4450 27770
rect 4502 27718 4514 27770
rect 4566 27718 4578 27770
rect 4630 27718 12096 27770
rect 12148 27718 12160 27770
rect 12212 27718 12224 27770
rect 12276 27718 12288 27770
rect 12340 27718 12352 27770
rect 12404 27718 19870 27770
rect 19922 27718 19934 27770
rect 19986 27718 19998 27770
rect 20050 27718 20062 27770
rect 20114 27718 20126 27770
rect 20178 27718 27644 27770
rect 27696 27718 27708 27770
rect 27760 27718 27772 27770
rect 27824 27718 27836 27770
rect 27888 27718 27900 27770
rect 27952 27718 31648 27770
rect 552 27696 31648 27718
rect 14369 27659 14427 27665
rect 14369 27625 14381 27659
rect 14415 27656 14427 27659
rect 14458 27656 14464 27668
rect 14415 27628 14464 27656
rect 14415 27625 14427 27628
rect 14369 27619 14427 27625
rect 14458 27616 14464 27628
rect 14516 27616 14522 27668
rect 16298 27616 16304 27668
rect 16356 27656 16362 27668
rect 18138 27656 18144 27668
rect 16356 27628 18144 27656
rect 16356 27616 16362 27628
rect 18138 27616 18144 27628
rect 18196 27616 18202 27668
rect 23290 27616 23296 27668
rect 23348 27656 23354 27668
rect 23348 27628 24624 27656
rect 23348 27616 23354 27628
rect 11885 27591 11943 27597
rect 11885 27557 11897 27591
rect 11931 27588 11943 27591
rect 15102 27588 15108 27600
rect 11931 27560 12112 27588
rect 11931 27557 11943 27560
rect 11885 27551 11943 27557
rect 11701 27523 11759 27529
rect 11701 27489 11713 27523
rect 11747 27489 11759 27523
rect 11701 27483 11759 27489
rect 11716 27452 11744 27483
rect 11790 27480 11796 27532
rect 11848 27520 11854 27532
rect 12084 27529 12112 27560
rect 13832 27560 15108 27588
rect 11977 27523 12035 27529
rect 11977 27520 11989 27523
rect 11848 27492 11989 27520
rect 11848 27480 11854 27492
rect 11977 27489 11989 27492
rect 12023 27489 12035 27523
rect 11977 27483 12035 27489
rect 12069 27523 12127 27529
rect 12069 27489 12081 27523
rect 12115 27520 12127 27523
rect 12526 27520 12532 27532
rect 12115 27492 12532 27520
rect 12115 27489 12127 27492
rect 12069 27483 12127 27489
rect 12526 27480 12532 27492
rect 12584 27520 12590 27532
rect 13262 27520 13268 27532
rect 12584 27492 13268 27520
rect 12584 27480 12590 27492
rect 13262 27480 13268 27492
rect 13320 27520 13326 27532
rect 13722 27520 13728 27532
rect 13320 27492 13728 27520
rect 13320 27480 13326 27492
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 13832 27529 13860 27560
rect 13818 27523 13876 27529
rect 13818 27489 13830 27523
rect 13864 27489 13876 27523
rect 13818 27483 13876 27489
rect 13998 27480 14004 27532
rect 14056 27480 14062 27532
rect 14476 27529 14504 27560
rect 15102 27548 15108 27560
rect 15160 27548 15166 27600
rect 16758 27548 16764 27600
rect 16816 27548 16822 27600
rect 18230 27548 18236 27600
rect 18288 27548 18294 27600
rect 21634 27548 21640 27600
rect 21692 27548 21698 27600
rect 21729 27591 21787 27597
rect 21729 27557 21741 27591
rect 21775 27588 21787 27591
rect 22189 27591 22247 27597
rect 22189 27588 22201 27591
rect 21775 27560 22201 27588
rect 21775 27557 21787 27560
rect 21729 27551 21787 27557
rect 22189 27557 22201 27560
rect 22235 27557 22247 27591
rect 22189 27551 22247 27557
rect 23658 27548 23664 27600
rect 23716 27588 23722 27600
rect 23716 27560 23888 27588
rect 23716 27548 23722 27560
rect 14093 27523 14151 27529
rect 14093 27489 14105 27523
rect 14139 27489 14151 27523
rect 14093 27483 14151 27489
rect 14231 27523 14289 27529
rect 14231 27489 14243 27523
rect 14277 27520 14289 27523
rect 14461 27523 14519 27529
rect 14277 27492 14412 27520
rect 14277 27489 14289 27492
rect 14231 27483 14289 27489
rect 12345 27455 12403 27461
rect 11716 27424 12296 27452
rect 11790 27344 11796 27396
rect 11848 27384 11854 27396
rect 12268 27393 12296 27424
rect 12345 27421 12357 27455
rect 12391 27452 12403 27455
rect 13170 27452 13176 27464
rect 12391 27424 13176 27452
rect 12391 27421 12403 27424
rect 12345 27415 12403 27421
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 12161 27387 12219 27393
rect 12161 27384 12173 27387
rect 11848 27356 12173 27384
rect 11848 27344 11854 27356
rect 12161 27353 12173 27356
rect 12207 27353 12219 27387
rect 12161 27347 12219 27353
rect 12253 27387 12311 27393
rect 12253 27353 12265 27387
rect 12299 27353 12311 27387
rect 14108 27384 14136 27483
rect 14384 27452 14412 27492
rect 14461 27489 14473 27523
rect 14507 27489 14519 27523
rect 14461 27483 14519 27489
rect 14645 27523 14703 27529
rect 14645 27489 14657 27523
rect 14691 27520 14703 27523
rect 14734 27520 14740 27532
rect 14691 27492 14740 27520
rect 14691 27489 14703 27492
rect 14645 27483 14703 27489
rect 14734 27480 14740 27492
rect 14792 27480 14798 27532
rect 16669 27523 16727 27529
rect 16669 27489 16681 27523
rect 16715 27489 16727 27523
rect 16669 27483 16727 27489
rect 16853 27523 16911 27529
rect 16853 27489 16865 27523
rect 16899 27520 16911 27523
rect 17402 27520 17408 27532
rect 16899 27492 17408 27520
rect 16899 27489 16911 27492
rect 16853 27483 16911 27489
rect 14553 27455 14611 27461
rect 14553 27452 14565 27455
rect 14384 27424 14565 27452
rect 14553 27421 14565 27424
rect 14599 27421 14611 27455
rect 14553 27415 14611 27421
rect 15378 27412 15384 27464
rect 15436 27412 15442 27464
rect 15841 27455 15899 27461
rect 15841 27421 15853 27455
rect 15887 27452 15899 27455
rect 16482 27452 16488 27464
rect 15887 27424 16488 27452
rect 15887 27421 15899 27424
rect 15841 27415 15899 27421
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 16684 27452 16712 27483
rect 17402 27480 17408 27492
rect 17460 27480 17466 27532
rect 18690 27480 18696 27532
rect 18748 27480 18754 27532
rect 18949 27523 19007 27529
rect 18949 27520 18961 27523
rect 18800 27492 18961 27520
rect 17310 27452 17316 27464
rect 16684 27424 17316 27452
rect 17310 27412 17316 27424
rect 17368 27412 17374 27464
rect 17954 27412 17960 27464
rect 18012 27412 18018 27464
rect 18141 27455 18199 27461
rect 18141 27421 18153 27455
rect 18187 27421 18199 27455
rect 18800 27452 18828 27492
rect 18949 27489 18961 27492
rect 18995 27489 19007 27523
rect 18949 27483 19007 27489
rect 20438 27480 20444 27532
rect 20496 27480 20502 27532
rect 20530 27480 20536 27532
rect 20588 27480 20594 27532
rect 20993 27523 21051 27529
rect 20993 27489 21005 27523
rect 21039 27520 21051 27523
rect 21082 27520 21088 27532
rect 21039 27492 21088 27520
rect 21039 27489 21051 27492
rect 20993 27483 21051 27489
rect 21082 27480 21088 27492
rect 21140 27480 21146 27532
rect 21545 27523 21603 27529
rect 21545 27489 21557 27523
rect 21591 27489 21603 27523
rect 21867 27523 21925 27529
rect 21867 27520 21879 27523
rect 21545 27483 21603 27489
rect 21744 27492 21879 27520
rect 18141 27415 18199 27421
rect 18616 27424 18828 27452
rect 21560 27452 21588 27483
rect 21744 27464 21772 27492
rect 21867 27489 21879 27492
rect 21913 27520 21925 27523
rect 23290 27520 23296 27532
rect 21913 27492 23296 27520
rect 21913 27489 21925 27492
rect 21867 27483 21925 27489
rect 23290 27480 23296 27492
rect 23348 27480 23354 27532
rect 23860 27529 23888 27560
rect 23845 27523 23903 27529
rect 23845 27489 23857 27523
rect 23891 27489 23903 27523
rect 23845 27483 23903 27489
rect 24026 27480 24032 27532
rect 24084 27480 24090 27532
rect 24394 27520 24400 27532
rect 24136 27492 24400 27520
rect 21560 27424 21680 27452
rect 14274 27384 14280 27396
rect 12253 27347 12311 27353
rect 12406 27356 14280 27384
rect 11330 27276 11336 27328
rect 11388 27316 11394 27328
rect 11517 27319 11575 27325
rect 11517 27316 11529 27319
rect 11388 27288 11529 27316
rect 11388 27276 11394 27288
rect 11517 27285 11529 27288
rect 11563 27285 11575 27319
rect 11517 27279 11575 27285
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 12406 27316 12434 27356
rect 14274 27344 14280 27356
rect 14332 27344 14338 27396
rect 15102 27344 15108 27396
rect 15160 27384 15166 27396
rect 15657 27387 15715 27393
rect 15657 27384 15669 27387
rect 15160 27356 15669 27384
rect 15160 27344 15166 27356
rect 15657 27353 15669 27356
rect 15703 27353 15715 27387
rect 15657 27347 15715 27353
rect 12032 27288 12434 27316
rect 18156 27316 18184 27415
rect 18616 27393 18644 27424
rect 18601 27387 18659 27393
rect 18601 27353 18613 27387
rect 18647 27353 18659 27387
rect 21652 27384 21680 27424
rect 21726 27412 21732 27464
rect 21784 27412 21790 27464
rect 22005 27455 22063 27461
rect 22005 27421 22017 27455
rect 22051 27452 22063 27455
rect 22738 27452 22744 27464
rect 22051 27424 22744 27452
rect 22051 27421 22063 27424
rect 22005 27415 22063 27421
rect 22738 27412 22744 27424
rect 22796 27412 22802 27464
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27421 22891 27455
rect 22833 27415 22891 27421
rect 22462 27384 22468 27396
rect 21652 27356 22468 27384
rect 18601 27347 18659 27353
rect 22462 27344 22468 27356
rect 22520 27344 22526 27396
rect 22554 27344 22560 27396
rect 22612 27384 22618 27396
rect 22848 27384 22876 27415
rect 23474 27412 23480 27464
rect 23532 27452 23538 27464
rect 23753 27455 23811 27461
rect 23753 27452 23765 27455
rect 23532 27424 23765 27452
rect 23532 27412 23538 27424
rect 23753 27421 23765 27424
rect 23799 27452 23811 27455
rect 24136 27452 24164 27492
rect 24394 27480 24400 27492
rect 24452 27480 24458 27532
rect 24486 27480 24492 27532
rect 24544 27480 24550 27532
rect 24596 27520 24624 27628
rect 25038 27616 25044 27668
rect 25096 27616 25102 27668
rect 27518 27659 27576 27665
rect 27518 27625 27530 27659
rect 27564 27656 27576 27659
rect 27564 27628 27844 27656
rect 27564 27625 27576 27628
rect 27518 27619 27576 27625
rect 24854 27548 24860 27600
rect 24912 27588 24918 27600
rect 25317 27591 25375 27597
rect 25317 27588 25329 27591
rect 24912 27560 25329 27588
rect 24912 27548 24918 27560
rect 25317 27557 25329 27560
rect 25363 27557 25375 27591
rect 25317 27551 25375 27557
rect 27433 27591 27491 27597
rect 27433 27557 27445 27591
rect 27479 27588 27491 27591
rect 27709 27591 27767 27597
rect 27709 27588 27721 27591
rect 27479 27560 27721 27588
rect 27479 27557 27491 27560
rect 27433 27551 27491 27557
rect 27709 27557 27721 27560
rect 27755 27557 27767 27591
rect 27816 27588 27844 27628
rect 27816 27560 28580 27588
rect 27709 27551 27767 27557
rect 24765 27523 24823 27529
rect 24765 27520 24777 27523
rect 24596 27492 24777 27520
rect 24765 27489 24777 27492
rect 24811 27489 24823 27523
rect 25041 27523 25099 27529
rect 25041 27520 25053 27523
rect 24765 27483 24823 27489
rect 24964 27492 25053 27520
rect 23799 27424 24164 27452
rect 23799 27421 23811 27424
rect 23753 27415 23811 27421
rect 24210 27412 24216 27464
rect 24268 27452 24274 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24268 27424 24593 27452
rect 24268 27412 24274 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 24670 27384 24676 27396
rect 22612 27356 24676 27384
rect 22612 27344 22618 27356
rect 24670 27344 24676 27356
rect 24728 27344 24734 27396
rect 19794 27316 19800 27328
rect 18156 27288 19800 27316
rect 12032 27276 12038 27288
rect 19794 27276 19800 27288
rect 19852 27316 19858 27328
rect 20073 27319 20131 27325
rect 20073 27316 20085 27319
rect 19852 27288 20085 27316
rect 19852 27276 19858 27288
rect 20073 27285 20085 27288
rect 20119 27285 20131 27319
rect 20073 27279 20131 27285
rect 20254 27276 20260 27328
rect 20312 27276 20318 27328
rect 20806 27276 20812 27328
rect 20864 27276 20870 27328
rect 21361 27319 21419 27325
rect 21361 27285 21373 27319
rect 21407 27316 21419 27319
rect 21450 27316 21456 27328
rect 21407 27288 21456 27316
rect 21407 27285 21419 27288
rect 21361 27279 21419 27285
rect 21450 27276 21456 27288
rect 21508 27276 21514 27328
rect 22370 27276 22376 27328
rect 22428 27316 22434 27328
rect 22738 27316 22744 27328
rect 22428 27288 22744 27316
rect 22428 27276 22434 27288
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 23014 27276 23020 27328
rect 23072 27316 23078 27328
rect 23109 27319 23167 27325
rect 23109 27316 23121 27319
rect 23072 27288 23121 27316
rect 23072 27276 23078 27288
rect 23109 27285 23121 27288
rect 23155 27285 23167 27319
rect 23109 27279 23167 27285
rect 24118 27276 24124 27328
rect 24176 27316 24182 27328
rect 24213 27319 24271 27325
rect 24213 27316 24225 27319
rect 24176 27288 24225 27316
rect 24176 27276 24182 27288
rect 24213 27285 24225 27288
rect 24259 27285 24271 27319
rect 24213 27279 24271 27285
rect 24578 27276 24584 27328
rect 24636 27276 24642 27328
rect 24780 27316 24808 27483
rect 24964 27393 24992 27492
rect 25041 27489 25053 27492
rect 25087 27489 25099 27523
rect 25041 27483 25099 27489
rect 25130 27480 25136 27532
rect 25188 27480 25194 27532
rect 25222 27480 25228 27532
rect 25280 27520 25286 27532
rect 26973 27523 27031 27529
rect 26973 27520 26985 27523
rect 25280 27492 26985 27520
rect 25280 27480 25286 27492
rect 25774 27412 25780 27464
rect 25832 27412 25838 27464
rect 24949 27387 25007 27393
rect 24949 27353 24961 27387
rect 24995 27353 25007 27387
rect 24949 27347 25007 27353
rect 25792 27316 25820 27412
rect 25866 27344 25872 27396
rect 25924 27384 25930 27396
rect 26050 27384 26056 27396
rect 25924 27356 26056 27384
rect 25924 27344 25930 27356
rect 26050 27344 26056 27356
rect 26108 27344 26114 27396
rect 26160 27384 26188 27492
rect 26973 27489 26985 27492
rect 27019 27489 27031 27523
rect 26973 27483 27031 27489
rect 27341 27523 27399 27529
rect 27341 27489 27353 27523
rect 27387 27520 27399 27523
rect 27522 27520 27528 27532
rect 27387 27492 27528 27520
rect 27387 27489 27399 27492
rect 27341 27483 27399 27489
rect 27522 27480 27528 27492
rect 27580 27480 27586 27532
rect 27617 27523 27675 27529
rect 27617 27489 27629 27523
rect 27663 27520 27675 27523
rect 28350 27520 28356 27532
rect 27663 27492 28356 27520
rect 27663 27489 27675 27492
rect 27617 27483 27675 27489
rect 28350 27480 28356 27492
rect 28408 27480 28414 27532
rect 28552 27529 28580 27560
rect 28537 27523 28595 27529
rect 28537 27489 28549 27523
rect 28583 27489 28595 27523
rect 28537 27483 28595 27489
rect 26326 27412 26332 27464
rect 26384 27452 26390 27464
rect 26384 27424 26648 27452
rect 26384 27412 26390 27424
rect 26513 27387 26571 27393
rect 26513 27384 26525 27387
rect 26160 27356 26525 27384
rect 26513 27353 26525 27356
rect 26559 27353 26571 27387
rect 26620 27384 26648 27424
rect 26694 27412 26700 27464
rect 26752 27452 26758 27464
rect 26881 27455 26939 27461
rect 26881 27452 26893 27455
rect 26752 27424 26893 27452
rect 26752 27412 26758 27424
rect 26881 27421 26893 27424
rect 26927 27421 26939 27455
rect 27540 27452 27568 27480
rect 28074 27452 28080 27464
rect 27540 27424 28080 27452
rect 26881 27415 26939 27421
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28261 27455 28319 27461
rect 28261 27421 28273 27455
rect 28307 27421 28319 27455
rect 28261 27415 28319 27421
rect 27522 27384 27528 27396
rect 26620 27356 27528 27384
rect 26513 27347 26571 27353
rect 27522 27344 27528 27356
rect 27580 27384 27586 27396
rect 28276 27384 28304 27415
rect 27580 27356 28304 27384
rect 27580 27344 27586 27356
rect 24780 27288 25820 27316
rect 26237 27319 26295 27325
rect 26237 27285 26249 27319
rect 26283 27316 26295 27319
rect 26326 27316 26332 27328
rect 26283 27288 26332 27316
rect 26283 27285 26295 27288
rect 26237 27279 26295 27285
rect 26326 27276 26332 27288
rect 26384 27276 26390 27328
rect 26418 27276 26424 27328
rect 26476 27276 26482 27328
rect 26878 27276 26884 27328
rect 26936 27316 26942 27328
rect 27065 27319 27123 27325
rect 27065 27316 27077 27319
rect 26936 27288 27077 27316
rect 26936 27276 26942 27288
rect 27065 27285 27077 27288
rect 27111 27285 27123 27319
rect 27065 27279 27123 27285
rect 29086 27276 29092 27328
rect 29144 27276 29150 27328
rect 552 27226 31648 27248
rect 552 27174 3662 27226
rect 3714 27174 3726 27226
rect 3778 27174 3790 27226
rect 3842 27174 3854 27226
rect 3906 27174 3918 27226
rect 3970 27174 11436 27226
rect 11488 27174 11500 27226
rect 11552 27174 11564 27226
rect 11616 27174 11628 27226
rect 11680 27174 11692 27226
rect 11744 27174 19210 27226
rect 19262 27174 19274 27226
rect 19326 27174 19338 27226
rect 19390 27174 19402 27226
rect 19454 27174 19466 27226
rect 19518 27174 26984 27226
rect 27036 27174 27048 27226
rect 27100 27174 27112 27226
rect 27164 27174 27176 27226
rect 27228 27174 27240 27226
rect 27292 27174 31648 27226
rect 552 27152 31648 27174
rect 12526 27072 12532 27124
rect 12584 27072 12590 27124
rect 13998 27072 14004 27124
rect 14056 27112 14062 27124
rect 14553 27115 14611 27121
rect 14553 27112 14565 27115
rect 14056 27084 14565 27112
rect 14056 27072 14062 27084
rect 14553 27081 14565 27084
rect 14599 27081 14611 27115
rect 14553 27075 14611 27081
rect 20714 27072 20720 27124
rect 20772 27112 20778 27124
rect 21085 27115 21143 27121
rect 21085 27112 21097 27115
rect 20772 27084 21097 27112
rect 20772 27072 20778 27084
rect 21085 27081 21097 27084
rect 21131 27112 21143 27115
rect 24210 27112 24216 27124
rect 21131 27084 24216 27112
rect 21131 27081 21143 27084
rect 21085 27075 21143 27081
rect 24210 27072 24216 27084
rect 24268 27112 24274 27124
rect 26142 27112 26148 27124
rect 24268 27084 26148 27112
rect 24268 27072 24274 27084
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 26326 27072 26332 27124
rect 26384 27072 26390 27124
rect 26418 27072 26424 27124
rect 26476 27072 26482 27124
rect 26786 27072 26792 27124
rect 26844 27072 26850 27124
rect 14369 27047 14427 27053
rect 14369 27013 14381 27047
rect 14415 27044 14427 27047
rect 17770 27044 17776 27056
rect 14415 27016 17776 27044
rect 14415 27013 14427 27016
rect 14369 27007 14427 27013
rect 17770 27004 17776 27016
rect 17828 27004 17834 27056
rect 24946 27004 24952 27056
rect 25004 27044 25010 27056
rect 25869 27047 25927 27053
rect 25869 27044 25881 27047
rect 25004 27016 25881 27044
rect 25004 27004 25010 27016
rect 25869 27013 25881 27016
rect 25915 27044 25927 27047
rect 25915 27016 26924 27044
rect 25915 27013 25927 27016
rect 25869 27007 25927 27013
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26976 11023 26979
rect 11149 26979 11207 26985
rect 11149 26976 11161 26979
rect 11011 26948 11161 26976
rect 11011 26945 11023 26948
rect 10965 26939 11023 26945
rect 11149 26945 11161 26948
rect 11195 26945 11207 26979
rect 19521 26979 19579 26985
rect 11149 26939 11207 26945
rect 14292 26948 14780 26976
rect 14292 26920 14320 26948
rect 11057 26911 11115 26917
rect 11057 26877 11069 26911
rect 11103 26908 11115 26911
rect 11238 26908 11244 26920
rect 11103 26880 11244 26908
rect 11103 26877 11115 26880
rect 11057 26871 11115 26877
rect 11238 26868 11244 26880
rect 11296 26868 11302 26920
rect 11422 26917 11428 26920
rect 11416 26908 11428 26917
rect 11383 26880 11428 26908
rect 11416 26871 11428 26880
rect 11422 26868 11428 26871
rect 11480 26868 11486 26920
rect 13722 26868 13728 26920
rect 13780 26908 13786 26920
rect 14185 26911 14243 26917
rect 14185 26908 14197 26911
rect 13780 26880 14197 26908
rect 13780 26868 13786 26880
rect 14185 26877 14197 26880
rect 14231 26877 14243 26911
rect 14185 26871 14243 26877
rect 14274 26868 14280 26920
rect 14332 26868 14338 26920
rect 14550 26868 14556 26920
rect 14608 26868 14614 26920
rect 14752 26917 14780 26948
rect 19521 26945 19533 26979
rect 19567 26976 19579 26979
rect 19705 26979 19763 26985
rect 19705 26976 19717 26979
rect 19567 26948 19717 26976
rect 19567 26945 19579 26948
rect 19521 26939 19579 26945
rect 19705 26945 19717 26948
rect 19751 26945 19763 26979
rect 19705 26939 19763 26945
rect 22462 26936 22468 26988
rect 22520 26976 22526 26988
rect 25961 26979 26019 26985
rect 22520 26948 22968 26976
rect 22520 26936 22526 26948
rect 14737 26911 14795 26917
rect 14737 26877 14749 26911
rect 14783 26877 14795 26911
rect 14737 26871 14795 26877
rect 17034 26868 17040 26920
rect 17092 26908 17098 26920
rect 17497 26911 17555 26917
rect 17497 26908 17509 26911
rect 17092 26880 17509 26908
rect 17092 26868 17098 26880
rect 17497 26877 17509 26880
rect 17543 26877 17555 26911
rect 17497 26871 17555 26877
rect 17954 26868 17960 26920
rect 18012 26908 18018 26920
rect 18233 26911 18291 26917
rect 18233 26908 18245 26911
rect 18012 26880 18245 26908
rect 18012 26868 18018 26880
rect 18233 26877 18245 26880
rect 18279 26877 18291 26911
rect 18233 26871 18291 26877
rect 18506 26868 18512 26920
rect 18564 26908 18570 26920
rect 19245 26911 19303 26917
rect 19245 26908 19257 26911
rect 18564 26880 19257 26908
rect 18564 26868 18570 26880
rect 19245 26877 19257 26880
rect 19291 26877 19303 26911
rect 19245 26871 19303 26877
rect 19610 26868 19616 26920
rect 19668 26868 19674 26920
rect 19972 26911 20030 26917
rect 19972 26877 19984 26911
rect 20018 26908 20030 26911
rect 20254 26908 20260 26920
rect 20018 26880 20260 26908
rect 20018 26877 20030 26880
rect 19972 26871 20030 26877
rect 20254 26868 20260 26880
rect 20312 26868 20318 26920
rect 21174 26868 21180 26920
rect 21232 26868 21238 26920
rect 21450 26917 21456 26920
rect 21444 26908 21456 26917
rect 21411 26880 21456 26908
rect 21444 26871 21456 26880
rect 21450 26868 21456 26871
rect 21508 26868 21514 26920
rect 22738 26868 22744 26920
rect 22796 26908 22802 26920
rect 22940 26917 22968 26948
rect 25961 26945 25973 26979
rect 26007 26976 26019 26979
rect 26513 26979 26571 26985
rect 26513 26976 26525 26979
rect 26007 26948 26525 26976
rect 26007 26945 26019 26948
rect 25961 26939 26019 26945
rect 26513 26945 26525 26948
rect 26559 26945 26571 26979
rect 26513 26939 26571 26945
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 22796 26880 22845 26908
rect 22796 26868 22802 26880
rect 22833 26877 22845 26880
rect 22879 26877 22891 26911
rect 22833 26871 22891 26877
rect 22925 26911 22983 26917
rect 22925 26877 22937 26911
rect 22971 26877 22983 26911
rect 22925 26871 22983 26877
rect 23014 26868 23020 26920
rect 23072 26868 23078 26920
rect 23290 26868 23296 26920
rect 23348 26868 23354 26920
rect 23382 26868 23388 26920
rect 23440 26908 23446 26920
rect 24118 26917 24124 26920
rect 23477 26911 23535 26917
rect 23477 26908 23489 26911
rect 23440 26880 23489 26908
rect 23440 26868 23446 26880
rect 23477 26877 23489 26880
rect 23523 26877 23535 26911
rect 23477 26871 23535 26877
rect 23569 26911 23627 26917
rect 23569 26877 23581 26911
rect 23615 26908 23627 26911
rect 23845 26911 23903 26917
rect 23845 26908 23857 26911
rect 23615 26880 23857 26908
rect 23615 26877 23627 26880
rect 23569 26871 23627 26877
rect 23845 26877 23857 26880
rect 23891 26877 23903 26911
rect 24112 26908 24124 26917
rect 24079 26880 24124 26908
rect 23845 26871 23903 26877
rect 24112 26871 24124 26880
rect 24118 26868 24124 26871
rect 24176 26868 24182 26920
rect 24394 26868 24400 26920
rect 24452 26908 24458 26920
rect 25222 26908 25228 26920
rect 24452 26880 25228 26908
rect 24452 26868 24458 26880
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 25314 26868 25320 26920
rect 25372 26908 25378 26920
rect 26050 26908 26056 26920
rect 25372 26880 26056 26908
rect 25372 26868 25378 26880
rect 26050 26868 26056 26880
rect 26108 26868 26114 26920
rect 26237 26911 26295 26917
rect 26237 26877 26249 26911
rect 26283 26908 26295 26911
rect 26326 26908 26332 26920
rect 26283 26880 26332 26908
rect 26283 26877 26295 26880
rect 26237 26871 26295 26877
rect 26326 26868 26332 26880
rect 26384 26868 26390 26920
rect 26896 26917 26924 27016
rect 28813 26979 28871 26985
rect 28813 26945 28825 26979
rect 28859 26976 28871 26979
rect 29089 26979 29147 26985
rect 29089 26976 29101 26979
rect 28859 26948 29101 26976
rect 28859 26945 28871 26948
rect 28813 26939 28871 26945
rect 29089 26945 29101 26948
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 26881 26911 26939 26917
rect 26881 26877 26893 26911
rect 26927 26877 26939 26911
rect 26881 26871 26939 26877
rect 27982 26868 27988 26920
rect 28040 26908 28046 26920
rect 28997 26911 29055 26917
rect 28997 26908 29009 26911
rect 28040 26880 29009 26908
rect 28040 26868 28046 26880
rect 28997 26877 29009 26880
rect 29043 26877 29055 26911
rect 28997 26871 29055 26877
rect 14461 26843 14519 26849
rect 14461 26840 14473 26843
rect 14200 26812 14473 26840
rect 14200 26784 14228 26812
rect 14461 26809 14473 26812
rect 14507 26809 14519 26843
rect 14461 26803 14519 26809
rect 20530 26800 20536 26852
rect 20588 26840 20594 26852
rect 22370 26840 22376 26852
rect 20588 26812 22376 26840
rect 20588 26800 20594 26812
rect 22370 26800 22376 26812
rect 22428 26800 22434 26852
rect 23135 26843 23193 26849
rect 23135 26840 23147 26843
rect 22480 26812 23147 26840
rect 13906 26732 13912 26784
rect 13964 26772 13970 26784
rect 14182 26772 14188 26784
rect 13964 26744 14188 26772
rect 13964 26732 13970 26744
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 16942 26732 16948 26784
rect 17000 26732 17006 26784
rect 17494 26732 17500 26784
rect 17552 26772 17558 26784
rect 17681 26775 17739 26781
rect 17681 26772 17693 26775
rect 17552 26744 17693 26772
rect 17552 26732 17558 26744
rect 17681 26741 17693 26744
rect 17727 26741 17739 26775
rect 17681 26735 17739 26741
rect 18322 26732 18328 26784
rect 18380 26772 18386 26784
rect 18693 26775 18751 26781
rect 18693 26772 18705 26775
rect 18380 26744 18705 26772
rect 18380 26732 18386 26744
rect 18693 26741 18705 26744
rect 18739 26741 18751 26775
rect 18693 26735 18751 26741
rect 20990 26732 20996 26784
rect 21048 26772 21054 26784
rect 22002 26772 22008 26784
rect 21048 26744 22008 26772
rect 21048 26732 21054 26744
rect 22002 26732 22008 26744
rect 22060 26772 22066 26784
rect 22480 26772 22508 26812
rect 23135 26809 23147 26812
rect 23181 26809 23193 26843
rect 23135 26803 23193 26809
rect 22060 26744 22508 26772
rect 22060 26732 22066 26744
rect 22554 26732 22560 26784
rect 22612 26732 22618 26784
rect 22646 26732 22652 26784
rect 22704 26732 22710 26784
rect 22738 26732 22744 26784
rect 22796 26772 22802 26784
rect 23308 26772 23336 26868
rect 25501 26843 25559 26849
rect 25501 26809 25513 26843
rect 25547 26840 25559 26843
rect 26510 26840 26516 26852
rect 25547 26812 26516 26840
rect 25547 26809 25559 26812
rect 25501 26803 25559 26809
rect 26510 26800 26516 26812
rect 26568 26800 26574 26852
rect 28442 26840 28448 26852
rect 26620 26812 28448 26840
rect 22796 26744 23336 26772
rect 22796 26732 22802 26744
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 24578 26772 24584 26784
rect 23624 26744 24584 26772
rect 23624 26732 23630 26744
rect 24578 26732 24584 26744
rect 24636 26772 24642 26784
rect 24762 26772 24768 26784
rect 24636 26744 24768 26772
rect 24636 26732 24642 26744
rect 24762 26732 24768 26744
rect 24820 26732 24826 26784
rect 25225 26775 25283 26781
rect 25225 26741 25237 26775
rect 25271 26772 25283 26775
rect 25406 26772 25412 26784
rect 25271 26744 25412 26772
rect 25271 26741 25283 26744
rect 25225 26735 25283 26741
rect 25406 26732 25412 26744
rect 25464 26732 25470 26784
rect 25866 26732 25872 26784
rect 25924 26772 25930 26784
rect 26620 26772 26648 26812
rect 28442 26800 28448 26812
rect 28500 26800 28506 26852
rect 28568 26843 28626 26849
rect 28568 26809 28580 26843
rect 28614 26840 28626 26843
rect 29086 26840 29092 26852
rect 28614 26812 29092 26840
rect 28614 26809 28626 26812
rect 28568 26803 28626 26809
rect 29086 26800 29092 26812
rect 29144 26800 29150 26852
rect 25924 26744 26648 26772
rect 25924 26732 25930 26744
rect 26694 26732 26700 26784
rect 26752 26772 26758 26784
rect 26973 26775 27031 26781
rect 26973 26772 26985 26775
rect 26752 26744 26985 26772
rect 26752 26732 26758 26744
rect 26973 26741 26985 26744
rect 27019 26741 27031 26775
rect 26973 26735 27031 26741
rect 27433 26775 27491 26781
rect 27433 26741 27445 26775
rect 27479 26772 27491 26775
rect 27522 26772 27528 26784
rect 27479 26744 27528 26772
rect 27479 26741 27491 26744
rect 27433 26735 27491 26741
rect 27522 26732 27528 26744
rect 27580 26732 27586 26784
rect 552 26682 31648 26704
rect 552 26630 4322 26682
rect 4374 26630 4386 26682
rect 4438 26630 4450 26682
rect 4502 26630 4514 26682
rect 4566 26630 4578 26682
rect 4630 26630 12096 26682
rect 12148 26630 12160 26682
rect 12212 26630 12224 26682
rect 12276 26630 12288 26682
rect 12340 26630 12352 26682
rect 12404 26630 19870 26682
rect 19922 26630 19934 26682
rect 19986 26630 19998 26682
rect 20050 26630 20062 26682
rect 20114 26630 20126 26682
rect 20178 26630 27644 26682
rect 27696 26630 27708 26682
rect 27760 26630 27772 26682
rect 27824 26630 27836 26682
rect 27888 26630 27900 26682
rect 27952 26630 31648 26682
rect 552 26608 31648 26630
rect 13814 26528 13820 26580
rect 13872 26568 13878 26580
rect 14461 26571 14519 26577
rect 14461 26568 14473 26571
rect 13872 26540 14473 26568
rect 13872 26528 13878 26540
rect 14461 26537 14473 26540
rect 14507 26537 14519 26571
rect 14461 26531 14519 26537
rect 14734 26528 14740 26580
rect 14792 26528 14798 26580
rect 17034 26528 17040 26580
rect 17092 26528 17098 26580
rect 17310 26528 17316 26580
rect 17368 26568 17374 26580
rect 17405 26571 17463 26577
rect 17405 26568 17417 26571
rect 17368 26540 17417 26568
rect 17368 26528 17374 26540
rect 17405 26537 17417 26540
rect 17451 26537 17463 26571
rect 17405 26531 17463 26537
rect 17494 26528 17500 26580
rect 17552 26528 17558 26580
rect 18138 26528 18144 26580
rect 18196 26568 18202 26580
rect 18233 26571 18291 26577
rect 18233 26568 18245 26571
rect 18196 26540 18245 26568
rect 18196 26528 18202 26540
rect 18233 26537 18245 26540
rect 18279 26537 18291 26571
rect 18233 26531 18291 26537
rect 18322 26528 18328 26580
rect 18380 26528 18386 26580
rect 18414 26528 18420 26580
rect 18472 26568 18478 26580
rect 19061 26571 19119 26577
rect 19061 26568 19073 26571
rect 18472 26540 19073 26568
rect 18472 26528 18478 26540
rect 19061 26537 19073 26540
rect 19107 26537 19119 26571
rect 19061 26531 19119 26537
rect 19702 26528 19708 26580
rect 19760 26528 19766 26580
rect 20257 26571 20315 26577
rect 20257 26537 20269 26571
rect 20303 26568 20315 26571
rect 20438 26568 20444 26580
rect 20303 26540 20444 26568
rect 20303 26537 20315 26540
rect 20257 26531 20315 26537
rect 20438 26528 20444 26540
rect 20496 26528 20502 26580
rect 20548 26540 21128 26568
rect 15105 26503 15163 26509
rect 15105 26469 15117 26503
rect 15151 26500 15163 26503
rect 15286 26500 15292 26512
rect 15151 26472 15292 26500
rect 15151 26469 15163 26472
rect 15105 26463 15163 26469
rect 15286 26460 15292 26472
rect 15344 26460 15350 26512
rect 18432 26472 19288 26500
rect 16758 26392 16764 26444
rect 16816 26392 16822 26444
rect 12618 26324 12624 26376
rect 12676 26324 12682 26376
rect 12802 26324 12808 26376
rect 12860 26324 12866 26376
rect 13170 26324 13176 26376
rect 13228 26364 13234 26376
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 13228 26336 13553 26364
rect 13228 26324 13234 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13630 26324 13636 26376
rect 13688 26373 13694 26376
rect 13688 26367 13716 26373
rect 13704 26333 13716 26367
rect 13688 26327 13716 26333
rect 13817 26367 13875 26373
rect 13817 26333 13829 26367
rect 13863 26364 13875 26367
rect 14182 26364 14188 26376
rect 13863 26336 14188 26364
rect 13863 26333 13875 26336
rect 13817 26327 13875 26333
rect 13688 26324 13694 26327
rect 14182 26324 14188 26336
rect 14240 26324 14246 26376
rect 15194 26324 15200 26376
rect 15252 26324 15258 26376
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26333 15347 26367
rect 15289 26327 15347 26333
rect 17681 26367 17739 26373
rect 17681 26333 17693 26367
rect 17727 26364 17739 26367
rect 18046 26364 18052 26376
rect 17727 26336 18052 26364
rect 17727 26333 17739 26336
rect 17681 26327 17739 26333
rect 13265 26299 13323 26305
rect 13265 26265 13277 26299
rect 13311 26296 13323 26299
rect 15304 26296 15332 26327
rect 18046 26324 18052 26336
rect 18104 26364 18110 26376
rect 18432 26373 18460 26472
rect 19260 26373 19288 26472
rect 19610 26460 19616 26512
rect 19668 26500 19674 26512
rect 20346 26500 20352 26512
rect 19668 26472 20352 26500
rect 19668 26460 19674 26472
rect 20346 26460 20352 26472
rect 20404 26500 20410 26512
rect 20548 26500 20576 26540
rect 20404 26472 20576 26500
rect 20404 26460 20410 26472
rect 20438 26392 20444 26444
rect 20496 26392 20502 26444
rect 20533 26435 20591 26441
rect 20533 26401 20545 26435
rect 20579 26401 20591 26435
rect 20533 26395 20591 26401
rect 20625 26435 20683 26441
rect 20625 26401 20637 26435
rect 20671 26401 20683 26435
rect 20625 26395 20683 26401
rect 20763 26435 20821 26441
rect 20763 26401 20775 26435
rect 20809 26432 20821 26435
rect 20990 26432 20996 26444
rect 20809 26404 20996 26432
rect 20809 26401 20821 26404
rect 20763 26395 20821 26401
rect 18417 26367 18475 26373
rect 18417 26364 18429 26367
rect 18104 26336 18429 26364
rect 18104 26324 18110 26336
rect 18417 26333 18429 26336
rect 18463 26333 18475 26367
rect 18417 26327 18475 26333
rect 19153 26367 19211 26373
rect 19153 26333 19165 26367
rect 19199 26333 19211 26367
rect 19153 26327 19211 26333
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26333 19303 26367
rect 19245 26327 19303 26333
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26333 19947 26367
rect 19889 26327 19947 26333
rect 13311 26268 13400 26296
rect 13311 26265 13323 26268
rect 13265 26259 13323 26265
rect 13372 26228 13400 26268
rect 15120 26268 15332 26296
rect 13906 26228 13912 26240
rect 13372 26200 13912 26228
rect 13906 26188 13912 26200
rect 13964 26228 13970 26240
rect 15010 26228 15016 26240
rect 13964 26200 15016 26228
rect 13964 26188 13970 26200
rect 15010 26188 15016 26200
rect 15068 26228 15074 26240
rect 15120 26228 15148 26268
rect 18138 26256 18144 26308
rect 18196 26296 18202 26308
rect 18196 26268 18828 26296
rect 18196 26256 18202 26268
rect 15068 26200 15148 26228
rect 15068 26188 15074 26200
rect 16574 26188 16580 26240
rect 16632 26228 16638 26240
rect 16669 26231 16727 26237
rect 16669 26228 16681 26231
rect 16632 26200 16681 26228
rect 16632 26188 16638 26200
rect 16669 26197 16681 26200
rect 16715 26197 16727 26231
rect 16669 26191 16727 26197
rect 17862 26188 17868 26240
rect 17920 26188 17926 26240
rect 18690 26188 18696 26240
rect 18748 26188 18754 26240
rect 18800 26228 18828 26268
rect 19058 26256 19064 26308
rect 19116 26296 19122 26308
rect 19168 26296 19196 26327
rect 19536 26296 19564 26327
rect 19904 26296 19932 26327
rect 19116 26268 19564 26296
rect 19628 26268 19932 26296
rect 20548 26296 20576 26395
rect 20640 26364 20668 26395
rect 20990 26392 20996 26404
rect 21048 26392 21054 26444
rect 21100 26432 21128 26540
rect 21174 26528 21180 26580
rect 21232 26568 21238 26580
rect 21361 26571 21419 26577
rect 21361 26568 21373 26571
rect 21232 26540 21373 26568
rect 21232 26528 21238 26540
rect 21361 26537 21373 26540
rect 21407 26537 21419 26571
rect 22278 26568 22284 26580
rect 21361 26531 21419 26537
rect 21468 26540 22284 26568
rect 21468 26441 21496 26540
rect 22278 26528 22284 26540
rect 22336 26568 22342 26580
rect 23106 26568 23112 26580
rect 22336 26540 23112 26568
rect 22336 26528 22342 26540
rect 23106 26528 23112 26540
rect 23164 26568 23170 26580
rect 23290 26568 23296 26580
rect 23164 26540 23296 26568
rect 23164 26528 23170 26540
rect 23290 26528 23296 26540
rect 23348 26528 23354 26580
rect 24026 26528 24032 26580
rect 24084 26568 24090 26580
rect 24121 26571 24179 26577
rect 24121 26568 24133 26571
rect 24084 26540 24133 26568
rect 24084 26528 24090 26540
rect 24121 26537 24133 26540
rect 24167 26537 24179 26571
rect 24121 26531 24179 26537
rect 26602 26528 26608 26580
rect 26660 26568 26666 26580
rect 27065 26571 27123 26577
rect 27065 26568 27077 26571
rect 26660 26540 27077 26568
rect 26660 26528 26666 26540
rect 27065 26537 27077 26540
rect 27111 26537 27123 26571
rect 28166 26568 28172 26580
rect 27065 26531 27123 26537
rect 28000 26540 28172 26568
rect 22186 26500 22192 26512
rect 21744 26472 22192 26500
rect 21744 26441 21772 26472
rect 22186 26460 22192 26472
rect 22244 26460 22250 26512
rect 22646 26460 22652 26512
rect 22704 26460 22710 26512
rect 22830 26460 22836 26512
rect 22888 26500 22894 26512
rect 23615 26503 23673 26509
rect 23615 26500 23627 26503
rect 22888 26472 23627 26500
rect 22888 26460 22894 26472
rect 23615 26469 23627 26472
rect 23661 26469 23673 26503
rect 23615 26463 23673 26469
rect 23845 26503 23903 26509
rect 23845 26469 23857 26503
rect 23891 26500 23903 26503
rect 24486 26500 24492 26512
rect 23891 26472 24492 26500
rect 23891 26469 23903 26472
rect 23845 26463 23903 26469
rect 24486 26460 24492 26472
rect 24544 26500 24550 26512
rect 25498 26500 25504 26512
rect 24544 26472 25504 26500
rect 24544 26460 24550 26472
rect 25498 26460 25504 26472
rect 25556 26460 25562 26512
rect 26694 26460 26700 26512
rect 26752 26460 26758 26512
rect 26786 26460 26792 26512
rect 26844 26460 26850 26512
rect 27617 26503 27675 26509
rect 27617 26469 27629 26503
rect 27663 26500 27675 26503
rect 27706 26500 27712 26512
rect 27663 26472 27712 26500
rect 27663 26469 27675 26472
rect 27617 26463 27675 26469
rect 27706 26460 27712 26472
rect 27764 26460 27770 26512
rect 27833 26503 27891 26509
rect 27833 26469 27845 26503
rect 27879 26500 27891 26503
rect 28000 26500 28028 26540
rect 28166 26528 28172 26540
rect 28224 26528 28230 26580
rect 28350 26528 28356 26580
rect 28408 26528 28414 26580
rect 27879 26472 28028 26500
rect 27879 26469 27891 26472
rect 27833 26463 27891 26469
rect 21453 26435 21511 26441
rect 21453 26432 21465 26435
rect 21100 26404 21465 26432
rect 21453 26401 21465 26404
rect 21499 26401 21511 26435
rect 21453 26395 21511 26401
rect 21729 26435 21787 26441
rect 21729 26401 21741 26435
rect 21775 26401 21787 26435
rect 21729 26395 21787 26401
rect 21996 26435 22054 26441
rect 21996 26401 22008 26435
rect 22042 26432 22054 26435
rect 22664 26432 22692 26460
rect 22042 26404 22692 26432
rect 22042 26401 22054 26404
rect 21996 26395 22054 26401
rect 23382 26392 23388 26444
rect 23440 26432 23446 26444
rect 23753 26435 23811 26441
rect 23753 26432 23765 26435
rect 23440 26404 23765 26432
rect 23440 26392 23446 26404
rect 23753 26401 23765 26404
rect 23799 26401 23811 26435
rect 23753 26395 23811 26401
rect 23937 26435 23995 26441
rect 23937 26401 23949 26435
rect 23983 26401 23995 26435
rect 23937 26395 23995 26401
rect 20640 26336 20852 26364
rect 20824 26308 20852 26336
rect 20898 26324 20904 26376
rect 20956 26324 20962 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26364 23535 26367
rect 23566 26364 23572 26376
rect 23523 26336 23572 26364
rect 23523 26333 23535 26336
rect 23477 26327 23535 26333
rect 23566 26324 23572 26336
rect 23624 26324 23630 26376
rect 20714 26296 20720 26308
rect 20548 26268 20720 26296
rect 19116 26256 19122 26268
rect 18874 26228 18880 26240
rect 18800 26200 18880 26228
rect 18874 26188 18880 26200
rect 18932 26228 18938 26240
rect 19628 26228 19656 26268
rect 20714 26256 20720 26268
rect 20772 26256 20778 26308
rect 20806 26256 20812 26308
rect 20864 26296 20870 26308
rect 21634 26296 21640 26308
rect 20864 26268 21640 26296
rect 20864 26256 20870 26268
rect 21634 26256 21640 26268
rect 21692 26256 21698 26308
rect 18932 26200 19656 26228
rect 18932 26188 18938 26200
rect 19794 26188 19800 26240
rect 19852 26228 19858 26240
rect 19889 26231 19947 26237
rect 19889 26228 19901 26231
rect 19852 26200 19901 26228
rect 19852 26188 19858 26200
rect 19889 26197 19901 26200
rect 19935 26197 19947 26231
rect 19889 26191 19947 26197
rect 23109 26231 23167 26237
rect 23109 26197 23121 26231
rect 23155 26228 23167 26231
rect 23474 26228 23480 26240
rect 23155 26200 23480 26228
rect 23155 26197 23167 26200
rect 23109 26191 23167 26197
rect 23474 26188 23480 26200
rect 23532 26188 23538 26240
rect 23566 26188 23572 26240
rect 23624 26228 23630 26240
rect 23750 26228 23756 26240
rect 23624 26200 23756 26228
rect 23624 26188 23630 26200
rect 23750 26188 23756 26200
rect 23808 26228 23814 26240
rect 23952 26228 23980 26395
rect 26326 26392 26332 26444
rect 26384 26392 26390 26444
rect 26418 26392 26424 26444
rect 26476 26392 26482 26444
rect 26510 26392 26516 26444
rect 26568 26432 26574 26444
rect 26568 26404 26613 26432
rect 26568 26392 26574 26404
rect 26344 26364 26372 26392
rect 26804 26364 26832 26460
rect 26878 26392 26884 26444
rect 26936 26441 26942 26444
rect 26936 26432 26944 26441
rect 26936 26404 26981 26432
rect 26936 26395 26944 26404
rect 26936 26392 26942 26395
rect 27522 26392 27528 26444
rect 27580 26432 27586 26444
rect 28077 26435 28135 26441
rect 28077 26432 28089 26435
rect 27580 26404 28089 26432
rect 27580 26392 27586 26404
rect 28077 26401 28089 26404
rect 28123 26401 28135 26435
rect 28077 26395 28135 26401
rect 28169 26435 28227 26441
rect 28169 26401 28181 26435
rect 28215 26401 28227 26435
rect 28169 26395 28227 26401
rect 27890 26364 27896 26376
rect 26344 26336 26740 26364
rect 26804 26336 27896 26364
rect 26050 26256 26056 26308
rect 26108 26296 26114 26308
rect 26326 26296 26332 26308
rect 26108 26268 26332 26296
rect 26108 26256 26114 26268
rect 26326 26256 26332 26268
rect 26384 26256 26390 26308
rect 26712 26296 26740 26336
rect 27890 26324 27896 26336
rect 27948 26324 27954 26376
rect 28184 26364 28212 26395
rect 28092 26336 28212 26364
rect 28092 26308 28120 26336
rect 28258 26324 28264 26376
rect 28316 26364 28322 26376
rect 28353 26367 28411 26373
rect 28353 26364 28365 26367
rect 28316 26336 28365 26364
rect 28316 26324 28322 26336
rect 28353 26333 28365 26336
rect 28399 26333 28411 26367
rect 28353 26327 28411 26333
rect 26786 26296 26792 26308
rect 26712 26268 26792 26296
rect 26786 26256 26792 26268
rect 26844 26256 26850 26308
rect 27985 26299 28043 26305
rect 27985 26265 27997 26299
rect 28031 26296 28043 26299
rect 28074 26296 28080 26308
rect 28031 26268 28080 26296
rect 28031 26265 28043 26268
rect 27985 26259 28043 26265
rect 28074 26256 28080 26268
rect 28132 26256 28138 26308
rect 28166 26256 28172 26308
rect 28224 26296 28230 26308
rect 28442 26296 28448 26308
rect 28224 26268 28448 26296
rect 28224 26256 28230 26268
rect 28442 26256 28448 26268
rect 28500 26256 28506 26308
rect 23808 26200 23980 26228
rect 27801 26231 27859 26237
rect 23808 26188 23814 26200
rect 27801 26197 27813 26231
rect 27847 26228 27859 26231
rect 28902 26228 28908 26240
rect 27847 26200 28908 26228
rect 27847 26197 27859 26200
rect 27801 26191 27859 26197
rect 28902 26188 28908 26200
rect 28960 26188 28966 26240
rect 552 26138 31648 26160
rect 552 26086 3662 26138
rect 3714 26086 3726 26138
rect 3778 26086 3790 26138
rect 3842 26086 3854 26138
rect 3906 26086 3918 26138
rect 3970 26086 11436 26138
rect 11488 26086 11500 26138
rect 11552 26086 11564 26138
rect 11616 26086 11628 26138
rect 11680 26086 11692 26138
rect 11744 26086 19210 26138
rect 19262 26086 19274 26138
rect 19326 26086 19338 26138
rect 19390 26086 19402 26138
rect 19454 26086 19466 26138
rect 19518 26086 26984 26138
rect 27036 26086 27048 26138
rect 27100 26086 27112 26138
rect 27164 26086 27176 26138
rect 27228 26086 27240 26138
rect 27292 26086 31648 26138
rect 552 26064 31648 26086
rect 12986 25984 12992 26036
rect 13044 25984 13050 26036
rect 14461 26027 14519 26033
rect 14461 25993 14473 26027
rect 14507 26024 14519 26027
rect 14550 26024 14556 26036
rect 14507 25996 14556 26024
rect 14507 25993 14519 25996
rect 14461 25987 14519 25993
rect 14550 25984 14556 25996
rect 14608 25984 14614 26036
rect 15286 25984 15292 26036
rect 15344 25984 15350 26036
rect 15378 25984 15384 26036
rect 15436 26024 15442 26036
rect 15841 26027 15899 26033
rect 15841 26024 15853 26027
rect 15436 25996 15853 26024
rect 15436 25984 15442 25996
rect 15841 25993 15853 25996
rect 15887 25993 15899 26027
rect 16758 26024 16764 26036
rect 15841 25987 15899 25993
rect 16224 25996 16764 26024
rect 13004 25956 13032 25984
rect 13357 25959 13415 25965
rect 13004 25928 13308 25956
rect 12618 25848 12624 25900
rect 12676 25888 12682 25900
rect 12989 25891 13047 25897
rect 12989 25888 13001 25891
rect 12676 25860 13001 25888
rect 12676 25848 12682 25860
rect 12989 25857 13001 25860
rect 13035 25857 13047 25891
rect 13280 25888 13308 25928
rect 13357 25925 13369 25959
rect 13403 25956 13415 25959
rect 13403 25928 15884 25956
rect 13403 25925 13415 25928
rect 13357 25919 13415 25925
rect 13541 25891 13599 25897
rect 13541 25888 13553 25891
rect 13280 25860 13553 25888
rect 12989 25851 13047 25857
rect 13541 25857 13553 25860
rect 13587 25888 13599 25891
rect 13630 25888 13636 25900
rect 13587 25860 13636 25888
rect 13587 25857 13599 25860
rect 13541 25851 13599 25857
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 15010 25848 15016 25900
rect 15068 25848 15074 25900
rect 15381 25891 15439 25897
rect 15381 25888 15393 25891
rect 15120 25860 15393 25888
rect 11330 25780 11336 25832
rect 11388 25820 11394 25832
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 11388 25792 12173 25820
rect 11388 25780 11394 25792
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 12802 25780 12808 25832
rect 12860 25820 12866 25832
rect 12897 25823 12955 25829
rect 12897 25820 12909 25823
rect 12860 25792 12909 25820
rect 12860 25780 12866 25792
rect 12897 25789 12909 25792
rect 12943 25789 12955 25823
rect 12897 25783 12955 25789
rect 13170 25780 13176 25832
rect 13228 25780 13234 25832
rect 15120 25820 15148 25860
rect 15381 25857 15393 25860
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 14752 25792 15148 25820
rect 11882 25644 11888 25696
rect 11940 25684 11946 25696
rect 12069 25687 12127 25693
rect 12069 25684 12081 25687
rect 11940 25656 12081 25684
rect 11940 25644 11946 25656
rect 12069 25653 12081 25656
rect 12115 25653 12127 25687
rect 12069 25647 12127 25653
rect 14182 25644 14188 25696
rect 14240 25644 14246 25696
rect 14274 25644 14280 25696
rect 14332 25684 14338 25696
rect 14752 25684 14780 25792
rect 15194 25780 15200 25832
rect 15252 25820 15258 25832
rect 15565 25823 15623 25829
rect 15565 25820 15577 25823
rect 15252 25792 15577 25820
rect 15252 25780 15258 25792
rect 15565 25789 15577 25792
rect 15611 25820 15623 25823
rect 15746 25820 15752 25832
rect 15611 25792 15752 25820
rect 15611 25789 15623 25792
rect 15565 25783 15623 25789
rect 15746 25780 15752 25792
rect 15804 25780 15810 25832
rect 15856 25829 15884 25928
rect 16224 25829 16252 25996
rect 16758 25984 16764 25996
rect 16816 26024 16822 26036
rect 17126 26024 17132 26036
rect 16816 25996 17132 26024
rect 16816 25984 16822 25996
rect 17126 25984 17132 25996
rect 17184 26024 17190 26036
rect 17184 25996 18276 26024
rect 17184 25984 17190 25996
rect 17770 25916 17776 25968
rect 17828 25956 17834 25968
rect 17828 25928 18092 25956
rect 17828 25916 17834 25928
rect 17954 25848 17960 25900
rect 18012 25848 18018 25900
rect 15841 25823 15899 25829
rect 15841 25789 15853 25823
rect 15887 25789 15899 25823
rect 15841 25783 15899 25789
rect 16025 25823 16083 25829
rect 16025 25789 16037 25823
rect 16071 25789 16083 25823
rect 16025 25783 16083 25789
rect 16209 25823 16267 25829
rect 16209 25789 16221 25823
rect 16255 25789 16267 25823
rect 16209 25783 16267 25789
rect 16485 25823 16543 25829
rect 16485 25789 16497 25823
rect 16531 25820 16543 25823
rect 16574 25820 16580 25832
rect 16531 25792 16580 25820
rect 16531 25789 16543 25792
rect 16485 25783 16543 25789
rect 14829 25755 14887 25761
rect 14829 25721 14841 25755
rect 14875 25752 14887 25755
rect 15289 25755 15347 25761
rect 15289 25752 15301 25755
rect 14875 25724 15301 25752
rect 14875 25721 14887 25724
rect 14829 25715 14887 25721
rect 15289 25721 15301 25724
rect 15335 25752 15347 25755
rect 15470 25752 15476 25764
rect 15335 25724 15476 25752
rect 15335 25721 15347 25724
rect 15289 25715 15347 25721
rect 15470 25712 15476 25724
rect 15528 25712 15534 25764
rect 16040 25752 16068 25783
rect 16574 25780 16580 25792
rect 16632 25780 16638 25832
rect 16752 25823 16810 25829
rect 16752 25789 16764 25823
rect 16798 25820 16810 25823
rect 17862 25820 17868 25832
rect 16798 25792 17868 25820
rect 16798 25789 16810 25792
rect 16752 25783 16810 25789
rect 17862 25780 17868 25792
rect 17920 25780 17926 25832
rect 18064 25820 18092 25928
rect 18248 25888 18276 25996
rect 18506 25984 18512 26036
rect 18564 25984 18570 26036
rect 20349 26027 20407 26033
rect 20349 25993 20361 26027
rect 20395 26024 20407 26027
rect 20990 26024 20996 26036
rect 20395 25996 20996 26024
rect 20395 25993 20407 25996
rect 20349 25987 20407 25993
rect 20990 25984 20996 25996
rect 21048 25984 21054 26036
rect 28810 25888 28816 25900
rect 18248 25860 18920 25888
rect 18892 25829 18920 25860
rect 27908 25860 28816 25888
rect 27908 25832 27936 25860
rect 28810 25848 28816 25860
rect 28868 25848 28874 25900
rect 18325 25823 18383 25829
rect 18325 25820 18337 25823
rect 18064 25792 18337 25820
rect 18325 25789 18337 25792
rect 18371 25789 18383 25823
rect 18325 25783 18383 25789
rect 18877 25823 18935 25829
rect 18877 25789 18889 25823
rect 18923 25789 18935 25823
rect 18877 25783 18935 25789
rect 19058 25780 19064 25832
rect 19116 25780 19122 25832
rect 19245 25823 19303 25829
rect 19245 25789 19257 25823
rect 19291 25789 19303 25823
rect 19245 25783 19303 25789
rect 18506 25752 18512 25764
rect 15764 25724 16068 25752
rect 17880 25724 18512 25752
rect 15764 25693 15792 25724
rect 14921 25687 14979 25693
rect 14921 25684 14933 25687
rect 14332 25656 14933 25684
rect 14332 25644 14338 25656
rect 14921 25653 14933 25656
rect 14967 25653 14979 25687
rect 14921 25647 14979 25653
rect 15749 25687 15807 25693
rect 15749 25653 15761 25687
rect 15795 25653 15807 25687
rect 15749 25647 15807 25653
rect 16301 25687 16359 25693
rect 16301 25653 16313 25687
rect 16347 25684 16359 25687
rect 16482 25684 16488 25696
rect 16347 25656 16488 25684
rect 16347 25653 16359 25656
rect 16301 25647 16359 25653
rect 16482 25644 16488 25656
rect 16540 25644 16546 25696
rect 17880 25693 17908 25724
rect 18506 25712 18512 25724
rect 18564 25712 18570 25764
rect 18966 25712 18972 25764
rect 19024 25752 19030 25764
rect 19260 25752 19288 25783
rect 19794 25780 19800 25832
rect 19852 25780 19858 25832
rect 27890 25780 27896 25832
rect 27948 25780 27954 25832
rect 28074 25780 28080 25832
rect 28132 25820 28138 25832
rect 28169 25823 28227 25829
rect 28169 25820 28181 25823
rect 28132 25792 28181 25820
rect 28132 25780 28138 25792
rect 28169 25789 28181 25792
rect 28215 25789 28227 25823
rect 28169 25783 28227 25789
rect 19024 25724 19288 25752
rect 27709 25755 27767 25761
rect 19024 25712 19030 25724
rect 27709 25721 27721 25755
rect 27755 25752 27767 25755
rect 27755 25724 28212 25752
rect 27755 25721 27767 25724
rect 27709 25715 27767 25721
rect 28184 25696 28212 25724
rect 17865 25687 17923 25693
rect 17865 25653 17877 25687
rect 17911 25653 17923 25687
rect 17865 25647 17923 25653
rect 18138 25644 18144 25696
rect 18196 25644 18202 25696
rect 18322 25644 18328 25696
rect 18380 25684 18386 25696
rect 18785 25687 18843 25693
rect 18785 25684 18797 25687
rect 18380 25656 18797 25684
rect 18380 25644 18386 25656
rect 18785 25653 18797 25656
rect 18831 25653 18843 25687
rect 18785 25647 18843 25653
rect 21358 25644 21364 25696
rect 21416 25684 21422 25696
rect 23198 25684 23204 25696
rect 21416 25656 23204 25684
rect 21416 25644 21422 25656
rect 23198 25644 23204 25656
rect 23256 25644 23262 25696
rect 27522 25644 27528 25696
rect 27580 25684 27586 25696
rect 28077 25687 28135 25693
rect 28077 25684 28089 25687
rect 27580 25656 28089 25684
rect 27580 25644 27586 25656
rect 28077 25653 28089 25656
rect 28123 25653 28135 25687
rect 28077 25647 28135 25653
rect 28166 25644 28172 25696
rect 28224 25644 28230 25696
rect 552 25594 31648 25616
rect 552 25542 4322 25594
rect 4374 25542 4386 25594
rect 4438 25542 4450 25594
rect 4502 25542 4514 25594
rect 4566 25542 4578 25594
rect 4630 25542 12096 25594
rect 12148 25542 12160 25594
rect 12212 25542 12224 25594
rect 12276 25542 12288 25594
rect 12340 25542 12352 25594
rect 12404 25542 19870 25594
rect 19922 25542 19934 25594
rect 19986 25542 19998 25594
rect 20050 25542 20062 25594
rect 20114 25542 20126 25594
rect 20178 25542 27644 25594
rect 27696 25542 27708 25594
rect 27760 25542 27772 25594
rect 27824 25542 27836 25594
rect 27888 25542 27900 25594
rect 27952 25542 31648 25594
rect 552 25520 31648 25542
rect 13170 25440 13176 25492
rect 13228 25480 13234 25492
rect 13265 25483 13323 25489
rect 13265 25480 13277 25483
rect 13228 25452 13277 25480
rect 13228 25440 13234 25452
rect 13265 25449 13277 25452
rect 13311 25449 13323 25483
rect 13265 25443 13323 25449
rect 17865 25483 17923 25489
rect 17865 25449 17877 25483
rect 17911 25480 17923 25483
rect 17954 25480 17960 25492
rect 17911 25452 17960 25480
rect 17911 25449 17923 25452
rect 17865 25443 17923 25449
rect 11882 25304 11888 25356
rect 11940 25304 11946 25356
rect 12152 25347 12210 25353
rect 12152 25313 12164 25347
rect 12198 25344 12210 25347
rect 13078 25344 13084 25356
rect 12198 25316 13084 25344
rect 12198 25313 12210 25316
rect 12152 25307 12210 25313
rect 13078 25304 13084 25316
rect 13136 25304 13142 25356
rect 13280 25344 13308 25443
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 24213 25483 24271 25489
rect 24213 25449 24225 25483
rect 24259 25480 24271 25483
rect 24854 25480 24860 25492
rect 24259 25452 24860 25480
rect 24259 25449 24271 25452
rect 24213 25443 24271 25449
rect 24854 25440 24860 25452
rect 24912 25440 24918 25492
rect 25685 25483 25743 25489
rect 25685 25449 25697 25483
rect 25731 25480 25743 25483
rect 26418 25480 26424 25492
rect 25731 25452 26424 25480
rect 25731 25449 25743 25452
rect 25685 25443 25743 25449
rect 26418 25440 26424 25452
rect 26476 25440 26482 25492
rect 14182 25372 14188 25424
rect 14240 25412 14246 25424
rect 14553 25415 14611 25421
rect 14553 25412 14565 25415
rect 14240 25384 14565 25412
rect 14240 25372 14246 25384
rect 14553 25381 14565 25384
rect 14599 25381 14611 25415
rect 14553 25375 14611 25381
rect 14737 25415 14795 25421
rect 14737 25381 14749 25415
rect 14783 25412 14795 25415
rect 14829 25415 14887 25421
rect 14829 25412 14841 25415
rect 14783 25384 14841 25412
rect 14783 25381 14795 25384
rect 14737 25375 14795 25381
rect 14829 25381 14841 25384
rect 14875 25412 14887 25415
rect 15194 25412 15200 25424
rect 14875 25384 15200 25412
rect 14875 25381 14887 25384
rect 14829 25375 14887 25381
rect 15194 25372 15200 25384
rect 15252 25372 15258 25424
rect 16752 25415 16810 25421
rect 16752 25381 16764 25415
rect 16798 25412 16810 25415
rect 16942 25412 16948 25424
rect 16798 25384 16948 25412
rect 16798 25381 16810 25384
rect 16752 25375 16810 25381
rect 16942 25372 16948 25384
rect 17000 25372 17006 25424
rect 18592 25415 18650 25421
rect 18592 25381 18604 25415
rect 18638 25412 18650 25415
rect 18690 25412 18696 25424
rect 18638 25384 18696 25412
rect 18638 25381 18650 25384
rect 18592 25375 18650 25381
rect 18690 25372 18696 25384
rect 18748 25372 18754 25424
rect 21634 25372 21640 25424
rect 21692 25412 21698 25424
rect 22741 25415 22799 25421
rect 22741 25412 22753 25415
rect 21692 25384 22753 25412
rect 21692 25372 21698 25384
rect 22741 25381 22753 25384
rect 22787 25412 22799 25415
rect 23382 25412 23388 25424
rect 22787 25384 23388 25412
rect 22787 25381 22799 25384
rect 22741 25375 22799 25381
rect 23382 25372 23388 25384
rect 23440 25372 23446 25424
rect 24118 25412 24124 25424
rect 23860 25384 24124 25412
rect 13633 25347 13691 25353
rect 13633 25344 13645 25347
rect 13280 25316 13645 25344
rect 13633 25313 13645 25316
rect 13679 25313 13691 25347
rect 13633 25307 13691 25313
rect 15013 25347 15071 25353
rect 15013 25313 15025 25347
rect 15059 25344 15071 25347
rect 15289 25347 15347 25353
rect 15289 25344 15301 25347
rect 15059 25316 15301 25344
rect 15059 25313 15071 25316
rect 15013 25307 15071 25313
rect 15289 25313 15301 25316
rect 15335 25313 15347 25347
rect 15289 25307 15347 25313
rect 16206 25304 16212 25356
rect 16264 25344 16270 25356
rect 16393 25347 16451 25353
rect 16393 25344 16405 25347
rect 16264 25316 16405 25344
rect 16264 25304 16270 25316
rect 16393 25313 16405 25316
rect 16439 25313 16451 25347
rect 16393 25307 16451 25313
rect 16482 25304 16488 25356
rect 16540 25304 16546 25356
rect 18322 25304 18328 25356
rect 18380 25304 18386 25356
rect 20346 25304 20352 25356
rect 20404 25344 20410 25356
rect 20533 25347 20591 25353
rect 20533 25344 20545 25347
rect 20404 25316 20545 25344
rect 20404 25304 20410 25316
rect 20533 25313 20545 25316
rect 20579 25313 20591 25347
rect 20533 25307 20591 25313
rect 22189 25347 22247 25353
rect 22189 25313 22201 25347
rect 22235 25344 22247 25347
rect 22278 25344 22284 25356
rect 22235 25316 22284 25344
rect 22235 25313 22247 25316
rect 22189 25307 22247 25313
rect 22278 25304 22284 25316
rect 22336 25304 22342 25356
rect 22557 25347 22615 25353
rect 22557 25313 22569 25347
rect 22603 25313 22615 25347
rect 22557 25307 22615 25313
rect 22649 25347 22707 25353
rect 22649 25313 22661 25347
rect 22695 25313 22707 25347
rect 22649 25307 22707 25313
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 15933 25279 15991 25285
rect 15933 25276 15945 25279
rect 15436 25248 15945 25276
rect 15436 25236 15442 25248
rect 15933 25245 15945 25248
rect 15979 25276 15991 25279
rect 16022 25276 16028 25288
rect 15979 25248 16028 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16022 25236 16028 25248
rect 16080 25236 16086 25288
rect 21450 25236 21456 25288
rect 21508 25276 21514 25288
rect 22572 25276 22600 25307
rect 21508 25248 22600 25276
rect 21508 25236 21514 25248
rect 13998 25168 14004 25220
rect 14056 25208 14062 25220
rect 14369 25211 14427 25217
rect 14369 25208 14381 25211
rect 14056 25180 14381 25208
rect 14056 25168 14062 25180
rect 14369 25177 14381 25180
rect 14415 25177 14427 25211
rect 14369 25171 14427 25177
rect 14277 25143 14335 25149
rect 14277 25109 14289 25143
rect 14323 25140 14335 25143
rect 14642 25140 14648 25152
rect 14323 25112 14648 25140
rect 14323 25109 14335 25112
rect 14277 25103 14335 25109
rect 14642 25100 14648 25112
rect 14700 25100 14706 25152
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 15562 25140 15568 25152
rect 15243 25112 15568 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 15562 25100 15568 25112
rect 15620 25100 15626 25152
rect 16206 25100 16212 25152
rect 16264 25100 16270 25152
rect 19058 25100 19064 25152
rect 19116 25140 19122 25152
rect 19705 25143 19763 25149
rect 19705 25140 19717 25143
rect 19116 25112 19717 25140
rect 19116 25100 19122 25112
rect 19705 25109 19717 25112
rect 19751 25109 19763 25143
rect 19705 25103 19763 25109
rect 20254 25100 20260 25152
rect 20312 25140 20318 25152
rect 20441 25143 20499 25149
rect 20441 25140 20453 25143
rect 20312 25112 20453 25140
rect 20312 25100 20318 25112
rect 20441 25109 20453 25112
rect 20487 25109 20499 25143
rect 20441 25103 20499 25109
rect 22094 25100 22100 25152
rect 22152 25100 22158 25152
rect 22370 25100 22376 25152
rect 22428 25100 22434 25152
rect 22572 25140 22600 25248
rect 22664 25208 22692 25307
rect 22830 25304 22836 25356
rect 22888 25353 22894 25356
rect 22888 25347 22917 25353
rect 22905 25344 22917 25347
rect 23247 25347 23305 25353
rect 23247 25344 23259 25347
rect 22905 25316 23259 25344
rect 22905 25313 22917 25316
rect 22888 25307 22917 25313
rect 23247 25313 23259 25316
rect 23293 25313 23305 25347
rect 23247 25307 23305 25313
rect 22888 25304 22894 25307
rect 23474 25304 23480 25356
rect 23532 25304 23538 25356
rect 23566 25304 23572 25356
rect 23624 25304 23630 25356
rect 23860 25353 23888 25384
rect 24118 25372 24124 25384
rect 24176 25372 24182 25424
rect 24581 25415 24639 25421
rect 24581 25381 24593 25415
rect 24627 25412 24639 25415
rect 25222 25412 25228 25424
rect 24627 25384 25228 25412
rect 24627 25381 24639 25384
rect 24581 25375 24639 25381
rect 25222 25372 25228 25384
rect 25280 25412 25286 25424
rect 25317 25415 25375 25421
rect 25317 25412 25329 25415
rect 25280 25384 25329 25412
rect 25280 25372 25286 25384
rect 25317 25381 25329 25384
rect 25363 25381 25375 25415
rect 25317 25375 25375 25381
rect 25409 25415 25467 25421
rect 25409 25381 25421 25415
rect 25455 25412 25467 25415
rect 26142 25412 26148 25424
rect 25455 25384 26148 25412
rect 25455 25381 25467 25384
rect 25409 25375 25467 25381
rect 26142 25372 26148 25384
rect 26200 25372 26206 25424
rect 23845 25347 23903 25353
rect 23845 25313 23857 25347
rect 23891 25313 23903 25347
rect 24489 25347 24547 25353
rect 24489 25344 24501 25347
rect 23845 25307 23903 25313
rect 23952 25316 24501 25344
rect 23014 25236 23020 25288
rect 23072 25236 23078 25288
rect 23109 25279 23167 25285
rect 23109 25245 23121 25279
rect 23155 25276 23167 25279
rect 23492 25276 23520 25304
rect 23952 25285 23980 25316
rect 24489 25313 24501 25316
rect 24535 25313 24547 25347
rect 24489 25307 24547 25313
rect 25133 25347 25191 25353
rect 25133 25313 25145 25347
rect 25179 25344 25191 25347
rect 25501 25347 25559 25353
rect 25179 25316 25360 25344
rect 25179 25313 25191 25316
rect 25133 25307 25191 25313
rect 25332 25288 25360 25316
rect 25501 25313 25513 25347
rect 25547 25313 25559 25347
rect 25501 25307 25559 25313
rect 27709 25347 27767 25353
rect 27709 25313 27721 25347
rect 27755 25344 27767 25347
rect 27982 25344 27988 25356
rect 27755 25316 27988 25344
rect 27755 25313 27767 25316
rect 27709 25307 27767 25313
rect 23937 25279 23995 25285
rect 23937 25276 23949 25279
rect 23155 25248 23244 25276
rect 23492 25248 23949 25276
rect 23155 25245 23167 25248
rect 23109 25239 23167 25245
rect 23216 25220 23244 25248
rect 23937 25245 23949 25248
rect 23983 25245 23995 25279
rect 23937 25239 23995 25245
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 22922 25208 22928 25220
rect 22664 25180 22928 25208
rect 22922 25168 22928 25180
rect 22980 25168 22986 25220
rect 23198 25168 23204 25220
rect 23256 25168 23262 25220
rect 24486 25168 24492 25220
rect 24544 25208 24550 25220
rect 24670 25208 24676 25220
rect 24544 25180 24676 25208
rect 24544 25168 24550 25180
rect 24670 25168 24676 25180
rect 24728 25208 24734 25220
rect 25516 25208 25544 25307
rect 27982 25304 27988 25316
rect 28040 25344 28046 25356
rect 28626 25344 28632 25356
rect 28040 25316 28632 25344
rect 28040 25304 28046 25316
rect 28626 25304 28632 25316
rect 28684 25304 28690 25356
rect 24728 25180 25544 25208
rect 24728 25168 24734 25180
rect 23566 25140 23572 25152
rect 22572 25112 23572 25140
rect 23566 25100 23572 25112
rect 23624 25100 23630 25152
rect 23750 25100 23756 25152
rect 23808 25100 23814 25152
rect 24026 25100 24032 25152
rect 24084 25140 24090 25152
rect 24854 25140 24860 25152
rect 24084 25112 24860 25140
rect 24084 25100 24090 25112
rect 24854 25100 24860 25112
rect 24912 25100 24918 25152
rect 27614 25100 27620 25152
rect 27672 25100 27678 25152
rect 552 25050 31648 25072
rect 552 24998 3662 25050
rect 3714 24998 3726 25050
rect 3778 24998 3790 25050
rect 3842 24998 3854 25050
rect 3906 24998 3918 25050
rect 3970 24998 11436 25050
rect 11488 24998 11500 25050
rect 11552 24998 11564 25050
rect 11616 24998 11628 25050
rect 11680 24998 11692 25050
rect 11744 24998 19210 25050
rect 19262 24998 19274 25050
rect 19326 24998 19338 25050
rect 19390 24998 19402 25050
rect 19454 24998 19466 25050
rect 19518 24998 26984 25050
rect 27036 24998 27048 25050
rect 27100 24998 27112 25050
rect 27164 24998 27176 25050
rect 27228 24998 27240 25050
rect 27292 24998 31648 25050
rect 552 24976 31648 24998
rect 12986 24896 12992 24948
rect 13044 24896 13050 24948
rect 16022 24896 16028 24948
rect 16080 24896 16086 24948
rect 21726 24896 21732 24948
rect 21784 24936 21790 24948
rect 22830 24936 22836 24948
rect 21784 24908 22836 24936
rect 21784 24896 21790 24908
rect 22830 24896 22836 24908
rect 22888 24896 22894 24948
rect 22922 24896 22928 24948
rect 22980 24936 22986 24948
rect 23293 24939 23351 24945
rect 23293 24936 23305 24939
rect 22980 24908 23305 24936
rect 22980 24896 22986 24908
rect 23293 24905 23305 24908
rect 23339 24936 23351 24939
rect 24026 24936 24032 24948
rect 23339 24908 24032 24936
rect 23339 24905 23351 24908
rect 23293 24899 23351 24905
rect 24026 24896 24032 24908
rect 24084 24896 24090 24948
rect 27249 24939 27307 24945
rect 27249 24905 27261 24939
rect 27295 24936 27307 24939
rect 27430 24936 27436 24948
rect 27295 24908 27436 24936
rect 27295 24905 27307 24908
rect 27249 24899 27307 24905
rect 27430 24896 27436 24908
rect 27488 24896 27494 24948
rect 28810 24896 28816 24948
rect 28868 24896 28874 24948
rect 17954 24868 17960 24880
rect 17788 24840 17960 24868
rect 13832 24772 14780 24800
rect 13832 24744 13860 24772
rect 11330 24692 11336 24744
rect 11388 24692 11394 24744
rect 11425 24735 11483 24741
rect 11425 24701 11437 24735
rect 11471 24732 11483 24735
rect 11609 24735 11667 24741
rect 11609 24732 11621 24735
rect 11471 24704 11621 24732
rect 11471 24701 11483 24704
rect 11425 24695 11483 24701
rect 11609 24701 11621 24704
rect 11655 24701 11667 24735
rect 11609 24695 11667 24701
rect 13814 24692 13820 24744
rect 13872 24692 13878 24744
rect 13906 24692 13912 24744
rect 13964 24692 13970 24744
rect 13998 24692 14004 24744
rect 14056 24692 14062 24744
rect 14185 24735 14243 24741
rect 14185 24701 14197 24735
rect 14231 24732 14243 24735
rect 14231 24704 14320 24732
rect 14231 24701 14243 24704
rect 14185 24695 14243 24701
rect 11876 24667 11934 24673
rect 11876 24633 11888 24667
rect 11922 24664 11934 24667
rect 13541 24667 13599 24673
rect 13541 24664 13553 24667
rect 11922 24636 13553 24664
rect 11922 24633 11934 24636
rect 11876 24627 11934 24633
rect 13541 24633 13553 24636
rect 13587 24633 13599 24667
rect 13541 24627 13599 24633
rect 13722 24556 13728 24608
rect 13780 24596 13786 24608
rect 14292 24596 14320 24704
rect 14366 24692 14372 24744
rect 14424 24692 14430 24744
rect 14461 24735 14519 24741
rect 14461 24701 14473 24735
rect 14507 24732 14519 24735
rect 14645 24735 14703 24741
rect 14645 24732 14657 24735
rect 14507 24704 14657 24732
rect 14507 24701 14519 24704
rect 14461 24695 14519 24701
rect 14645 24701 14657 24704
rect 14691 24701 14703 24735
rect 14752 24732 14780 24772
rect 17678 24760 17684 24812
rect 17736 24760 17742 24812
rect 17788 24809 17816 24840
rect 17954 24828 17960 24840
rect 18012 24828 18018 24880
rect 24857 24871 24915 24877
rect 24857 24837 24869 24871
rect 24903 24868 24915 24871
rect 26602 24868 26608 24880
rect 24903 24840 26608 24868
rect 24903 24837 24915 24840
rect 24857 24831 24915 24837
rect 26602 24828 26608 24840
rect 26660 24828 26666 24880
rect 17773 24803 17831 24809
rect 17773 24769 17785 24803
rect 17819 24769 17831 24803
rect 17773 24763 17831 24769
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24769 18107 24803
rect 18049 24763 18107 24769
rect 18233 24803 18291 24809
rect 18233 24769 18245 24803
rect 18279 24800 18291 24803
rect 18506 24800 18512 24812
rect 18279 24772 18512 24800
rect 18279 24769 18291 24772
rect 18233 24763 18291 24769
rect 14752 24704 16620 24732
rect 14645 24695 14703 24701
rect 14912 24667 14970 24673
rect 14912 24633 14924 24667
rect 14958 24664 14970 24667
rect 15010 24664 15016 24676
rect 14958 24636 15016 24664
rect 14958 24633 14970 24636
rect 14912 24627 14970 24633
rect 15010 24624 15016 24636
rect 15068 24624 15074 24676
rect 16592 24664 16620 24704
rect 17954 24692 17960 24744
rect 18012 24732 18018 24744
rect 18064 24732 18092 24763
rect 18506 24760 18512 24772
rect 18564 24760 18570 24812
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19024 24772 19288 24800
rect 19024 24760 19030 24772
rect 18984 24732 19012 24760
rect 18012 24704 19012 24732
rect 18012 24692 18018 24704
rect 19058 24692 19064 24744
rect 19116 24692 19122 24744
rect 19260 24741 19288 24772
rect 20254 24760 20260 24812
rect 20312 24760 20318 24812
rect 24486 24760 24492 24812
rect 24544 24760 24550 24812
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24800 25835 24803
rect 25823 24772 26924 24800
rect 25823 24769 25835 24772
rect 25777 24763 25835 24769
rect 19245 24735 19303 24741
rect 19245 24701 19257 24735
rect 19291 24701 19303 24735
rect 19245 24695 19303 24701
rect 19794 24692 19800 24744
rect 19852 24692 19858 24744
rect 21913 24735 21971 24741
rect 21913 24701 21925 24735
rect 21959 24732 21971 24735
rect 22002 24732 22008 24744
rect 21959 24704 22008 24732
rect 21959 24701 21971 24704
rect 21913 24695 21971 24701
rect 22002 24692 22008 24704
rect 22060 24692 22066 24744
rect 23106 24692 23112 24744
rect 23164 24732 23170 24744
rect 23385 24735 23443 24741
rect 23385 24732 23397 24735
rect 23164 24704 23397 24732
rect 23164 24692 23170 24704
rect 23385 24701 23397 24704
rect 23431 24701 23443 24735
rect 23385 24695 23443 24701
rect 23750 24692 23756 24744
rect 23808 24732 23814 24744
rect 24029 24735 24087 24741
rect 24029 24732 24041 24735
rect 23808 24704 24041 24732
rect 23808 24692 23814 24704
rect 24029 24701 24041 24704
rect 24075 24701 24087 24735
rect 24029 24695 24087 24701
rect 24213 24735 24271 24741
rect 24213 24701 24225 24735
rect 24259 24701 24271 24735
rect 24213 24695 24271 24701
rect 20254 24664 20260 24676
rect 16592 24636 20260 24664
rect 20254 24624 20260 24636
rect 20312 24624 20318 24676
rect 20346 24624 20352 24676
rect 20404 24664 20410 24676
rect 20502 24667 20560 24673
rect 20502 24664 20514 24667
rect 20404 24636 20514 24664
rect 20404 24624 20410 24636
rect 20502 24633 20514 24636
rect 20548 24633 20560 24667
rect 21726 24664 21732 24676
rect 20502 24627 20560 24633
rect 21560 24636 21732 24664
rect 15286 24596 15292 24608
rect 13780 24568 15292 24596
rect 13780 24556 13786 24568
rect 15286 24556 15292 24568
rect 15344 24596 15350 24608
rect 16206 24596 16212 24608
rect 15344 24568 16212 24596
rect 15344 24556 15350 24568
rect 16206 24556 16212 24568
rect 16264 24556 16270 24608
rect 19981 24599 20039 24605
rect 19981 24565 19993 24599
rect 20027 24596 20039 24599
rect 21560 24596 21588 24636
rect 21726 24624 21732 24636
rect 21784 24624 21790 24676
rect 22180 24667 22238 24673
rect 22180 24633 22192 24667
rect 22226 24664 22238 24667
rect 22278 24664 22284 24676
rect 22226 24636 22284 24664
rect 22226 24633 22238 24636
rect 22180 24627 22238 24633
rect 22278 24624 22284 24636
rect 22336 24624 22342 24676
rect 23658 24624 23664 24676
rect 23716 24664 23722 24676
rect 24228 24664 24256 24695
rect 25038 24692 25044 24744
rect 25096 24692 25102 24744
rect 25222 24692 25228 24744
rect 25280 24692 25286 24744
rect 25314 24692 25320 24744
rect 25372 24692 25378 24744
rect 25409 24735 25467 24741
rect 25409 24701 25421 24735
rect 25455 24732 25467 24735
rect 25498 24732 25504 24744
rect 25455 24704 25504 24732
rect 25455 24701 25467 24704
rect 25409 24695 25467 24701
rect 25498 24692 25504 24704
rect 25556 24692 25562 24744
rect 25590 24692 25596 24744
rect 25648 24692 25654 24744
rect 25869 24735 25927 24741
rect 25869 24732 25881 24735
rect 25700 24704 25881 24732
rect 23716 24636 24256 24664
rect 23716 24624 23722 24636
rect 24670 24624 24676 24676
rect 24728 24664 24734 24676
rect 25700 24664 25728 24704
rect 25869 24701 25881 24704
rect 25915 24701 25927 24735
rect 25869 24695 25927 24701
rect 26050 24692 26056 24744
rect 26108 24692 26114 24744
rect 26145 24735 26203 24741
rect 26145 24701 26157 24735
rect 26191 24701 26203 24735
rect 26145 24695 26203 24701
rect 26237 24735 26295 24741
rect 26237 24701 26249 24735
rect 26283 24701 26295 24735
rect 26237 24695 26295 24701
rect 26421 24735 26479 24741
rect 26421 24701 26433 24735
rect 26467 24732 26479 24735
rect 26786 24732 26792 24744
rect 26467 24704 26792 24732
rect 26467 24701 26479 24704
rect 26421 24695 26479 24701
rect 24728 24636 25728 24664
rect 24728 24624 24734 24636
rect 25774 24624 25780 24676
rect 25832 24664 25838 24676
rect 26160 24664 26188 24695
rect 25832 24636 26188 24664
rect 25832 24624 25838 24636
rect 20027 24568 21588 24596
rect 20027 24565 20039 24568
rect 19981 24559 20039 24565
rect 21634 24556 21640 24608
rect 21692 24556 21698 24608
rect 22462 24556 22468 24608
rect 22520 24596 22526 24608
rect 23014 24596 23020 24608
rect 22520 24568 23020 24596
rect 22520 24556 22526 24568
rect 23014 24556 23020 24568
rect 23072 24556 23078 24608
rect 23474 24556 23480 24608
rect 23532 24556 23538 24608
rect 23750 24556 23756 24608
rect 23808 24596 23814 24608
rect 23845 24599 23903 24605
rect 23845 24596 23857 24599
rect 23808 24568 23857 24596
rect 23808 24556 23814 24568
rect 23845 24565 23857 24568
rect 23891 24565 23903 24599
rect 23845 24559 23903 24565
rect 24949 24599 25007 24605
rect 24949 24565 24961 24599
rect 24995 24596 25007 24599
rect 25406 24596 25412 24608
rect 24995 24568 25412 24596
rect 24995 24565 25007 24568
rect 24949 24559 25007 24565
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 26252 24596 26280 24695
rect 26786 24692 26792 24704
rect 26844 24692 26850 24744
rect 26896 24741 26924 24772
rect 26881 24735 26939 24741
rect 26881 24701 26893 24735
rect 26927 24701 26939 24735
rect 26881 24695 26939 24701
rect 27433 24735 27491 24741
rect 27433 24701 27445 24735
rect 27479 24732 27491 24735
rect 27522 24732 27528 24744
rect 27479 24704 27528 24732
rect 27479 24701 27491 24704
rect 27433 24695 27491 24701
rect 27522 24692 27528 24704
rect 27580 24692 27586 24744
rect 26326 24624 26332 24676
rect 26384 24664 26390 24676
rect 26694 24664 26700 24676
rect 26384 24636 26700 24664
rect 26384 24624 26390 24636
rect 26694 24624 26700 24636
rect 26752 24624 26758 24676
rect 27678 24667 27736 24673
rect 27678 24664 27690 24667
rect 27540 24636 27690 24664
rect 27540 24608 27568 24636
rect 27678 24633 27690 24636
rect 27724 24633 27736 24667
rect 27678 24627 27736 24633
rect 26418 24596 26424 24608
rect 26252 24568 26424 24596
rect 26418 24556 26424 24568
rect 26476 24556 26482 24608
rect 26605 24599 26663 24605
rect 26605 24565 26617 24599
rect 26651 24596 26663 24599
rect 26973 24599 27031 24605
rect 26973 24596 26985 24599
rect 26651 24568 26985 24596
rect 26651 24565 26663 24568
rect 26605 24559 26663 24565
rect 26973 24565 26985 24568
rect 27019 24565 27031 24599
rect 26973 24559 27031 24565
rect 27062 24556 27068 24608
rect 27120 24556 27126 24608
rect 27522 24556 27528 24608
rect 27580 24556 27586 24608
rect 552 24506 31648 24528
rect 552 24454 4322 24506
rect 4374 24454 4386 24506
rect 4438 24454 4450 24506
rect 4502 24454 4514 24506
rect 4566 24454 4578 24506
rect 4630 24454 12096 24506
rect 12148 24454 12160 24506
rect 12212 24454 12224 24506
rect 12276 24454 12288 24506
rect 12340 24454 12352 24506
rect 12404 24454 19870 24506
rect 19922 24454 19934 24506
rect 19986 24454 19998 24506
rect 20050 24454 20062 24506
rect 20114 24454 20126 24506
rect 20178 24454 27644 24506
rect 27696 24454 27708 24506
rect 27760 24454 27772 24506
rect 27824 24454 27836 24506
rect 27888 24454 27900 24506
rect 27952 24454 31648 24506
rect 552 24432 31648 24454
rect 13078 24352 13084 24404
rect 13136 24352 13142 24404
rect 13372 24364 20300 24392
rect 13372 24265 13400 24364
rect 14461 24327 14519 24333
rect 14461 24324 14473 24327
rect 13556 24296 14473 24324
rect 13556 24265 13584 24296
rect 14461 24293 14473 24296
rect 14507 24293 14519 24327
rect 14461 24287 14519 24293
rect 14642 24284 14648 24336
rect 14700 24284 14706 24336
rect 15838 24324 15844 24336
rect 15488 24296 15844 24324
rect 13357 24259 13415 24265
rect 13357 24225 13369 24259
rect 13403 24225 13415 24259
rect 13357 24219 13415 24225
rect 13449 24259 13507 24265
rect 13449 24225 13461 24259
rect 13495 24225 13507 24259
rect 13449 24219 13507 24225
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 13464 24188 13492 24219
rect 13722 24216 13728 24268
rect 13780 24216 13786 24268
rect 14185 24259 14243 24265
rect 14185 24225 14197 24259
rect 14231 24256 14243 24259
rect 14274 24256 14280 24268
rect 14231 24228 14280 24256
rect 14231 24225 14243 24228
rect 14185 24219 14243 24225
rect 14274 24216 14280 24228
rect 14332 24216 14338 24268
rect 15488 24265 15516 24296
rect 15838 24284 15844 24296
rect 15896 24284 15902 24336
rect 20272 24324 20300 24364
rect 20346 24352 20352 24404
rect 20404 24352 20410 24404
rect 21634 24392 21640 24404
rect 21560 24364 21640 24392
rect 20990 24324 20996 24336
rect 20272 24296 20996 24324
rect 20990 24284 20996 24296
rect 21048 24324 21054 24336
rect 21560 24333 21588 24364
rect 21634 24352 21640 24364
rect 21692 24352 21698 24404
rect 22005 24395 22063 24401
rect 22005 24361 22017 24395
rect 22051 24392 22063 24395
rect 22278 24392 22284 24404
rect 22051 24364 22284 24392
rect 22051 24361 22063 24364
rect 22005 24355 22063 24361
rect 22278 24352 22284 24364
rect 22336 24352 22342 24404
rect 22649 24395 22707 24401
rect 22649 24361 22661 24395
rect 22695 24392 22707 24395
rect 23566 24392 23572 24404
rect 22695 24364 23572 24392
rect 22695 24361 22707 24364
rect 22649 24355 22707 24361
rect 23566 24352 23572 24364
rect 23624 24352 23630 24404
rect 24670 24352 24676 24404
rect 24728 24352 24734 24404
rect 25038 24352 25044 24404
rect 25096 24392 25102 24404
rect 25317 24395 25375 24401
rect 25317 24392 25329 24395
rect 25096 24364 25329 24392
rect 25096 24352 25102 24364
rect 25317 24361 25329 24364
rect 25363 24361 25375 24395
rect 25317 24355 25375 24361
rect 25498 24352 25504 24404
rect 25556 24352 25562 24404
rect 27522 24352 27528 24404
rect 27580 24352 27586 24404
rect 27709 24395 27767 24401
rect 27709 24361 27721 24395
rect 27755 24392 27767 24395
rect 28258 24392 28264 24404
rect 27755 24364 28264 24392
rect 27755 24361 27767 24364
rect 27709 24355 27767 24361
rect 28258 24352 28264 24364
rect 28316 24392 28322 24404
rect 28534 24392 28540 24404
rect 28316 24364 28540 24392
rect 28316 24352 28322 24364
rect 28534 24352 28540 24364
rect 28592 24352 28598 24404
rect 21545 24327 21603 24333
rect 21048 24296 21404 24324
rect 21048 24284 21054 24296
rect 14369 24259 14427 24265
rect 14369 24225 14381 24259
rect 14415 24256 14427 24259
rect 14829 24259 14887 24265
rect 14829 24256 14841 24259
rect 14415 24228 14841 24256
rect 14415 24225 14427 24228
rect 14369 24219 14427 24225
rect 14829 24225 14841 24228
rect 14875 24256 14887 24259
rect 15381 24259 15439 24265
rect 14875 24228 15056 24256
rect 14875 24225 14887 24228
rect 14829 24219 14887 24225
rect 13906 24188 13912 24200
rect 13464 24160 13912 24188
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 12986 24080 12992 24132
rect 13044 24120 13050 24132
rect 14384 24120 14412 24219
rect 13044 24092 14412 24120
rect 15028 24120 15056 24228
rect 15381 24225 15393 24259
rect 15427 24225 15439 24259
rect 15381 24219 15439 24225
rect 15473 24259 15531 24265
rect 15473 24225 15485 24259
rect 15519 24225 15531 24259
rect 15473 24219 15531 24225
rect 15396 24188 15424 24219
rect 15562 24216 15568 24268
rect 15620 24216 15626 24268
rect 15749 24259 15807 24265
rect 15749 24225 15761 24259
rect 15795 24256 15807 24259
rect 16206 24256 16212 24268
rect 15795 24228 16212 24256
rect 15795 24225 15807 24228
rect 15749 24219 15807 24225
rect 16206 24216 16212 24228
rect 16264 24216 16270 24268
rect 16390 24216 16396 24268
rect 16448 24216 16454 24268
rect 16482 24216 16488 24268
rect 16540 24256 16546 24268
rect 16577 24259 16635 24265
rect 16577 24256 16589 24259
rect 16540 24228 16589 24256
rect 16540 24216 16546 24228
rect 16577 24225 16589 24228
rect 16623 24225 16635 24259
rect 16577 24219 16635 24225
rect 20533 24259 20591 24265
rect 20533 24225 20545 24259
rect 20579 24256 20591 24259
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 20579 24228 21281 24256
rect 20579 24225 20591 24228
rect 20533 24219 20591 24225
rect 21269 24225 21281 24228
rect 21315 24225 21327 24259
rect 21269 24219 21327 24225
rect 18966 24188 18972 24200
rect 15396 24160 18972 24188
rect 18966 24148 18972 24160
rect 19024 24148 19030 24200
rect 20717 24191 20775 24197
rect 20717 24157 20729 24191
rect 20763 24157 20775 24191
rect 21376 24188 21404 24296
rect 21545 24293 21557 24327
rect 21591 24293 21603 24327
rect 21545 24287 21603 24293
rect 21726 24284 21732 24336
rect 21784 24333 21790 24336
rect 21784 24327 21813 24333
rect 21801 24293 21813 24327
rect 22370 24324 22376 24336
rect 21784 24287 21813 24293
rect 22204 24296 22376 24324
rect 21784 24284 21790 24287
rect 21450 24216 21456 24268
rect 21508 24216 21514 24268
rect 21634 24216 21640 24268
rect 21692 24216 21698 24268
rect 22204 24265 22232 24296
rect 22370 24284 22376 24296
rect 22428 24284 22434 24336
rect 23474 24284 23480 24336
rect 23532 24324 23538 24336
rect 25516 24324 25544 24352
rect 25685 24327 25743 24333
rect 25685 24324 25697 24327
rect 23532 24296 24072 24324
rect 25516 24296 25697 24324
rect 23532 24284 23538 24296
rect 22189 24259 22247 24265
rect 22189 24225 22201 24259
rect 22235 24225 22247 24259
rect 22189 24219 22247 24225
rect 23750 24216 23756 24268
rect 23808 24265 23814 24268
rect 24044 24265 24072 24296
rect 25685 24293 25697 24296
rect 25731 24293 25743 24327
rect 25685 24287 25743 24293
rect 26142 24284 26148 24336
rect 26200 24324 26206 24336
rect 26513 24327 26571 24333
rect 26513 24324 26525 24327
rect 26200 24296 26525 24324
rect 26200 24284 26206 24296
rect 26513 24293 26525 24296
rect 26559 24293 26571 24327
rect 26513 24287 26571 24293
rect 27338 24284 27344 24336
rect 27396 24284 27402 24336
rect 27614 24284 27620 24336
rect 27672 24324 27678 24336
rect 28442 24324 28448 24336
rect 27672 24296 28448 24324
rect 27672 24284 27678 24296
rect 28442 24284 28448 24296
rect 28500 24284 28506 24336
rect 23808 24256 23820 24265
rect 24029 24259 24087 24265
rect 23808 24228 23853 24256
rect 23808 24219 23820 24228
rect 24029 24225 24041 24259
rect 24075 24225 24087 24259
rect 24029 24219 24087 24225
rect 23808 24216 23814 24219
rect 24302 24216 24308 24268
rect 24360 24216 24366 24268
rect 24949 24259 25007 24265
rect 24949 24225 24961 24259
rect 24995 24256 25007 24259
rect 24995 24228 25360 24256
rect 24995 24225 25007 24228
rect 24949 24219 25007 24225
rect 21726 24188 21732 24200
rect 21376 24160 21732 24188
rect 20717 24151 20775 24157
rect 15194 24120 15200 24132
rect 15028 24092 15200 24120
rect 13044 24080 13050 24092
rect 15194 24080 15200 24092
rect 15252 24120 15258 24132
rect 16482 24120 16488 24132
rect 15252 24092 16488 24120
rect 15252 24080 15258 24092
rect 16482 24080 16488 24092
rect 16540 24080 16546 24132
rect 20732 24120 20760 24151
rect 21726 24148 21732 24160
rect 21784 24188 21790 24200
rect 21913 24191 21971 24197
rect 21913 24188 21925 24191
rect 21784 24160 21925 24188
rect 21784 24148 21790 24160
rect 21913 24157 21925 24160
rect 21959 24157 21971 24191
rect 21913 24151 21971 24157
rect 22373 24191 22431 24197
rect 22373 24157 22385 24191
rect 22419 24157 22431 24191
rect 22373 24151 22431 24157
rect 21358 24120 21364 24132
rect 20732 24092 21364 24120
rect 21358 24080 21364 24092
rect 21416 24120 21422 24132
rect 22388 24120 22416 24151
rect 24118 24148 24124 24200
rect 24176 24188 24182 24200
rect 24213 24191 24271 24197
rect 24213 24188 24225 24191
rect 24176 24160 24225 24188
rect 24176 24148 24182 24160
rect 24213 24157 24225 24160
rect 24259 24157 24271 24191
rect 24213 24151 24271 24157
rect 24854 24148 24860 24200
rect 24912 24148 24918 24200
rect 21416 24092 22416 24120
rect 25332 24120 25360 24228
rect 25406 24216 25412 24268
rect 25464 24216 25470 24268
rect 25501 24259 25559 24265
rect 25501 24225 25513 24259
rect 25547 24256 25559 24259
rect 25590 24256 25596 24268
rect 25547 24228 25596 24256
rect 25547 24225 25559 24228
rect 25501 24219 25559 24225
rect 25516 24188 25544 24219
rect 25590 24216 25596 24228
rect 25648 24216 25654 24268
rect 25774 24216 25780 24268
rect 25832 24216 25838 24268
rect 25869 24259 25927 24265
rect 25869 24225 25881 24259
rect 25915 24256 25927 24259
rect 26050 24256 26056 24268
rect 25915 24228 26056 24256
rect 25915 24225 25927 24228
rect 25869 24219 25927 24225
rect 26050 24216 26056 24228
rect 26108 24216 26114 24268
rect 26237 24259 26295 24265
rect 26237 24225 26249 24259
rect 26283 24225 26295 24259
rect 26237 24219 26295 24225
rect 26145 24191 26203 24197
rect 26145 24188 26157 24191
rect 25516 24160 26157 24188
rect 26145 24157 26157 24160
rect 26191 24157 26203 24191
rect 26252 24188 26280 24219
rect 26418 24216 26424 24268
rect 26476 24256 26482 24268
rect 26602 24256 26608 24268
rect 26476 24228 26608 24256
rect 26476 24216 26482 24228
rect 26602 24216 26608 24228
rect 26660 24216 26666 24268
rect 27356 24256 27384 24284
rect 27522 24256 27528 24268
rect 27356 24228 27528 24256
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 28169 24259 28227 24265
rect 28169 24256 28181 24259
rect 28092 24228 28181 24256
rect 27338 24188 27344 24200
rect 26252 24160 27344 24188
rect 26145 24151 26203 24157
rect 27338 24148 27344 24160
rect 27396 24148 27402 24200
rect 28092 24132 28120 24228
rect 28169 24225 28181 24228
rect 28215 24225 28227 24259
rect 28169 24219 28227 24225
rect 28350 24216 28356 24268
rect 28408 24256 28414 24268
rect 28718 24256 28724 24268
rect 28408 24228 28724 24256
rect 28408 24216 28414 24228
rect 28718 24216 28724 24228
rect 28776 24216 28782 24268
rect 26234 24120 26240 24132
rect 25332 24092 26240 24120
rect 21416 24080 21422 24092
rect 13998 24012 14004 24064
rect 14056 24012 14062 24064
rect 15010 24012 15016 24064
rect 15068 24052 15074 24064
rect 15105 24055 15163 24061
rect 15105 24052 15117 24055
rect 15068 24024 15117 24052
rect 15068 24012 15074 24024
rect 15105 24021 15117 24024
rect 15151 24021 15163 24055
rect 15105 24015 15163 24021
rect 16209 24055 16267 24061
rect 16209 24021 16221 24055
rect 16255 24052 16267 24055
rect 16298 24052 16304 24064
rect 16255 24024 16304 24052
rect 16255 24021 16267 24024
rect 16209 24015 16267 24021
rect 16298 24012 16304 24024
rect 16356 24012 16362 24064
rect 22388 24052 22416 24092
rect 26234 24080 26240 24092
rect 26292 24080 26298 24132
rect 28074 24080 28080 24132
rect 28132 24080 28138 24132
rect 23658 24052 23664 24064
rect 22388 24024 23664 24052
rect 23658 24012 23664 24024
rect 23716 24012 23722 24064
rect 25409 24055 25467 24061
rect 25409 24021 25421 24055
rect 25455 24052 25467 24055
rect 27062 24052 27068 24064
rect 25455 24024 27068 24052
rect 25455 24021 25467 24024
rect 25409 24015 25467 24021
rect 27062 24012 27068 24024
rect 27120 24012 27126 24064
rect 27709 24055 27767 24061
rect 27709 24021 27721 24055
rect 27755 24052 27767 24055
rect 28166 24052 28172 24064
rect 27755 24024 28172 24052
rect 27755 24021 27767 24024
rect 27709 24015 27767 24021
rect 28166 24012 28172 24024
rect 28224 24012 28230 24064
rect 28350 24012 28356 24064
rect 28408 24052 28414 24064
rect 28537 24055 28595 24061
rect 28537 24052 28549 24055
rect 28408 24024 28549 24052
rect 28408 24012 28414 24024
rect 28537 24021 28549 24024
rect 28583 24021 28595 24055
rect 28537 24015 28595 24021
rect 552 23962 31648 23984
rect 552 23910 3662 23962
rect 3714 23910 3726 23962
rect 3778 23910 3790 23962
rect 3842 23910 3854 23962
rect 3906 23910 3918 23962
rect 3970 23910 11436 23962
rect 11488 23910 11500 23962
rect 11552 23910 11564 23962
rect 11616 23910 11628 23962
rect 11680 23910 11692 23962
rect 11744 23910 19210 23962
rect 19262 23910 19274 23962
rect 19326 23910 19338 23962
rect 19390 23910 19402 23962
rect 19454 23910 19466 23962
rect 19518 23910 26984 23962
rect 27036 23910 27048 23962
rect 27100 23910 27112 23962
rect 27164 23910 27176 23962
rect 27228 23910 27240 23962
rect 27292 23910 31648 23962
rect 552 23888 31648 23910
rect 16390 23808 16396 23860
rect 16448 23808 16454 23860
rect 19702 23848 19708 23860
rect 16500 23820 19708 23848
rect 13630 23740 13636 23792
rect 13688 23780 13694 23792
rect 13688 23752 14320 23780
rect 13688 23740 13694 23752
rect 13357 23715 13415 23721
rect 13357 23681 13369 23715
rect 13403 23712 13415 23715
rect 14182 23712 14188 23724
rect 13403 23684 14188 23712
rect 13403 23681 13415 23684
rect 13357 23675 13415 23681
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 14292 23721 14320 23752
rect 15396 23752 15884 23780
rect 14277 23715 14335 23721
rect 14277 23681 14289 23715
rect 14323 23681 14335 23715
rect 14277 23675 14335 23681
rect 11330 23604 11336 23656
rect 11388 23644 11394 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 11388 23616 12541 23644
rect 11388 23604 11394 23616
rect 12529 23613 12541 23616
rect 12575 23644 12587 23647
rect 14366 23644 14372 23656
rect 12575 23616 14372 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 14366 23604 14372 23616
rect 14424 23644 14430 23656
rect 15396 23653 15424 23752
rect 15856 23712 15884 23752
rect 16114 23740 16120 23792
rect 16172 23780 16178 23792
rect 16500 23780 16528 23820
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 20346 23808 20352 23860
rect 20404 23848 20410 23860
rect 20806 23848 20812 23860
rect 20404 23820 20812 23848
rect 20404 23808 20410 23820
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 25958 23808 25964 23860
rect 26016 23848 26022 23860
rect 26973 23851 27031 23857
rect 26973 23848 26985 23851
rect 26016 23820 26985 23848
rect 26016 23808 26022 23820
rect 26973 23817 26985 23820
rect 27019 23817 27031 23851
rect 26973 23811 27031 23817
rect 27893 23851 27951 23857
rect 27893 23817 27905 23851
rect 27939 23848 27951 23851
rect 28074 23848 28080 23860
rect 27939 23820 28080 23848
rect 27939 23817 27951 23820
rect 27893 23811 27951 23817
rect 28074 23808 28080 23820
rect 28132 23808 28138 23860
rect 28350 23808 28356 23860
rect 28408 23808 28414 23860
rect 28718 23808 28724 23860
rect 28776 23848 28782 23860
rect 30377 23851 30435 23857
rect 30377 23848 30389 23851
rect 28776 23820 30389 23848
rect 28776 23808 28782 23820
rect 30377 23817 30389 23820
rect 30423 23817 30435 23851
rect 30377 23811 30435 23817
rect 16172 23752 16528 23780
rect 16172 23740 16178 23752
rect 17034 23740 17040 23792
rect 17092 23780 17098 23792
rect 28442 23780 28448 23792
rect 17092 23752 20300 23780
rect 17092 23740 17098 23752
rect 17862 23712 17868 23724
rect 15856 23684 17868 23712
rect 17862 23672 17868 23684
rect 17920 23672 17926 23724
rect 19076 23684 19380 23712
rect 19076 23656 19104 23684
rect 15381 23647 15439 23653
rect 14424 23616 14688 23644
rect 14424 23604 14430 23616
rect 14660 23588 14688 23616
rect 15381 23613 15393 23647
rect 15427 23613 15439 23647
rect 15749 23647 15807 23653
rect 15749 23644 15761 23647
rect 15381 23607 15439 23613
rect 15672 23616 15761 23644
rect 12986 23536 12992 23588
rect 13044 23536 13050 23588
rect 13173 23579 13231 23585
rect 13173 23545 13185 23579
rect 13219 23576 13231 23579
rect 13219 23548 13492 23576
rect 13219 23545 13231 23548
rect 13173 23539 13231 23545
rect 12434 23468 12440 23520
rect 12492 23468 12498 23520
rect 13464 23508 13492 23548
rect 14642 23536 14648 23588
rect 14700 23536 14706 23588
rect 13725 23511 13783 23517
rect 13725 23508 13737 23511
rect 13464 23480 13737 23508
rect 13725 23477 13737 23480
rect 13771 23477 13783 23511
rect 13725 23471 13783 23477
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15252 23480 15485 23508
rect 15252 23468 15258 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15672 23508 15700 23616
rect 15749 23613 15761 23616
rect 15795 23613 15807 23647
rect 15749 23607 15807 23613
rect 15838 23604 15844 23656
rect 15896 23604 15902 23656
rect 15930 23604 15936 23656
rect 15988 23604 15994 23656
rect 16114 23604 16120 23656
rect 16172 23604 16178 23656
rect 16206 23604 16212 23656
rect 16264 23644 16270 23656
rect 16945 23647 17003 23653
rect 16945 23644 16957 23647
rect 16264 23616 16957 23644
rect 16264 23604 16270 23616
rect 16945 23613 16957 23616
rect 16991 23613 17003 23647
rect 16945 23607 17003 23613
rect 17126 23604 17132 23656
rect 17184 23604 17190 23656
rect 18782 23604 18788 23656
rect 18840 23644 18846 23656
rect 18937 23647 18995 23653
rect 18937 23644 18949 23647
rect 18840 23616 18949 23644
rect 18840 23604 18846 23616
rect 18937 23613 18949 23616
rect 18983 23613 18995 23647
rect 18937 23607 18995 23613
rect 19058 23604 19064 23656
rect 19116 23604 19122 23656
rect 19352 23653 19380 23684
rect 20272 23653 20300 23752
rect 27080 23752 28448 23780
rect 19153 23647 19211 23653
rect 19153 23613 19165 23647
rect 19199 23613 19211 23647
rect 19153 23607 19211 23613
rect 19337 23647 19395 23653
rect 19337 23613 19349 23647
rect 19383 23613 19395 23647
rect 19337 23607 19395 23613
rect 20257 23647 20315 23653
rect 20257 23613 20269 23647
rect 20303 23644 20315 23647
rect 24578 23644 24584 23656
rect 20303 23616 24584 23644
rect 20303 23613 20315 23616
rect 20257 23607 20315 23613
rect 15856 23576 15884 23604
rect 16482 23576 16488 23588
rect 15856 23548 16488 23576
rect 16482 23536 16488 23548
rect 16540 23576 16546 23588
rect 17681 23579 17739 23585
rect 17681 23576 17693 23579
rect 16540 23548 17693 23576
rect 16540 23536 16546 23548
rect 17681 23545 17693 23548
rect 17727 23545 17739 23579
rect 17681 23539 17739 23545
rect 17865 23579 17923 23585
rect 17865 23545 17877 23579
rect 17911 23576 17923 23579
rect 17954 23576 17960 23588
rect 17911 23548 17960 23576
rect 17911 23545 17923 23548
rect 17865 23539 17923 23545
rect 17954 23536 17960 23548
rect 18012 23536 18018 23588
rect 18049 23579 18107 23585
rect 18049 23545 18061 23579
rect 18095 23576 18107 23579
rect 18138 23576 18144 23588
rect 18095 23548 18144 23576
rect 18095 23545 18107 23548
rect 18049 23539 18107 23545
rect 18138 23536 18144 23548
rect 18196 23576 18202 23588
rect 19168 23576 19196 23607
rect 24578 23604 24584 23616
rect 24636 23604 24642 23656
rect 27080 23653 27108 23752
rect 28442 23740 28448 23752
rect 28500 23740 28506 23792
rect 27525 23715 27583 23721
rect 27525 23681 27537 23715
rect 27571 23712 27583 23715
rect 27614 23712 27620 23724
rect 27571 23684 27620 23712
rect 27571 23681 27583 23684
rect 27525 23675 27583 23681
rect 27614 23672 27620 23684
rect 27672 23712 27678 23724
rect 27985 23715 28043 23721
rect 27672 23684 27936 23712
rect 27672 23672 27678 23684
rect 27065 23647 27123 23653
rect 27065 23613 27077 23647
rect 27111 23613 27123 23647
rect 27065 23607 27123 23613
rect 27709 23647 27767 23653
rect 27709 23613 27721 23647
rect 27755 23613 27767 23647
rect 27908 23644 27936 23684
rect 27985 23681 27997 23715
rect 28031 23712 28043 23715
rect 28258 23712 28264 23724
rect 28031 23684 28264 23712
rect 28031 23681 28043 23684
rect 27985 23675 28043 23681
rect 28258 23672 28264 23684
rect 28316 23672 28322 23724
rect 28166 23644 28172 23656
rect 27908 23616 28172 23644
rect 27709 23607 27767 23613
rect 19242 23576 19248 23588
rect 18196 23548 18920 23576
rect 19168 23548 19248 23576
rect 18196 23536 18202 23548
rect 17034 23508 17040 23520
rect 15672 23480 17040 23508
rect 15473 23471 15531 23477
rect 17034 23468 17040 23480
rect 17092 23468 17098 23520
rect 17221 23511 17279 23517
rect 17221 23477 17233 23511
rect 17267 23508 17279 23511
rect 17586 23508 17592 23520
rect 17267 23480 17592 23508
rect 17267 23477 17279 23480
rect 17221 23471 17279 23477
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 18693 23511 18751 23517
rect 18693 23477 18705 23511
rect 18739 23508 18751 23511
rect 18782 23508 18788 23520
rect 18739 23480 18788 23508
rect 18739 23477 18751 23480
rect 18693 23471 18751 23477
rect 18782 23468 18788 23480
rect 18840 23468 18846 23520
rect 18892 23508 18920 23548
rect 19242 23536 19248 23548
rect 19300 23576 19306 23588
rect 19794 23576 19800 23588
rect 19300 23548 19800 23576
rect 19300 23536 19306 23548
rect 19794 23536 19800 23548
rect 19852 23536 19858 23588
rect 27724 23576 27752 23607
rect 28166 23604 28172 23616
rect 28224 23604 28230 23656
rect 28626 23604 28632 23656
rect 28684 23604 28690 23656
rect 28721 23647 28779 23653
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 28997 23647 29055 23653
rect 28997 23644 29009 23647
rect 28767 23616 29009 23644
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 28997 23613 29009 23616
rect 29043 23613 29055 23647
rect 28997 23607 29055 23613
rect 29242 23579 29300 23585
rect 29242 23576 29254 23579
rect 27724 23548 28120 23576
rect 28092 23520 28120 23548
rect 28552 23548 29254 23576
rect 19150 23508 19156 23520
rect 18892 23480 19156 23508
rect 19150 23468 19156 23480
rect 19208 23468 19214 23520
rect 28074 23468 28080 23520
rect 28132 23468 28138 23520
rect 28350 23468 28356 23520
rect 28408 23468 28414 23520
rect 28552 23517 28580 23548
rect 29242 23545 29254 23548
rect 29288 23545 29300 23579
rect 29242 23539 29300 23545
rect 28537 23511 28595 23517
rect 28537 23477 28549 23511
rect 28583 23477 28595 23511
rect 28537 23471 28595 23477
rect 552 23418 31648 23440
rect 552 23366 4322 23418
rect 4374 23366 4386 23418
rect 4438 23366 4450 23418
rect 4502 23366 4514 23418
rect 4566 23366 4578 23418
rect 4630 23366 12096 23418
rect 12148 23366 12160 23418
rect 12212 23366 12224 23418
rect 12276 23366 12288 23418
rect 12340 23366 12352 23418
rect 12404 23366 19870 23418
rect 19922 23366 19934 23418
rect 19986 23366 19998 23418
rect 20050 23366 20062 23418
rect 20114 23366 20126 23418
rect 20178 23366 27644 23418
rect 27696 23366 27708 23418
rect 27760 23366 27772 23418
rect 27824 23366 27836 23418
rect 27888 23366 27900 23418
rect 27952 23366 31648 23418
rect 552 23344 31648 23366
rect 12618 23264 12624 23316
rect 12676 23304 12682 23316
rect 13630 23304 13636 23316
rect 12676 23276 13636 23304
rect 12676 23264 12682 23276
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 14366 23304 14372 23316
rect 14200 23276 14372 23304
rect 12520 23239 12578 23245
rect 12520 23205 12532 23239
rect 12566 23236 12578 23239
rect 13725 23239 13783 23245
rect 13725 23236 13737 23239
rect 12566 23208 13737 23236
rect 12566 23205 12578 23208
rect 12520 23199 12578 23205
rect 13725 23205 13737 23208
rect 13771 23205 13783 23239
rect 13725 23199 13783 23205
rect 13906 23196 13912 23248
rect 13964 23236 13970 23248
rect 14200 23236 14228 23276
rect 14366 23264 14372 23276
rect 14424 23304 14430 23316
rect 14424 23276 15424 23304
rect 14424 23264 14430 23276
rect 15286 23236 15292 23248
rect 13964 23208 14228 23236
rect 14384 23208 15292 23236
rect 13964 23196 13970 23208
rect 12253 23171 12311 23177
rect 12253 23137 12265 23171
rect 12299 23168 12311 23171
rect 12342 23168 12348 23180
rect 12299 23140 12348 23168
rect 12299 23137 12311 23140
rect 12253 23131 12311 23137
rect 12342 23128 12348 23140
rect 12400 23128 12406 23180
rect 14108 23177 14136 23208
rect 14001 23171 14059 23177
rect 14001 23137 14013 23171
rect 14047 23137 14059 23171
rect 14001 23131 14059 23137
rect 14093 23171 14151 23177
rect 14093 23137 14105 23171
rect 14139 23137 14151 23171
rect 14093 23131 14151 23137
rect 14016 23100 14044 23131
rect 14182 23128 14188 23180
rect 14240 23128 14246 23180
rect 14384 23177 14412 23208
rect 15286 23196 15292 23208
rect 15344 23196 15350 23248
rect 15396 23236 15424 23276
rect 15746 23264 15752 23316
rect 15804 23304 15810 23316
rect 16206 23304 16212 23316
rect 15804 23276 16212 23304
rect 15804 23264 15810 23276
rect 16206 23264 16212 23276
rect 16264 23264 16270 23316
rect 17862 23264 17868 23316
rect 17920 23304 17926 23316
rect 22186 23304 22192 23316
rect 17920 23276 22192 23304
rect 17920 23264 17926 23276
rect 22186 23264 22192 23276
rect 22244 23304 22250 23316
rect 23382 23304 23388 23316
rect 22244 23276 23388 23304
rect 22244 23264 22250 23276
rect 16482 23236 16488 23248
rect 15396 23208 16488 23236
rect 16482 23196 16488 23208
rect 16540 23196 16546 23248
rect 17126 23196 17132 23248
rect 17184 23236 17190 23248
rect 17678 23236 17684 23248
rect 17184 23208 17684 23236
rect 17184 23196 17190 23208
rect 17678 23196 17684 23208
rect 17736 23236 17742 23248
rect 22002 23236 22008 23248
rect 17736 23208 19564 23236
rect 17736 23196 17742 23208
rect 14369 23171 14427 23177
rect 14369 23137 14381 23171
rect 14415 23137 14427 23171
rect 14369 23131 14427 23137
rect 14642 23128 14648 23180
rect 14700 23128 14706 23180
rect 16850 23128 16856 23180
rect 16908 23168 16914 23180
rect 17322 23171 17380 23177
rect 17322 23168 17334 23171
rect 16908 23140 17334 23168
rect 16908 23128 16914 23140
rect 17322 23137 17334 23140
rect 17368 23137 17380 23171
rect 17322 23131 17380 23137
rect 17586 23128 17592 23180
rect 17644 23128 17650 23180
rect 17880 23177 17908 23208
rect 17865 23171 17923 23177
rect 17865 23137 17877 23171
rect 17911 23137 17923 23171
rect 17865 23131 17923 23137
rect 18690 23128 18696 23180
rect 18748 23168 18754 23180
rect 18874 23168 18880 23180
rect 18748 23140 18880 23168
rect 18748 23128 18754 23140
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 19150 23128 19156 23180
rect 19208 23128 19214 23180
rect 19536 23177 19564 23208
rect 19996 23208 22008 23236
rect 19521 23171 19579 23177
rect 19521 23137 19533 23171
rect 19567 23168 19579 23171
rect 19613 23171 19671 23177
rect 19613 23168 19625 23171
rect 19567 23140 19625 23168
rect 19567 23137 19579 23140
rect 19521 23131 19579 23137
rect 19613 23137 19625 23140
rect 19659 23137 19671 23171
rect 19613 23131 19671 23137
rect 19702 23128 19708 23180
rect 19760 23168 19766 23180
rect 19889 23171 19947 23177
rect 19889 23168 19901 23171
rect 19760 23140 19901 23168
rect 19760 23128 19766 23140
rect 19889 23137 19901 23140
rect 19935 23137 19947 23171
rect 19889 23131 19947 23137
rect 14826 23100 14832 23112
rect 14016 23072 14832 23100
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23100 19303 23103
rect 19996 23100 20024 23208
rect 20732 23180 20760 23208
rect 22002 23196 22008 23208
rect 22060 23196 22066 23248
rect 22296 23245 22324 23276
rect 23382 23264 23388 23276
rect 23440 23304 23446 23316
rect 23440 23276 25084 23304
rect 23440 23264 23446 23276
rect 22281 23239 22339 23245
rect 22281 23205 22293 23239
rect 22327 23205 22339 23239
rect 22281 23199 22339 23205
rect 23106 23196 23112 23248
rect 23164 23236 23170 23248
rect 25056 23245 25084 23276
rect 26786 23264 26792 23316
rect 26844 23304 26850 23316
rect 27430 23304 27436 23316
rect 26844 23276 27436 23304
rect 26844 23264 26850 23276
rect 27430 23264 27436 23276
rect 27488 23304 27494 23316
rect 27525 23307 27583 23313
rect 27525 23304 27537 23307
rect 27488 23276 27537 23304
rect 27488 23264 27494 23276
rect 27525 23273 27537 23276
rect 27571 23273 27583 23307
rect 28718 23304 28724 23316
rect 27525 23267 27583 23273
rect 28368 23276 28724 23304
rect 25041 23239 25099 23245
rect 23164 23208 23520 23236
rect 23164 23196 23170 23208
rect 20073 23171 20131 23177
rect 20073 23137 20085 23171
rect 20119 23137 20131 23171
rect 20073 23131 20131 23137
rect 19291 23072 20024 23100
rect 20088 23100 20116 23131
rect 20714 23128 20720 23180
rect 20772 23128 20778 23180
rect 20990 23128 20996 23180
rect 21048 23128 21054 23180
rect 21266 23128 21272 23180
rect 21324 23128 21330 23180
rect 21358 23128 21364 23180
rect 21416 23168 21422 23180
rect 21729 23171 21787 23177
rect 21729 23168 21741 23171
rect 21416 23140 21741 23168
rect 21416 23128 21422 23140
rect 21729 23137 21741 23140
rect 21775 23137 21787 23171
rect 21729 23131 21787 23137
rect 21913 23171 21971 23177
rect 21913 23137 21925 23171
rect 21959 23137 21971 23171
rect 21913 23131 21971 23137
rect 21450 23100 21456 23112
rect 20088 23072 21456 23100
rect 19291 23069 19303 23072
rect 19245 23063 19303 23069
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 21634 23060 21640 23112
rect 21692 23100 21698 23112
rect 21928 23100 21956 23131
rect 22094 23128 22100 23180
rect 22152 23168 22158 23180
rect 22554 23168 22560 23180
rect 22152 23140 22560 23168
rect 22152 23128 22158 23140
rect 22554 23128 22560 23140
rect 22612 23128 22618 23180
rect 23492 23177 23520 23208
rect 25041 23205 25053 23239
rect 25087 23205 25099 23239
rect 25041 23199 25099 23205
rect 25406 23196 25412 23248
rect 25464 23236 25470 23248
rect 27982 23236 27988 23248
rect 25464 23208 27016 23236
rect 25464 23196 25470 23208
rect 23477 23171 23535 23177
rect 23477 23137 23489 23171
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 24026 23128 24032 23180
rect 24084 23128 24090 23180
rect 24121 23171 24179 23177
rect 24121 23137 24133 23171
rect 24167 23137 24179 23171
rect 24121 23131 24179 23137
rect 21692 23072 21956 23100
rect 22572 23100 22600 23128
rect 24136 23100 24164 23131
rect 24210 23128 24216 23180
rect 24268 23128 24274 23180
rect 24351 23171 24409 23177
rect 24351 23137 24363 23171
rect 24397 23168 24409 23171
rect 24670 23168 24676 23180
rect 24397 23140 24676 23168
rect 24397 23137 24409 23140
rect 24351 23131 24409 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 26988 23177 27016 23208
rect 27632 23208 27988 23236
rect 27632 23180 27660 23208
rect 27982 23196 27988 23208
rect 28040 23196 28046 23248
rect 28074 23196 28080 23248
rect 28132 23245 28138 23248
rect 28368 23245 28396 23276
rect 28718 23264 28724 23276
rect 28776 23264 28782 23316
rect 28132 23239 28195 23245
rect 28132 23205 28149 23239
rect 28183 23205 28195 23239
rect 28132 23199 28195 23205
rect 28353 23239 28411 23245
rect 28353 23205 28365 23239
rect 28399 23205 28411 23239
rect 28353 23199 28411 23205
rect 28132 23196 28138 23199
rect 28534 23196 28540 23248
rect 28592 23196 28598 23248
rect 28736 23236 28764 23264
rect 28736 23208 29040 23236
rect 26605 23171 26663 23177
rect 26605 23137 26617 23171
rect 26651 23137 26663 23171
rect 26605 23131 26663 23137
rect 26973 23171 27031 23177
rect 26973 23137 26985 23171
rect 27019 23137 27031 23171
rect 26973 23131 27031 23137
rect 22572 23072 24164 23100
rect 21692 23060 21698 23072
rect 24486 23060 24492 23112
rect 24544 23060 24550 23112
rect 25869 23103 25927 23109
rect 25869 23069 25881 23103
rect 25915 23100 25927 23103
rect 26326 23100 26332 23112
rect 25915 23072 26332 23100
rect 25915 23069 25927 23072
rect 25869 23063 25927 23069
rect 26326 23060 26332 23072
rect 26384 23060 26390 23112
rect 26620 23100 26648 23131
rect 27614 23128 27620 23180
rect 27672 23128 27678 23180
rect 27709 23171 27767 23177
rect 27709 23137 27721 23171
rect 27755 23168 27767 23171
rect 28902 23168 28908 23180
rect 27755 23140 28908 23168
rect 27755 23137 27767 23140
rect 27709 23131 27767 23137
rect 28902 23128 28908 23140
rect 28960 23128 28966 23180
rect 27341 23103 27399 23109
rect 27341 23100 27353 23103
rect 26620 23072 27353 23100
rect 27341 23069 27353 23072
rect 27387 23100 27399 23103
rect 28810 23100 28816 23112
rect 27387 23072 28816 23100
rect 27387 23069 27399 23072
rect 27341 23063 27399 23069
rect 28810 23060 28816 23072
rect 28868 23060 28874 23112
rect 29012 23100 29040 23208
rect 28920 23072 29040 23100
rect 19610 23032 19616 23044
rect 17604 23004 19616 23032
rect 16574 22924 16580 22976
rect 16632 22964 16638 22976
rect 17604 22964 17632 23004
rect 19610 22992 19616 23004
rect 19668 22992 19674 23044
rect 20346 22992 20352 23044
rect 20404 23032 20410 23044
rect 20717 23035 20775 23041
rect 20717 23032 20729 23035
rect 20404 23004 20729 23032
rect 20404 22992 20410 23004
rect 20717 23001 20729 23004
rect 20763 23001 20775 23035
rect 20717 22995 20775 23001
rect 22278 22992 22284 23044
rect 22336 23032 22342 23044
rect 23845 23035 23903 23041
rect 23845 23032 23857 23035
rect 22336 23004 23857 23032
rect 22336 22992 22342 23004
rect 23845 23001 23857 23004
rect 23891 23001 23903 23035
rect 23845 22995 23903 23001
rect 26878 22992 26884 23044
rect 26936 23032 26942 23044
rect 27430 23032 27436 23044
rect 26936 23004 27436 23032
rect 26936 22992 26942 23004
rect 27430 22992 27436 23004
rect 27488 22992 27494 23044
rect 27985 23035 28043 23041
rect 27985 23001 27997 23035
rect 28031 23032 28043 23035
rect 28258 23032 28264 23044
rect 28031 23004 28264 23032
rect 28031 23001 28043 23004
rect 27985 22995 28043 23001
rect 28258 22992 28264 23004
rect 28316 22992 28322 23044
rect 28350 22992 28356 23044
rect 28408 23032 28414 23044
rect 28718 23032 28724 23044
rect 28408 23004 28724 23032
rect 28408 22992 28414 23004
rect 28718 22992 28724 23004
rect 28776 22992 28782 23044
rect 16632 22936 17632 22964
rect 16632 22924 16638 22936
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 18932 22936 19441 22964
rect 18932 22924 18938 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 19429 22927 19487 22933
rect 19702 22924 19708 22976
rect 19760 22924 19766 22976
rect 19978 22924 19984 22976
rect 20036 22924 20042 22976
rect 21174 22924 21180 22976
rect 21232 22964 21238 22976
rect 21361 22967 21419 22973
rect 21361 22964 21373 22967
rect 21232 22936 21373 22964
rect 21232 22924 21238 22936
rect 21361 22933 21373 22936
rect 21407 22933 21419 22967
rect 21361 22927 21419 22933
rect 23106 22924 23112 22976
rect 23164 22964 23170 22976
rect 23385 22967 23443 22973
rect 23385 22964 23397 22967
rect 23164 22936 23397 22964
rect 23164 22924 23170 22936
rect 23385 22933 23397 22936
rect 23431 22933 23443 22967
rect 23385 22927 23443 22933
rect 25314 22924 25320 22976
rect 25372 22964 25378 22976
rect 26513 22967 26571 22973
rect 26513 22964 26525 22967
rect 25372 22936 26525 22964
rect 25372 22924 25378 22936
rect 26513 22933 26525 22936
rect 26559 22933 26571 22967
rect 26513 22927 26571 22933
rect 26602 22924 26608 22976
rect 26660 22964 26666 22976
rect 27065 22967 27123 22973
rect 27065 22964 27077 22967
rect 26660 22936 27077 22964
rect 26660 22924 26666 22936
rect 27065 22933 27077 22936
rect 27111 22933 27123 22967
rect 27065 22927 27123 22933
rect 27893 22967 27951 22973
rect 27893 22933 27905 22967
rect 27939 22964 27951 22967
rect 28074 22964 28080 22976
rect 27939 22936 28080 22964
rect 27939 22933 27951 22936
rect 27893 22927 27951 22933
rect 28074 22924 28080 22936
rect 28132 22924 28138 22976
rect 28166 22924 28172 22976
rect 28224 22924 28230 22976
rect 28810 22924 28816 22976
rect 28868 22964 28874 22976
rect 28920 22964 28948 23072
rect 28868 22936 28948 22964
rect 28868 22924 28874 22936
rect 552 22874 31648 22896
rect 552 22822 3662 22874
rect 3714 22822 3726 22874
rect 3778 22822 3790 22874
rect 3842 22822 3854 22874
rect 3906 22822 3918 22874
rect 3970 22822 11436 22874
rect 11488 22822 11500 22874
rect 11552 22822 11564 22874
rect 11616 22822 11628 22874
rect 11680 22822 11692 22874
rect 11744 22822 19210 22874
rect 19262 22822 19274 22874
rect 19326 22822 19338 22874
rect 19390 22822 19402 22874
rect 19454 22822 19466 22874
rect 19518 22822 26984 22874
rect 27036 22822 27048 22874
rect 27100 22822 27112 22874
rect 27164 22822 27176 22874
rect 27228 22822 27240 22874
rect 27292 22822 31648 22874
rect 552 22800 31648 22822
rect 16114 22760 16120 22772
rect 14200 22732 16120 22760
rect 13357 22695 13415 22701
rect 13357 22661 13369 22695
rect 13403 22692 13415 22695
rect 14090 22692 14096 22704
rect 13403 22664 14096 22692
rect 13403 22661 13415 22664
rect 13357 22655 13415 22661
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 14200 22624 14228 22732
rect 16114 22720 16120 22732
rect 16172 22720 16178 22772
rect 16850 22720 16856 22772
rect 16908 22720 16914 22772
rect 19702 22760 19708 22772
rect 19352 22732 19708 22760
rect 13832 22596 14228 22624
rect 14292 22596 14688 22624
rect 13832 22565 13860 22596
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 12667 22528 13553 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 13541 22525 13553 22528
rect 13587 22525 13599 22559
rect 13541 22519 13599 22525
rect 13817 22559 13875 22565
rect 13817 22525 13829 22559
rect 13863 22525 13875 22559
rect 13817 22519 13875 22525
rect 12986 22448 12992 22500
rect 13044 22448 13050 22500
rect 13173 22491 13231 22497
rect 13173 22457 13185 22491
rect 13219 22457 13231 22491
rect 13556 22488 13584 22519
rect 13998 22516 14004 22568
rect 14056 22516 14062 22568
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22525 14151 22559
rect 14093 22519 14151 22525
rect 14185 22559 14243 22565
rect 14185 22525 14197 22559
rect 14231 22558 14243 22559
rect 14292 22558 14320 22596
rect 14231 22530 14320 22558
rect 14231 22525 14243 22530
rect 14185 22519 14243 22525
rect 13906 22488 13912 22500
rect 13556 22460 13912 22488
rect 13173 22451 13231 22457
rect 12710 22380 12716 22432
rect 12768 22380 12774 22432
rect 12802 22380 12808 22432
rect 12860 22420 12866 22432
rect 13188 22420 13216 22451
rect 13906 22448 13912 22460
rect 13964 22448 13970 22500
rect 14108 22488 14136 22519
rect 14550 22516 14556 22568
rect 14608 22516 14614 22568
rect 14660 22556 14688 22596
rect 17678 22584 17684 22636
rect 17736 22624 17742 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 17736 22596 17877 22624
rect 17736 22584 17742 22596
rect 17865 22593 17877 22596
rect 17911 22593 17923 22627
rect 17865 22587 17923 22593
rect 17954 22584 17960 22636
rect 18012 22624 18018 22636
rect 19352 22633 19380 22732
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 20717 22763 20775 22769
rect 20717 22729 20729 22763
rect 20763 22760 20775 22763
rect 21266 22760 21272 22772
rect 20763 22732 21272 22760
rect 20763 22729 20775 22732
rect 20717 22723 20775 22729
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 21450 22720 21456 22772
rect 21508 22720 21514 22772
rect 21818 22760 21824 22772
rect 21551 22732 21824 22760
rect 20990 22652 20996 22704
rect 21048 22692 21054 22704
rect 21551 22692 21579 22732
rect 21818 22720 21824 22732
rect 21876 22760 21882 22772
rect 21876 22732 24624 22760
rect 21876 22720 21882 22732
rect 22094 22692 22100 22704
rect 21048 22664 21579 22692
rect 21836 22664 22100 22692
rect 21048 22652 21054 22664
rect 19337 22627 19395 22633
rect 18012 22596 18368 22624
rect 18012 22584 18018 22596
rect 14820 22559 14878 22565
rect 14660 22528 14780 22556
rect 14366 22488 14372 22500
rect 14108 22460 14372 22488
rect 14366 22448 14372 22460
rect 14424 22448 14430 22500
rect 14752 22488 14780 22528
rect 14820 22525 14832 22559
rect 14866 22556 14878 22559
rect 15194 22556 15200 22568
rect 14866 22528 15200 22556
rect 14866 22525 14878 22528
rect 14820 22519 14878 22525
rect 15194 22516 15200 22528
rect 15252 22516 15258 22568
rect 15286 22516 15292 22568
rect 15344 22556 15350 22568
rect 16209 22559 16267 22565
rect 16209 22556 16221 22559
rect 15344 22528 16221 22556
rect 15344 22516 15350 22528
rect 16209 22525 16221 22528
rect 16255 22525 16267 22559
rect 16209 22519 16267 22525
rect 16298 22516 16304 22568
rect 16356 22556 16362 22568
rect 16393 22559 16451 22565
rect 16393 22556 16405 22559
rect 16356 22528 16405 22556
rect 16356 22516 16362 22528
rect 16393 22525 16405 22528
rect 16439 22525 16451 22559
rect 16393 22519 16451 22525
rect 16482 22516 16488 22568
rect 16540 22516 16546 22568
rect 16574 22516 16580 22568
rect 16632 22516 16638 22568
rect 17129 22559 17187 22565
rect 17129 22525 17141 22559
rect 17175 22556 17187 22559
rect 17770 22556 17776 22568
rect 17175 22528 17776 22556
rect 17175 22525 17187 22528
rect 17129 22519 17187 22525
rect 17770 22516 17776 22528
rect 17828 22516 17834 22568
rect 18138 22516 18144 22568
rect 18196 22516 18202 22568
rect 18340 22565 18368 22596
rect 19337 22593 19349 22627
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 20346 22584 20352 22636
rect 20404 22624 20410 22636
rect 20404 22596 21312 22624
rect 20404 22584 20410 22596
rect 18325 22559 18383 22565
rect 18325 22525 18337 22559
rect 18371 22556 18383 22559
rect 18414 22556 18420 22568
rect 18371 22528 18420 22556
rect 18371 22525 18383 22528
rect 18325 22519 18383 22525
rect 18414 22516 18420 22528
rect 18472 22516 18478 22568
rect 18690 22516 18696 22568
rect 18748 22516 18754 22568
rect 18782 22516 18788 22568
rect 18840 22556 18846 22568
rect 18877 22559 18935 22565
rect 18877 22556 18889 22559
rect 18840 22528 18889 22556
rect 18840 22516 18846 22528
rect 18877 22525 18889 22528
rect 18923 22525 18935 22559
rect 18877 22519 18935 22525
rect 19604 22559 19662 22565
rect 19604 22525 19616 22559
rect 19650 22556 19662 22559
rect 19978 22556 19984 22568
rect 19650 22528 19984 22556
rect 19650 22525 19662 22528
rect 19604 22519 19662 22525
rect 19978 22516 19984 22528
rect 20036 22516 20042 22568
rect 20806 22516 20812 22568
rect 20864 22516 20870 22568
rect 21082 22516 21088 22568
rect 21140 22516 21146 22568
rect 21174 22516 21180 22568
rect 21232 22516 21238 22568
rect 21284 22565 21312 22596
rect 21836 22565 21864 22664
rect 22094 22652 22100 22664
rect 22152 22652 22158 22704
rect 22186 22652 22192 22704
rect 22244 22692 22250 22704
rect 22738 22692 22744 22704
rect 22244 22664 22744 22692
rect 22244 22652 22250 22664
rect 22738 22652 22744 22664
rect 22796 22692 22802 22704
rect 24486 22692 24492 22704
rect 22796 22664 24492 22692
rect 22796 22652 22802 22664
rect 24486 22652 24492 22664
rect 24544 22652 24550 22704
rect 23845 22627 23903 22633
rect 23845 22624 23857 22627
rect 21928 22596 23857 22624
rect 21928 22565 21956 22596
rect 23845 22593 23857 22596
rect 23891 22593 23903 22627
rect 23845 22587 23903 22593
rect 21269 22559 21327 22565
rect 21269 22525 21281 22559
rect 21315 22556 21327 22559
rect 21729 22559 21787 22565
rect 21729 22556 21741 22559
rect 21315 22528 21741 22556
rect 21315 22525 21327 22528
rect 21269 22519 21327 22525
rect 21729 22525 21741 22528
rect 21775 22525 21787 22559
rect 21729 22519 21787 22525
rect 21821 22559 21879 22565
rect 21821 22525 21833 22559
rect 21867 22525 21879 22559
rect 21821 22519 21879 22525
rect 21913 22559 21971 22565
rect 21913 22525 21925 22559
rect 21959 22525 21971 22559
rect 21913 22519 21971 22525
rect 22002 22516 22008 22568
rect 22060 22565 22066 22568
rect 22060 22559 22089 22565
rect 22077 22525 22089 22559
rect 22060 22519 22089 22525
rect 22060 22516 22066 22519
rect 22186 22516 22192 22568
rect 22244 22516 22250 22568
rect 22925 22559 22983 22565
rect 22925 22525 22937 22559
rect 22971 22556 22983 22559
rect 23014 22556 23020 22568
rect 22971 22528 23020 22556
rect 22971 22525 22983 22528
rect 22925 22519 22983 22525
rect 23014 22516 23020 22528
rect 23072 22516 23078 22568
rect 23400 22528 24348 22556
rect 17402 22488 17408 22500
rect 14752 22460 17408 22488
rect 17402 22448 17408 22460
rect 17460 22448 17466 22500
rect 20714 22448 20720 22500
rect 20772 22488 20778 22500
rect 20947 22491 21005 22497
rect 20947 22488 20959 22491
rect 20772 22460 20959 22488
rect 20772 22448 20778 22460
rect 20947 22457 20959 22460
rect 20993 22457 21005 22491
rect 21192 22488 21220 22516
rect 23400 22488 23428 22528
rect 21192 22460 23428 22488
rect 23477 22491 23535 22497
rect 20947 22451 21005 22457
rect 23477 22457 23489 22491
rect 23523 22457 23535 22491
rect 24320 22488 24348 22528
rect 24394 22516 24400 22568
rect 24452 22516 24458 22568
rect 24596 22565 24624 22732
rect 27430 22652 27436 22704
rect 27488 22652 27494 22704
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 27154 22624 27160 22636
rect 26384 22596 27160 22624
rect 26384 22584 26390 22596
rect 24581 22559 24639 22565
rect 24581 22525 24593 22559
rect 24627 22525 24639 22559
rect 24581 22519 24639 22525
rect 24670 22516 24676 22568
rect 24728 22556 24734 22568
rect 24765 22559 24823 22565
rect 24765 22556 24777 22559
rect 24728 22528 24777 22556
rect 24728 22516 24734 22528
rect 24765 22525 24777 22528
rect 24811 22525 24823 22559
rect 26988 22542 27016 22596
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27448 22624 27476 22652
rect 27448 22596 27660 22624
rect 27249 22559 27307 22565
rect 27249 22556 27261 22559
rect 24765 22519 24823 22525
rect 27080 22528 27261 22556
rect 24320 22460 25084 22488
rect 23477 22451 23535 22457
rect 12860 22392 13216 22420
rect 13633 22423 13691 22429
rect 12860 22380 12866 22392
rect 13633 22389 13645 22423
rect 13679 22420 13691 22423
rect 13998 22420 14004 22432
rect 13679 22392 14004 22420
rect 13679 22389 13691 22392
rect 13633 22383 13691 22389
rect 13998 22380 14004 22392
rect 14056 22380 14062 22432
rect 14458 22380 14464 22432
rect 14516 22380 14522 22432
rect 15470 22380 15476 22432
rect 15528 22420 15534 22432
rect 15933 22423 15991 22429
rect 15933 22420 15945 22423
rect 15528 22392 15945 22420
rect 15528 22380 15534 22392
rect 15933 22389 15945 22392
rect 15979 22420 15991 22423
rect 16206 22420 16212 22432
rect 15979 22392 16212 22420
rect 15979 22389 15991 22392
rect 15933 22383 15991 22389
rect 16206 22380 16212 22392
rect 16264 22380 16270 22432
rect 16298 22380 16304 22432
rect 16356 22420 16362 22432
rect 18233 22423 18291 22429
rect 18233 22420 18245 22423
rect 16356 22392 18245 22420
rect 16356 22380 16362 22392
rect 18233 22389 18245 22392
rect 18279 22389 18291 22423
rect 18233 22383 18291 22389
rect 18969 22423 19027 22429
rect 18969 22389 18981 22423
rect 19015 22420 19027 22423
rect 20438 22420 20444 22432
rect 19015 22392 20444 22420
rect 19015 22389 19027 22392
rect 18969 22383 19027 22389
rect 20438 22380 20444 22392
rect 20496 22380 20502 22432
rect 21542 22380 21548 22432
rect 21600 22380 21606 22432
rect 23198 22380 23204 22432
rect 23256 22420 23262 22432
rect 23385 22423 23443 22429
rect 23385 22420 23397 22423
rect 23256 22392 23397 22420
rect 23256 22380 23262 22392
rect 23385 22389 23397 22392
rect 23431 22389 23443 22423
rect 23492 22420 23520 22451
rect 23658 22420 23664 22432
rect 23492 22392 23664 22420
rect 23385 22383 23443 22389
rect 23658 22380 23664 22392
rect 23716 22380 23722 22432
rect 24026 22380 24032 22432
rect 24084 22420 24090 22432
rect 24673 22423 24731 22429
rect 24673 22420 24685 22423
rect 24084 22392 24685 22420
rect 24084 22380 24090 22392
rect 24673 22389 24685 22392
rect 24719 22420 24731 22423
rect 24762 22420 24768 22432
rect 24719 22392 24768 22420
rect 24719 22389 24731 22392
rect 24673 22383 24731 22389
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 25056 22420 25084 22460
rect 25130 22448 25136 22500
rect 25188 22488 25194 22500
rect 27080 22488 27108 22528
rect 27249 22525 27261 22528
rect 27295 22525 27307 22559
rect 27249 22519 27307 22525
rect 27342 22559 27400 22565
rect 27342 22525 27354 22559
rect 27388 22525 27400 22559
rect 27342 22519 27400 22525
rect 25188 22460 27108 22488
rect 25188 22448 25194 22460
rect 27154 22448 27160 22500
rect 27212 22488 27218 22500
rect 27356 22488 27384 22519
rect 27430 22516 27436 22568
rect 27488 22565 27494 22568
rect 27632 22565 27660 22596
rect 27488 22559 27537 22565
rect 27488 22525 27491 22559
rect 27525 22558 27537 22559
rect 27614 22559 27672 22565
rect 27525 22528 27561 22558
rect 27525 22525 27537 22528
rect 27488 22519 27537 22525
rect 27614 22525 27626 22559
rect 27660 22525 27672 22559
rect 27614 22519 27672 22525
rect 27714 22559 27772 22565
rect 27714 22525 27726 22559
rect 27760 22525 27772 22559
rect 27714 22519 27772 22525
rect 27488 22516 27494 22519
rect 27729 22488 27757 22519
rect 28626 22516 28632 22568
rect 28684 22556 28690 22568
rect 28721 22559 28779 22565
rect 28721 22556 28733 22559
rect 28684 22528 28733 22556
rect 28684 22516 28690 22528
rect 28721 22525 28733 22528
rect 28767 22556 28779 22559
rect 28994 22556 29000 22568
rect 28767 22528 29000 22556
rect 28767 22525 28779 22528
rect 28721 22519 28779 22525
rect 28994 22516 29000 22528
rect 29052 22516 29058 22568
rect 27212 22460 27384 22488
rect 27693 22460 27757 22488
rect 27212 22448 27218 22460
rect 26786 22420 26792 22432
rect 25056 22392 26792 22420
rect 26786 22380 26792 22392
rect 26844 22420 26850 22432
rect 27693 22420 27721 22460
rect 26844 22392 27721 22420
rect 27893 22423 27951 22429
rect 26844 22380 26850 22392
rect 27893 22389 27905 22423
rect 27939 22420 27951 22423
rect 27982 22420 27988 22432
rect 27939 22392 27988 22420
rect 27939 22389 27951 22392
rect 27893 22383 27951 22389
rect 27982 22380 27988 22392
rect 28040 22380 28046 22432
rect 28442 22380 28448 22432
rect 28500 22420 28506 22432
rect 28629 22423 28687 22429
rect 28629 22420 28641 22423
rect 28500 22392 28641 22420
rect 28500 22380 28506 22392
rect 28629 22389 28641 22392
rect 28675 22389 28687 22423
rect 28629 22383 28687 22389
rect 552 22330 31648 22352
rect 552 22278 4322 22330
rect 4374 22278 4386 22330
rect 4438 22278 4450 22330
rect 4502 22278 4514 22330
rect 4566 22278 4578 22330
rect 4630 22278 12096 22330
rect 12148 22278 12160 22330
rect 12212 22278 12224 22330
rect 12276 22278 12288 22330
rect 12340 22278 12352 22330
rect 12404 22278 19870 22330
rect 19922 22278 19934 22330
rect 19986 22278 19998 22330
rect 20050 22278 20062 22330
rect 20114 22278 20126 22330
rect 20178 22278 27644 22330
rect 27696 22278 27708 22330
rect 27760 22278 27772 22330
rect 27824 22278 27836 22330
rect 27888 22278 27900 22330
rect 27952 22278 31648 22330
rect 552 22256 31648 22278
rect 12529 22219 12587 22225
rect 12529 22185 12541 22219
rect 12575 22216 12587 22219
rect 12802 22216 12808 22228
rect 12575 22188 12808 22216
rect 12575 22185 12587 22188
rect 12529 22179 12587 22185
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 13906 22176 13912 22228
rect 13964 22216 13970 22228
rect 14642 22216 14648 22228
rect 13964 22188 14648 22216
rect 13964 22176 13970 22188
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 18782 22216 18788 22228
rect 18616 22188 18788 22216
rect 12710 22108 12716 22160
rect 12768 22148 12774 22160
rect 14268 22151 14326 22157
rect 12768 22120 13952 22148
rect 12768 22108 12774 22120
rect 13630 22040 13636 22092
rect 13688 22089 13694 22092
rect 13924 22089 13952 22120
rect 14268 22117 14280 22151
rect 14314 22148 14326 22151
rect 14458 22148 14464 22160
rect 14314 22120 14464 22148
rect 14314 22117 14326 22120
rect 14268 22111 14326 22117
rect 14458 22108 14464 22120
rect 14516 22108 14522 22160
rect 15473 22151 15531 22157
rect 15473 22117 15485 22151
rect 15519 22148 15531 22151
rect 16298 22148 16304 22160
rect 15519 22120 16304 22148
rect 15519 22117 15531 22120
rect 15473 22111 15531 22117
rect 16298 22108 16304 22120
rect 16356 22108 16362 22160
rect 18616 22157 18644 22188
rect 18782 22176 18788 22188
rect 18840 22176 18846 22228
rect 20165 22219 20223 22225
rect 20165 22185 20177 22219
rect 20211 22185 20223 22219
rect 20165 22179 20223 22185
rect 18601 22151 18659 22157
rect 18601 22148 18613 22151
rect 17420 22120 17908 22148
rect 13688 22043 13700 22089
rect 13909 22083 13967 22089
rect 13909 22049 13921 22083
rect 13955 22049 13967 22083
rect 13909 22043 13967 22049
rect 13688 22040 13694 22043
rect 13998 22040 14004 22092
rect 14056 22040 14062 22092
rect 15657 22083 15715 22089
rect 15657 22049 15669 22083
rect 15703 22080 15715 22083
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 15703 22052 16129 22080
rect 15703 22049 15715 22052
rect 15657 22043 15715 22049
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16117 22043 16175 22049
rect 16206 22040 16212 22092
rect 16264 22080 16270 22092
rect 16669 22083 16727 22089
rect 16669 22080 16681 22083
rect 16264 22052 16681 22080
rect 16264 22040 16270 22052
rect 16669 22049 16681 22052
rect 16715 22049 16727 22083
rect 16669 22043 16727 22049
rect 17310 22040 17316 22092
rect 17368 22040 17374 22092
rect 17420 22089 17448 22120
rect 17405 22083 17463 22089
rect 17405 22049 17417 22083
rect 17451 22049 17463 22083
rect 17405 22043 17463 22049
rect 17497 22083 17555 22089
rect 17497 22049 17509 22083
rect 17543 22080 17555 22083
rect 17586 22080 17592 22092
rect 17543 22052 17592 22080
rect 17543 22049 17555 22052
rect 17497 22043 17555 22049
rect 15841 22015 15899 22021
rect 15841 21981 15853 22015
rect 15887 22012 15899 22015
rect 15930 22012 15936 22024
rect 15887 21984 15936 22012
rect 15887 21981 15899 21984
rect 15841 21975 15899 21981
rect 15930 21972 15936 21984
rect 15988 21972 15994 22024
rect 17420 22012 17448 22043
rect 17586 22040 17592 22052
rect 17644 22040 17650 22092
rect 17681 22083 17739 22089
rect 17681 22049 17693 22083
rect 17727 22049 17739 22083
rect 17681 22043 17739 22049
rect 16546 21984 17448 22012
rect 16546 21956 16574 21984
rect 15562 21904 15568 21956
rect 15620 21944 15626 21956
rect 16482 21944 16488 21956
rect 15620 21916 16488 21944
rect 15620 21904 15626 21916
rect 16482 21904 16488 21916
rect 16540 21916 16574 21956
rect 16540 21904 16546 21916
rect 14274 21836 14280 21888
rect 14332 21876 14338 21888
rect 15381 21879 15439 21885
rect 15381 21876 15393 21879
rect 14332 21848 15393 21876
rect 14332 21836 14338 21848
rect 15381 21845 15393 21848
rect 15427 21845 15439 21879
rect 15381 21839 15439 21845
rect 17037 21879 17095 21885
rect 17037 21845 17049 21879
rect 17083 21876 17095 21879
rect 17126 21876 17132 21888
rect 17083 21848 17132 21876
rect 17083 21845 17095 21848
rect 17037 21839 17095 21845
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 17696 21876 17724 22043
rect 17880 22012 17908 22120
rect 17972 22120 18613 22148
rect 17972 22089 18000 22120
rect 18601 22117 18613 22120
rect 18647 22117 18659 22151
rect 18601 22111 18659 22117
rect 18966 22108 18972 22160
rect 19024 22148 19030 22160
rect 20180 22148 20208 22179
rect 20438 22176 20444 22228
rect 20496 22216 20502 22228
rect 23474 22216 23480 22228
rect 20496 22188 23480 22216
rect 20496 22176 20502 22188
rect 23474 22176 23480 22188
rect 23532 22216 23538 22228
rect 24670 22216 24676 22228
rect 23532 22188 24676 22216
rect 23532 22176 23538 22188
rect 24670 22176 24676 22188
rect 24728 22176 24734 22228
rect 25130 22176 25136 22228
rect 25188 22176 25194 22228
rect 25314 22176 25320 22228
rect 25372 22176 25378 22228
rect 27430 22216 27436 22228
rect 26068 22188 27436 22216
rect 21542 22157 21548 22160
rect 20533 22151 20591 22157
rect 20533 22148 20545 22151
rect 19024 22120 19196 22148
rect 20180 22120 20545 22148
rect 19024 22108 19030 22120
rect 17957 22083 18015 22089
rect 17957 22049 17969 22083
rect 18003 22049 18015 22083
rect 17957 22043 18015 22049
rect 18141 22083 18199 22089
rect 18141 22049 18153 22083
rect 18187 22080 18199 22083
rect 18414 22080 18420 22092
rect 18187 22052 18420 22080
rect 18187 22049 18199 22052
rect 18141 22043 18199 22049
rect 18414 22040 18420 22052
rect 18472 22040 18478 22092
rect 18785 22083 18843 22089
rect 18785 22049 18797 22083
rect 18831 22080 18843 22083
rect 18874 22080 18880 22092
rect 18831 22052 18880 22080
rect 18831 22049 18843 22052
rect 18785 22043 18843 22049
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 19058 22089 19064 22092
rect 19052 22043 19064 22089
rect 19058 22040 19064 22043
rect 19116 22040 19122 22092
rect 19168 22080 19196 22120
rect 20533 22117 20545 22120
rect 20579 22148 20591 22151
rect 21536 22148 21548 22157
rect 20579 22120 21404 22148
rect 21503 22120 21548 22148
rect 20579 22117 20591 22120
rect 20533 22111 20591 22117
rect 19168 22052 19840 22080
rect 18233 22015 18291 22021
rect 18233 22012 18245 22015
rect 17880 21984 18245 22012
rect 18233 21981 18245 21984
rect 18279 21981 18291 22015
rect 19812 22012 19840 22052
rect 20162 22040 20168 22092
rect 20220 22080 20226 22092
rect 20438 22080 20444 22092
rect 20220 22052 20444 22080
rect 20220 22040 20226 22052
rect 20438 22040 20444 22052
rect 20496 22040 20502 22092
rect 20625 22083 20683 22089
rect 20625 22049 20637 22083
rect 20671 22049 20683 22083
rect 20625 22043 20683 22049
rect 19812 21984 20392 22012
rect 18233 21975 18291 21981
rect 17865 21947 17923 21953
rect 17865 21913 17877 21947
rect 17911 21944 17923 21947
rect 17954 21944 17960 21956
rect 17911 21916 17960 21944
rect 17911 21913 17923 21916
rect 17865 21907 17923 21913
rect 17954 21904 17960 21916
rect 18012 21904 18018 21956
rect 19978 21876 19984 21888
rect 17696 21848 19984 21876
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 20254 21836 20260 21888
rect 20312 21836 20318 21888
rect 20364 21876 20392 21984
rect 20438 21904 20444 21956
rect 20496 21944 20502 21956
rect 20640 21944 20668 22043
rect 20714 22040 20720 22092
rect 20772 22089 20778 22092
rect 20772 22083 20801 22089
rect 20789 22049 20801 22083
rect 21376 22080 21404 22120
rect 21536 22111 21548 22120
rect 21542 22108 21548 22111
rect 21600 22108 21606 22160
rect 23198 22108 23204 22160
rect 23256 22148 23262 22160
rect 23354 22151 23412 22157
rect 23354 22148 23366 22151
rect 23256 22120 23366 22148
rect 23256 22108 23262 22120
rect 23354 22117 23366 22120
rect 23400 22117 23412 22151
rect 23354 22111 23412 22117
rect 25958 22108 25964 22160
rect 26016 22108 26022 22160
rect 26068 22092 26096 22188
rect 27430 22176 27436 22188
rect 27488 22176 27494 22228
rect 28166 22216 28172 22228
rect 27908 22188 28172 22216
rect 26421 22151 26479 22157
rect 26421 22117 26433 22151
rect 26467 22148 26479 22151
rect 26602 22148 26608 22160
rect 26467 22120 26608 22148
rect 26467 22117 26479 22120
rect 26421 22111 26479 22117
rect 26602 22108 26608 22120
rect 26660 22108 26666 22160
rect 27154 22148 27160 22160
rect 26712 22120 27160 22148
rect 22830 22080 22836 22092
rect 21376 22052 22836 22080
rect 20772 22043 20801 22049
rect 20772 22040 20778 22043
rect 22830 22040 22836 22052
rect 22888 22040 22894 22092
rect 23106 22040 23112 22092
rect 23164 22040 23170 22092
rect 24394 22080 24400 22092
rect 23216 22052 24400 22080
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 22012 20959 22015
rect 20947 21984 21036 22012
rect 20947 21981 20959 21984
rect 20901 21975 20959 21981
rect 20496 21916 20668 21944
rect 20496 21904 20502 21916
rect 21008 21876 21036 21984
rect 21266 21972 21272 22024
rect 21324 21972 21330 22024
rect 23216 22012 23244 22052
rect 24394 22040 24400 22052
rect 24452 22080 24458 22092
rect 25225 22083 25283 22089
rect 25225 22080 25237 22083
rect 24452 22052 25237 22080
rect 24452 22040 24458 22052
rect 25225 22049 25237 22052
rect 25271 22080 25283 22083
rect 25498 22080 25504 22092
rect 25271 22052 25504 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 25498 22040 25504 22052
rect 25556 22040 25562 22092
rect 26050 22040 26056 22092
rect 26108 22040 26114 22092
rect 26237 22083 26295 22089
rect 26237 22049 26249 22083
rect 26283 22080 26295 22083
rect 26326 22080 26332 22092
rect 26283 22052 26332 22080
rect 26283 22049 26295 22052
rect 26237 22043 26295 22049
rect 26326 22040 26332 22052
rect 26384 22080 26390 22092
rect 26712 22080 26740 22120
rect 27154 22108 27160 22120
rect 27212 22108 27218 22160
rect 27798 22108 27804 22160
rect 27856 22148 27862 22160
rect 27908 22148 27936 22188
rect 28166 22176 28172 22188
rect 28224 22176 28230 22228
rect 27856 22120 27936 22148
rect 27856 22108 27862 22120
rect 28031 22117 28089 22123
rect 28031 22114 28043 22117
rect 28016 22092 28043 22114
rect 26384 22052 26740 22080
rect 26384 22040 26390 22052
rect 26786 22040 26792 22092
rect 26844 22040 26850 22092
rect 26881 22083 26939 22089
rect 26881 22049 26893 22083
rect 26927 22080 26939 22083
rect 26970 22080 26976 22092
rect 26927 22052 26976 22080
rect 26927 22049 26939 22052
rect 26881 22043 26939 22049
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 27341 22083 27399 22089
rect 27341 22049 27353 22083
rect 27387 22080 27399 22083
rect 27522 22080 27528 22092
rect 27387 22052 27528 22080
rect 27387 22049 27399 22052
rect 27341 22043 27399 22049
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 27617 22083 27675 22089
rect 27617 22049 27629 22083
rect 27663 22080 27675 22083
rect 27890 22080 27896 22092
rect 27663 22052 27896 22080
rect 27663 22049 27675 22052
rect 27617 22043 27675 22049
rect 27890 22040 27896 22052
rect 27948 22040 27954 22092
rect 27982 22040 27988 22092
rect 28040 22083 28043 22092
rect 28077 22083 28089 22117
rect 28040 22077 28089 22083
rect 28040 22040 28046 22077
rect 28442 22040 28448 22092
rect 28500 22040 28506 22092
rect 28718 22089 28724 22092
rect 28712 22043 28724 22089
rect 28718 22040 28724 22043
rect 28776 22040 28782 22092
rect 23150 21984 23244 22012
rect 24673 22015 24731 22021
rect 22649 21947 22707 21953
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 23150 21944 23178 21984
rect 24673 21981 24685 22015
rect 24719 22012 24731 22015
rect 26418 22012 26424 22024
rect 24719 21984 26424 22012
rect 24719 21981 24731 21984
rect 24673 21975 24731 21981
rect 26418 21972 26424 21984
rect 26476 22012 26482 22024
rect 26513 22015 26571 22021
rect 26513 22012 26525 22015
rect 26476 21984 26525 22012
rect 26476 21972 26482 21984
rect 26513 21981 26525 21984
rect 26559 21981 26571 22015
rect 26513 21975 26571 21981
rect 27430 21972 27436 22024
rect 27488 21972 27494 22024
rect 25041 21947 25099 21953
rect 25041 21944 25053 21947
rect 22695 21916 23178 21944
rect 24044 21916 25053 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 22738 21876 22744 21888
rect 20364 21848 22744 21876
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 22830 21836 22836 21888
rect 22888 21876 22894 21888
rect 24044 21876 24072 21916
rect 25041 21913 25053 21916
rect 25087 21944 25099 21947
rect 25406 21944 25412 21956
rect 25087 21916 25412 21944
rect 25087 21913 25099 21916
rect 25041 21907 25099 21913
rect 25406 21904 25412 21916
rect 25464 21904 25470 21956
rect 25501 21947 25559 21953
rect 25501 21913 25513 21947
rect 25547 21944 25559 21947
rect 26053 21947 26111 21953
rect 26053 21944 26065 21947
rect 25547 21916 26065 21944
rect 25547 21913 25559 21916
rect 25501 21907 25559 21913
rect 26053 21913 26065 21916
rect 26099 21913 26111 21947
rect 26694 21944 26700 21956
rect 26053 21907 26111 21913
rect 26160 21916 26700 21944
rect 22888 21848 24072 21876
rect 24489 21879 24547 21885
rect 22888 21836 22894 21848
rect 24489 21845 24501 21879
rect 24535 21876 24547 21879
rect 24854 21876 24860 21888
rect 24535 21848 24860 21876
rect 24535 21845 24547 21848
rect 24489 21839 24547 21845
rect 24854 21836 24860 21848
rect 24912 21836 24918 21888
rect 25590 21836 25596 21888
rect 25648 21836 25654 21888
rect 25685 21879 25743 21885
rect 25685 21845 25697 21879
rect 25731 21876 25743 21879
rect 26160 21876 26188 21916
rect 26694 21904 26700 21916
rect 26752 21904 26758 21956
rect 27065 21947 27123 21953
rect 27065 21913 27077 21947
rect 27111 21944 27123 21947
rect 27111 21916 27384 21944
rect 27111 21913 27123 21916
rect 27065 21907 27123 21913
rect 25731 21848 26188 21876
rect 25731 21845 25743 21848
rect 25685 21839 25743 21845
rect 26418 21836 26424 21888
rect 26476 21876 26482 21888
rect 27356 21885 27384 21916
rect 27157 21879 27215 21885
rect 27157 21876 27169 21879
rect 26476 21848 27169 21876
rect 26476 21836 26482 21848
rect 27157 21845 27169 21848
rect 27203 21845 27215 21879
rect 27157 21839 27215 21845
rect 27341 21879 27399 21885
rect 27341 21845 27353 21879
rect 27387 21845 27399 21879
rect 27341 21839 27399 21845
rect 27985 21879 28043 21885
rect 27985 21845 27997 21879
rect 28031 21876 28043 21879
rect 28074 21876 28080 21888
rect 28031 21848 28080 21876
rect 28031 21845 28043 21848
rect 27985 21839 28043 21845
rect 28074 21836 28080 21848
rect 28132 21836 28138 21888
rect 28169 21879 28227 21885
rect 28169 21845 28181 21879
rect 28215 21876 28227 21879
rect 28350 21876 28356 21888
rect 28215 21848 28356 21876
rect 28215 21845 28227 21848
rect 28169 21839 28227 21845
rect 28350 21836 28356 21848
rect 28408 21836 28414 21888
rect 28442 21836 28448 21888
rect 28500 21876 28506 21888
rect 29825 21879 29883 21885
rect 29825 21876 29837 21879
rect 28500 21848 29837 21876
rect 28500 21836 28506 21848
rect 29825 21845 29837 21848
rect 29871 21845 29883 21879
rect 29825 21839 29883 21845
rect 552 21786 31648 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 11436 21786
rect 11488 21734 11500 21786
rect 11552 21734 11564 21786
rect 11616 21734 11628 21786
rect 11680 21734 11692 21786
rect 11744 21734 19210 21786
rect 19262 21734 19274 21786
rect 19326 21734 19338 21786
rect 19390 21734 19402 21786
rect 19454 21734 19466 21786
rect 19518 21734 26984 21786
rect 27036 21734 27048 21786
rect 27100 21734 27112 21786
rect 27164 21734 27176 21786
rect 27228 21734 27240 21786
rect 27292 21734 31648 21786
rect 552 21712 31648 21734
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13630 21672 13636 21684
rect 13587 21644 13636 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 14550 21632 14556 21684
rect 14608 21672 14614 21684
rect 14737 21675 14795 21681
rect 14737 21672 14749 21675
rect 14608 21644 14749 21672
rect 14608 21632 14614 21644
rect 14737 21641 14749 21644
rect 14783 21641 14795 21675
rect 17770 21672 17776 21684
rect 14737 21635 14795 21641
rect 16684 21644 17776 21672
rect 14366 21536 14372 21548
rect 13924 21508 14372 21536
rect 13924 21477 13952 21508
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 15378 21536 15384 21548
rect 14568 21508 15384 21536
rect 13817 21471 13875 21477
rect 13817 21437 13829 21471
rect 13863 21437 13875 21471
rect 13817 21431 13875 21437
rect 13909 21471 13967 21477
rect 13909 21437 13921 21471
rect 13955 21437 13967 21471
rect 13909 21431 13967 21437
rect 14001 21471 14059 21477
rect 14001 21437 14013 21471
rect 14047 21468 14059 21471
rect 14090 21468 14096 21480
rect 14047 21440 14096 21468
rect 14047 21437 14059 21440
rect 14001 21431 14059 21437
rect 13832 21400 13860 21431
rect 14090 21428 14096 21440
rect 14148 21428 14154 21480
rect 14185 21471 14243 21477
rect 14185 21437 14197 21471
rect 14231 21468 14243 21471
rect 14568 21468 14596 21508
rect 15378 21496 15384 21508
rect 15436 21496 15442 21548
rect 16684 21536 16712 21644
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 19429 21675 19487 21681
rect 19429 21672 19441 21675
rect 19116 21644 19441 21672
rect 19116 21632 19122 21644
rect 19429 21641 19441 21644
rect 19475 21641 19487 21675
rect 19429 21635 19487 21641
rect 20070 21632 20076 21684
rect 20128 21672 20134 21684
rect 20438 21672 20444 21684
rect 20128 21644 20444 21672
rect 20128 21632 20134 21644
rect 20438 21632 20444 21644
rect 20496 21632 20502 21684
rect 21266 21632 21272 21684
rect 21324 21672 21330 21684
rect 21453 21675 21511 21681
rect 21453 21672 21465 21675
rect 21324 21644 21465 21672
rect 21324 21632 21330 21644
rect 21453 21641 21465 21644
rect 21499 21641 21511 21675
rect 22094 21672 22100 21684
rect 21453 21635 21511 21641
rect 21652 21644 22100 21672
rect 20254 21564 20260 21616
rect 20312 21564 20318 21616
rect 20272 21536 20300 21564
rect 16592 21508 16712 21536
rect 19628 21508 20300 21536
rect 14231 21440 14596 21468
rect 14231 21437 14243 21440
rect 14185 21431 14243 21437
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 16592 21477 16620 21508
rect 17126 21477 17132 21480
rect 14829 21471 14887 21477
rect 14829 21468 14841 21471
rect 14700 21440 14841 21468
rect 14700 21428 14706 21440
rect 14829 21437 14841 21440
rect 14875 21437 14887 21471
rect 14829 21431 14887 21437
rect 16393 21471 16451 21477
rect 16393 21437 16405 21471
rect 16439 21468 16451 21471
rect 16577 21471 16635 21477
rect 16577 21468 16589 21471
rect 16439 21440 16589 21468
rect 16439 21437 16451 21440
rect 16393 21431 16451 21437
rect 16577 21437 16589 21440
rect 16623 21437 16635 21471
rect 16577 21431 16635 21437
rect 16669 21471 16727 21477
rect 16669 21437 16681 21471
rect 16715 21468 16727 21471
rect 16853 21471 16911 21477
rect 16853 21468 16865 21471
rect 16715 21440 16865 21468
rect 16715 21437 16727 21440
rect 16669 21431 16727 21437
rect 16853 21437 16865 21440
rect 16899 21437 16911 21471
rect 17120 21468 17132 21477
rect 17087 21440 17132 21468
rect 16853 21431 16911 21437
rect 17120 21431 17132 21440
rect 17126 21428 17132 21431
rect 17184 21428 17190 21480
rect 19628 21477 19656 21508
rect 19245 21471 19303 21477
rect 19245 21468 19257 21471
rect 18432 21440 19257 21468
rect 15654 21400 15660 21412
rect 13832 21372 15660 21400
rect 15654 21360 15660 21372
rect 15712 21360 15718 21412
rect 18432 21344 18460 21440
rect 19245 21437 19257 21440
rect 19291 21437 19303 21471
rect 19245 21431 19303 21437
rect 19613 21471 19671 21477
rect 19613 21437 19625 21471
rect 19659 21437 19671 21471
rect 19613 21431 19671 21437
rect 19797 21471 19855 21477
rect 19797 21437 19809 21471
rect 19843 21437 19855 21471
rect 19797 21431 19855 21437
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21468 20315 21471
rect 20806 21468 20812 21480
rect 20303 21440 20812 21468
rect 20303 21437 20315 21440
rect 20257 21431 20315 21437
rect 19812 21344 19840 21431
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 21545 21471 21603 21477
rect 21545 21437 21557 21471
rect 21591 21468 21603 21471
rect 21652 21468 21680 21644
rect 22094 21632 22100 21644
rect 22152 21672 22158 21684
rect 23014 21672 23020 21684
rect 22152 21644 23020 21672
rect 22152 21632 22158 21644
rect 23014 21632 23020 21644
rect 23072 21632 23078 21684
rect 23198 21632 23204 21684
rect 23256 21632 23262 21684
rect 24210 21632 24216 21684
rect 24268 21672 24274 21684
rect 24489 21675 24547 21681
rect 24489 21672 24501 21675
rect 24268 21644 24501 21672
rect 24268 21632 24274 21644
rect 24489 21641 24501 21644
rect 24535 21641 24547 21675
rect 24489 21635 24547 21641
rect 25682 21632 25688 21684
rect 25740 21672 25746 21684
rect 26329 21675 26387 21681
rect 26329 21672 26341 21675
rect 25740 21644 26341 21672
rect 25740 21632 25746 21644
rect 26329 21641 26341 21644
rect 26375 21641 26387 21675
rect 26329 21635 26387 21641
rect 27246 21632 27252 21684
rect 27304 21672 27310 21684
rect 27614 21672 27620 21684
rect 27304 21644 27620 21672
rect 27304 21632 27310 21644
rect 27614 21632 27620 21644
rect 27672 21632 27678 21684
rect 28718 21632 28724 21684
rect 28776 21632 28782 21684
rect 23109 21607 23167 21613
rect 23109 21573 23121 21607
rect 23155 21573 23167 21607
rect 23109 21567 23167 21573
rect 23492 21576 25452 21604
rect 23124 21536 23152 21567
rect 23492 21536 23520 21576
rect 23124 21508 23520 21536
rect 23566 21496 23572 21548
rect 23624 21496 23630 21548
rect 23860 21545 23888 21576
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21505 23903 21539
rect 23845 21499 23903 21505
rect 24578 21496 24584 21548
rect 24636 21496 24642 21548
rect 24762 21496 24768 21548
rect 24820 21536 24826 21548
rect 25424 21536 25452 21576
rect 25498 21564 25504 21616
rect 25556 21604 25562 21616
rect 25556 21576 25820 21604
rect 25556 21564 25562 21576
rect 24820 21508 25084 21536
rect 25424 21508 25636 21536
rect 24820 21496 24826 21508
rect 21591 21440 21680 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 21726 21428 21732 21480
rect 21784 21428 21790 21480
rect 21996 21471 22054 21477
rect 21996 21437 22008 21471
rect 22042 21468 22054 21471
rect 22278 21468 22284 21480
rect 22042 21440 22284 21468
rect 22042 21437 22054 21440
rect 21996 21431 22054 21437
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 23198 21428 23204 21480
rect 23256 21468 23262 21480
rect 23385 21471 23443 21477
rect 23385 21468 23397 21471
rect 23256 21440 23397 21468
rect 23256 21428 23262 21440
rect 23385 21437 23397 21440
rect 23431 21437 23443 21471
rect 24857 21471 24915 21477
rect 24857 21468 24869 21471
rect 23385 21431 23443 21437
rect 23492 21465 24532 21468
rect 24596 21465 24869 21468
rect 23492 21440 24869 21465
rect 19978 21360 19984 21412
rect 20036 21400 20042 21412
rect 20036 21372 21588 21400
rect 20036 21360 20042 21372
rect 16114 21292 16120 21344
rect 16172 21332 16178 21344
rect 16301 21335 16359 21341
rect 16301 21332 16313 21335
rect 16172 21304 16313 21332
rect 16172 21292 16178 21304
rect 16301 21301 16313 21304
rect 16347 21301 16359 21335
rect 16301 21295 16359 21301
rect 18233 21335 18291 21341
rect 18233 21301 18245 21335
rect 18279 21332 18291 21335
rect 18414 21332 18420 21344
rect 18279 21304 18420 21332
rect 18279 21301 18291 21304
rect 18233 21295 18291 21301
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 18690 21292 18696 21344
rect 18748 21292 18754 21344
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 20073 21335 20131 21341
rect 20073 21332 20085 21335
rect 19852 21304 20085 21332
rect 19852 21292 19858 21304
rect 20073 21301 20085 21304
rect 20119 21301 20131 21335
rect 20073 21295 20131 21301
rect 20162 21292 20168 21344
rect 20220 21332 20226 21344
rect 20622 21332 20628 21344
rect 20220 21304 20628 21332
rect 20220 21292 20226 21304
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 21560 21332 21588 21372
rect 21634 21360 21640 21412
rect 21692 21400 21698 21412
rect 23492 21400 23520 21440
rect 24504 21437 24624 21440
rect 24857 21437 24869 21440
rect 24903 21437 24915 21471
rect 24857 21431 24915 21437
rect 24946 21428 24952 21480
rect 25004 21428 25010 21480
rect 25056 21477 25084 21508
rect 25041 21471 25099 21477
rect 25041 21437 25053 21471
rect 25087 21437 25099 21471
rect 25041 21431 25099 21437
rect 25130 21428 25136 21480
rect 25188 21468 25194 21480
rect 25409 21471 25467 21477
rect 25409 21468 25421 21471
rect 25188 21440 25421 21468
rect 25188 21428 25194 21440
rect 25409 21437 25421 21440
rect 25455 21437 25467 21471
rect 25409 21431 25467 21437
rect 25498 21428 25504 21480
rect 25556 21468 25562 21480
rect 25608 21477 25636 21508
rect 25682 21496 25688 21548
rect 25740 21496 25746 21548
rect 25792 21545 25820 21576
rect 25958 21564 25964 21616
rect 26016 21604 26022 21616
rect 26016 21576 26280 21604
rect 26016 21564 26022 21576
rect 26252 21545 26280 21576
rect 26418 21564 26424 21616
rect 26476 21564 26482 21616
rect 27985 21607 28043 21613
rect 27985 21573 27997 21607
rect 28031 21604 28043 21607
rect 28166 21604 28172 21616
rect 28031 21576 28172 21604
rect 28031 21573 28043 21576
rect 27985 21567 28043 21573
rect 28166 21564 28172 21576
rect 28224 21604 28230 21616
rect 28442 21604 28448 21616
rect 28224 21576 28448 21604
rect 28224 21564 28230 21576
rect 28442 21564 28448 21576
rect 28500 21564 28506 21616
rect 25777 21539 25835 21545
rect 25777 21505 25789 21539
rect 25823 21505 25835 21539
rect 25777 21499 25835 21505
rect 26237 21539 26295 21545
rect 26237 21505 26249 21539
rect 26283 21505 26295 21539
rect 26237 21499 26295 21505
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21536 27307 21539
rect 27295 21508 28304 21536
rect 27295 21505 27307 21508
rect 27249 21499 27307 21505
rect 25593 21471 25651 21477
rect 25593 21468 25605 21471
rect 25556 21440 25605 21468
rect 25556 21428 25562 21440
rect 25593 21437 25605 21440
rect 25639 21437 25651 21471
rect 25593 21431 25651 21437
rect 25961 21471 26019 21477
rect 25961 21437 25973 21471
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 21692 21372 23520 21400
rect 21692 21360 21698 21372
rect 24670 21360 24676 21412
rect 24728 21409 24734 21412
rect 24728 21403 24777 21409
rect 24728 21369 24731 21403
rect 24765 21369 24777 21403
rect 24728 21363 24777 21369
rect 24728 21360 24734 21363
rect 25314 21360 25320 21412
rect 25372 21400 25378 21412
rect 25976 21400 26004 21431
rect 26510 21428 26516 21480
rect 26568 21428 26574 21480
rect 26786 21428 26792 21480
rect 26844 21468 26850 21480
rect 27157 21471 27215 21477
rect 27157 21468 27169 21471
rect 26844 21440 27169 21468
rect 26844 21428 26850 21440
rect 27157 21437 27169 21440
rect 27203 21468 27215 21471
rect 27433 21471 27491 21477
rect 27433 21468 27445 21471
rect 27203 21440 27445 21468
rect 27203 21437 27215 21440
rect 27157 21431 27215 21437
rect 27433 21437 27445 21440
rect 27479 21437 27491 21471
rect 27433 21431 27491 21437
rect 27798 21428 27804 21480
rect 27856 21428 27862 21480
rect 28276 21477 28304 21508
rect 28077 21471 28135 21477
rect 28077 21437 28089 21471
rect 28123 21437 28135 21471
rect 28077 21431 28135 21437
rect 28261 21471 28319 21477
rect 28261 21437 28273 21471
rect 28307 21437 28319 21471
rect 28261 21431 28319 21437
rect 25372 21372 26004 21400
rect 27617 21403 27675 21409
rect 25372 21360 25378 21372
rect 27617 21369 27629 21403
rect 27663 21400 27675 21403
rect 27982 21400 27988 21412
rect 27663 21372 27988 21400
rect 27663 21369 27675 21372
rect 27617 21363 27675 21369
rect 27982 21360 27988 21372
rect 28040 21360 28046 21412
rect 28092 21400 28120 21431
rect 28350 21428 28356 21480
rect 28408 21428 28414 21480
rect 28460 21477 28488 21564
rect 28445 21471 28503 21477
rect 28445 21437 28457 21471
rect 28491 21437 28503 21471
rect 28445 21431 28503 21437
rect 28994 21428 29000 21480
rect 29052 21428 29058 21480
rect 28534 21400 28540 21412
rect 28092 21372 28540 21400
rect 28534 21360 28540 21372
rect 28592 21360 28598 21412
rect 22370 21332 22376 21344
rect 21560 21304 22376 21332
rect 22370 21292 22376 21304
rect 22428 21332 22434 21344
rect 23566 21332 23572 21344
rect 22428 21304 23572 21332
rect 22428 21292 22434 21304
rect 23566 21292 23572 21304
rect 23624 21292 23630 21344
rect 23750 21292 23756 21344
rect 23808 21332 23814 21344
rect 25225 21335 25283 21341
rect 25225 21332 25237 21335
rect 23808 21304 25237 21332
rect 23808 21292 23814 21304
rect 25225 21301 25237 21304
rect 25271 21301 25283 21335
rect 25225 21295 25283 21301
rect 25682 21292 25688 21344
rect 25740 21332 25746 21344
rect 25866 21332 25872 21344
rect 25740 21304 25872 21332
rect 25740 21292 25746 21304
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 26142 21292 26148 21344
rect 26200 21292 26206 21344
rect 27709 21335 27767 21341
rect 27709 21301 27721 21335
rect 27755 21332 27767 21335
rect 28074 21332 28080 21344
rect 27755 21304 28080 21332
rect 27755 21301 27767 21304
rect 27709 21295 27767 21301
rect 28074 21292 28080 21304
rect 28132 21292 28138 21344
rect 28810 21292 28816 21344
rect 28868 21332 28874 21344
rect 29089 21335 29147 21341
rect 29089 21332 29101 21335
rect 28868 21304 29101 21332
rect 28868 21292 28874 21304
rect 29089 21301 29101 21304
rect 29135 21301 29147 21335
rect 29089 21295 29147 21301
rect 552 21242 31648 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 12096 21242
rect 12148 21190 12160 21242
rect 12212 21190 12224 21242
rect 12276 21190 12288 21242
rect 12340 21190 12352 21242
rect 12404 21190 19870 21242
rect 19922 21190 19934 21242
rect 19986 21190 19998 21242
rect 20050 21190 20062 21242
rect 20114 21190 20126 21242
rect 20178 21190 27644 21242
rect 27696 21190 27708 21242
rect 27760 21190 27772 21242
rect 27824 21190 27836 21242
rect 27888 21190 27900 21242
rect 27952 21190 31648 21242
rect 552 21168 31648 21190
rect 17586 21088 17592 21140
rect 17644 21088 17650 21140
rect 21726 21088 21732 21140
rect 21784 21128 21790 21140
rect 21913 21131 21971 21137
rect 21913 21128 21925 21131
rect 21784 21100 21925 21128
rect 21784 21088 21790 21100
rect 21913 21097 21925 21100
rect 21959 21097 21971 21131
rect 21913 21091 21971 21097
rect 22738 21088 22744 21140
rect 22796 21128 22802 21140
rect 23934 21128 23940 21140
rect 22796 21100 23940 21128
rect 22796 21088 22802 21100
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 25130 21088 25136 21140
rect 25188 21088 25194 21140
rect 25406 21088 25412 21140
rect 25464 21128 25470 21140
rect 26326 21128 26332 21140
rect 25464 21100 26332 21128
rect 25464 21088 25470 21100
rect 26326 21088 26332 21100
rect 26384 21088 26390 21140
rect 27246 21088 27252 21140
rect 27304 21128 27310 21140
rect 27706 21128 27712 21140
rect 27304 21100 27712 21128
rect 27304 21088 27310 21100
rect 27706 21088 27712 21100
rect 27764 21088 27770 21140
rect 27982 21088 27988 21140
rect 28040 21088 28046 21140
rect 30193 21131 30251 21137
rect 30193 21128 30205 21131
rect 28460 21100 30205 21128
rect 15933 21063 15991 21069
rect 15933 21029 15945 21063
rect 15979 21060 15991 21063
rect 16362 21063 16420 21069
rect 16362 21060 16374 21063
rect 15979 21032 16374 21060
rect 15979 21029 15991 21032
rect 15933 21023 15991 21029
rect 16362 21029 16374 21032
rect 16408 21029 16420 21063
rect 16362 21023 16420 21029
rect 17773 21063 17831 21069
rect 17773 21029 17785 21063
rect 17819 21060 17831 21063
rect 18690 21060 18696 21072
rect 17819 21032 18696 21060
rect 17819 21029 17831 21032
rect 17773 21023 17831 21029
rect 18690 21020 18696 21032
rect 18748 21020 18754 21072
rect 28460 21060 28488 21100
rect 30193 21097 30205 21100
rect 30239 21097 30251 21131
rect 30193 21091 30251 21097
rect 27448 21032 28488 21060
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20992 15347 20995
rect 15378 20992 15384 21004
rect 15335 20964 15384 20992
rect 15335 20961 15347 20964
rect 15289 20955 15347 20961
rect 15378 20952 15384 20964
rect 15436 20952 15442 21004
rect 15470 20952 15476 21004
rect 15528 20952 15534 21004
rect 15562 20952 15568 21004
rect 15620 20952 15626 21004
rect 15654 20952 15660 21004
rect 15712 20952 15718 21004
rect 16114 20952 16120 21004
rect 16172 20952 16178 21004
rect 16224 20964 17448 20992
rect 15672 20924 15700 20952
rect 16224 20924 16252 20964
rect 15672 20896 16252 20924
rect 17420 20924 17448 20964
rect 17586 20952 17592 21004
rect 17644 20992 17650 21004
rect 17954 20992 17960 21004
rect 17644 20964 17960 20992
rect 17644 20952 17650 20964
rect 17954 20952 17960 20964
rect 18012 20952 18018 21004
rect 22005 20995 22063 21001
rect 22005 20961 22017 20995
rect 22051 20992 22063 20995
rect 22094 20992 22100 21004
rect 22051 20964 22100 20992
rect 22051 20961 22063 20964
rect 22005 20955 22063 20961
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 24765 20995 24823 21001
rect 24765 20961 24777 20995
rect 24811 20992 24823 20995
rect 27338 20992 27344 21004
rect 24811 20964 27344 20992
rect 24811 20961 24823 20964
rect 24765 20955 24823 20961
rect 27338 20952 27344 20964
rect 27396 20992 27402 21004
rect 27448 21001 27476 21032
rect 27433 20995 27491 21001
rect 27433 20992 27445 20995
rect 27396 20964 27445 20992
rect 27396 20952 27402 20964
rect 27433 20961 27445 20964
rect 27479 20961 27491 20995
rect 27433 20955 27491 20961
rect 27617 20995 27675 21001
rect 27617 20961 27629 20995
rect 27663 20961 27675 20995
rect 27617 20955 27675 20961
rect 18598 20924 18604 20936
rect 17420 20896 18604 20924
rect 18598 20884 18604 20896
rect 18656 20884 18662 20936
rect 24854 20884 24860 20936
rect 24912 20884 24918 20936
rect 27632 20924 27660 20955
rect 27798 20952 27804 21004
rect 27856 20952 27862 21004
rect 28074 20952 28080 21004
rect 28132 20952 28138 21004
rect 28460 21001 28488 21032
rect 28721 21063 28779 21069
rect 28721 21029 28733 21063
rect 28767 21060 28779 21063
rect 29058 21063 29116 21069
rect 29058 21060 29070 21063
rect 28767 21032 29070 21060
rect 28767 21029 28779 21032
rect 28721 21023 28779 21029
rect 29058 21029 29070 21032
rect 29104 21029 29116 21063
rect 29058 21023 29116 21029
rect 28261 20995 28319 21001
rect 28261 20961 28273 20995
rect 28307 20961 28319 20995
rect 28261 20955 28319 20961
rect 28353 20995 28411 21001
rect 28353 20961 28365 20995
rect 28399 20961 28411 20995
rect 28353 20955 28411 20961
rect 28445 20995 28503 21001
rect 28445 20961 28457 20995
rect 28491 20961 28503 20995
rect 28445 20955 28503 20961
rect 27982 20924 27988 20936
rect 27632 20896 27988 20924
rect 27982 20884 27988 20896
rect 28040 20884 28046 20936
rect 17494 20748 17500 20800
rect 17552 20748 17558 20800
rect 23934 20748 23940 20800
rect 23992 20788 23998 20800
rect 24578 20788 24584 20800
rect 23992 20760 24584 20788
rect 23992 20748 23998 20760
rect 24578 20748 24584 20760
rect 24636 20748 24642 20800
rect 28276 20788 28304 20955
rect 28368 20856 28396 20955
rect 28810 20952 28816 21004
rect 28868 20952 28874 21004
rect 28442 20856 28448 20868
rect 28368 20828 28448 20856
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 28626 20788 28632 20800
rect 28276 20760 28632 20788
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 552 20698 31648 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 11436 20698
rect 11488 20646 11500 20698
rect 11552 20646 11564 20698
rect 11616 20646 11628 20698
rect 11680 20646 11692 20698
rect 11744 20646 19210 20698
rect 19262 20646 19274 20698
rect 19326 20646 19338 20698
rect 19390 20646 19402 20698
rect 19454 20646 19466 20698
rect 19518 20646 26984 20698
rect 27036 20646 27048 20698
rect 27100 20646 27112 20698
rect 27164 20646 27176 20698
rect 27228 20646 27240 20698
rect 27292 20646 31648 20698
rect 552 20624 31648 20646
rect 15470 20544 15476 20596
rect 15528 20584 15534 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 15528 20556 15853 20584
rect 15528 20544 15534 20556
rect 15841 20553 15853 20556
rect 15887 20553 15899 20587
rect 15841 20547 15899 20553
rect 20364 20556 22968 20584
rect 18230 20476 18236 20528
rect 18288 20516 18294 20528
rect 20364 20516 20392 20556
rect 18288 20488 20392 20516
rect 18288 20476 18294 20488
rect 20254 20448 20260 20460
rect 18892 20420 19656 20448
rect 18892 20392 18920 20420
rect 16025 20383 16083 20389
rect 16025 20349 16037 20383
rect 16071 20380 16083 20383
rect 16666 20380 16672 20392
rect 16071 20352 16672 20380
rect 16071 20349 16083 20352
rect 16025 20343 16083 20349
rect 16666 20340 16672 20352
rect 16724 20380 16730 20392
rect 17494 20380 17500 20392
rect 16724 20352 17500 20380
rect 16724 20340 16730 20352
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 17586 20340 17592 20392
rect 17644 20380 17650 20392
rect 17773 20383 17831 20389
rect 17773 20380 17785 20383
rect 17644 20352 17785 20380
rect 17644 20340 17650 20352
rect 17773 20349 17785 20352
rect 17819 20349 17831 20383
rect 17773 20343 17831 20349
rect 18417 20383 18475 20389
rect 18417 20349 18429 20383
rect 18463 20380 18475 20383
rect 18874 20380 18880 20392
rect 18463 20352 18880 20380
rect 18463 20349 18475 20352
rect 18417 20343 18475 20349
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 19242 20340 19248 20392
rect 19300 20340 19306 20392
rect 19628 20389 19656 20420
rect 19904 20420 20260 20448
rect 19904 20389 19932 20420
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 20364 20457 20392 20488
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 22940 20457 22968 20556
rect 25590 20544 25596 20596
rect 25648 20584 25654 20596
rect 25685 20587 25743 20593
rect 25685 20584 25697 20587
rect 25648 20556 25697 20584
rect 25648 20544 25654 20556
rect 25685 20553 25697 20556
rect 25731 20553 25743 20587
rect 25685 20547 25743 20553
rect 25774 20544 25780 20596
rect 25832 20584 25838 20596
rect 26145 20587 26203 20593
rect 26145 20584 26157 20587
rect 25832 20556 26157 20584
rect 25832 20544 25838 20556
rect 26145 20553 26157 20556
rect 26191 20553 26203 20587
rect 26145 20547 26203 20553
rect 28074 20544 28080 20596
rect 28132 20584 28138 20596
rect 28169 20587 28227 20593
rect 28169 20584 28181 20587
rect 28132 20556 28181 20584
rect 28132 20544 28138 20556
rect 28169 20553 28181 20556
rect 28215 20553 28227 20587
rect 28169 20547 28227 20553
rect 24946 20476 24952 20528
rect 25004 20516 25010 20528
rect 27798 20516 27804 20528
rect 25004 20488 27804 20516
rect 25004 20476 25010 20488
rect 27798 20476 27804 20488
rect 27856 20516 27862 20528
rect 28718 20516 28724 20528
rect 27856 20488 28724 20516
rect 27856 20476 27862 20488
rect 28718 20476 28724 20488
rect 28776 20476 28782 20528
rect 22925 20451 22983 20457
rect 20680 20420 22692 20448
rect 20680 20408 20686 20420
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 19889 20383 19947 20389
rect 19889 20349 19901 20383
rect 19935 20349 19947 20383
rect 19889 20343 19947 20349
rect 20073 20383 20131 20389
rect 20073 20349 20085 20383
rect 20119 20380 20131 20383
rect 20806 20380 20812 20392
rect 20119 20352 20812 20380
rect 20119 20349 20131 20352
rect 20073 20343 20131 20349
rect 20806 20340 20812 20352
rect 20864 20380 20870 20392
rect 21634 20380 21640 20392
rect 20864 20352 21640 20380
rect 20864 20340 20870 20352
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 22002 20340 22008 20392
rect 22060 20340 22066 20392
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20349 22523 20383
rect 22465 20343 22523 20349
rect 16209 20315 16267 20321
rect 16209 20281 16221 20315
rect 16255 20312 16267 20315
rect 16574 20312 16580 20324
rect 16255 20284 16580 20312
rect 16255 20281 16267 20284
rect 16209 20275 16267 20281
rect 16574 20272 16580 20284
rect 16632 20312 16638 20324
rect 17604 20312 17632 20340
rect 16632 20284 17632 20312
rect 17957 20315 18015 20321
rect 16632 20272 16638 20284
rect 17957 20281 17969 20315
rect 18003 20312 18015 20315
rect 18693 20315 18751 20321
rect 18693 20312 18705 20315
rect 18003 20284 18705 20312
rect 18003 20281 18015 20284
rect 17957 20275 18015 20281
rect 18693 20281 18705 20284
rect 18739 20281 18751 20315
rect 18693 20275 18751 20281
rect 19981 20315 20039 20321
rect 19981 20281 19993 20315
rect 20027 20281 20039 20315
rect 19981 20275 20039 20281
rect 20211 20315 20269 20321
rect 20211 20281 20223 20315
rect 20257 20312 20269 20315
rect 20714 20312 20720 20324
rect 20257 20284 20720 20312
rect 20257 20281 20269 20284
rect 20211 20275 20269 20281
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18141 20247 18199 20253
rect 18141 20244 18153 20247
rect 18104 20216 18153 20244
rect 18104 20204 18110 20216
rect 18141 20213 18153 20216
rect 18187 20213 18199 20247
rect 18141 20207 18199 20213
rect 18322 20204 18328 20256
rect 18380 20204 18386 20256
rect 19150 20204 19156 20256
rect 19208 20244 19214 20256
rect 19521 20247 19579 20253
rect 19521 20244 19533 20247
rect 19208 20216 19533 20244
rect 19208 20204 19214 20216
rect 19521 20213 19533 20216
rect 19567 20213 19579 20247
rect 19521 20207 19579 20213
rect 19702 20204 19708 20256
rect 19760 20204 19766 20256
rect 19996 20244 20024 20275
rect 20714 20272 20720 20284
rect 20772 20312 20778 20324
rect 21726 20312 21732 20324
rect 20772 20284 21732 20312
rect 20772 20272 20778 20284
rect 21726 20272 21732 20284
rect 21784 20272 21790 20324
rect 22480 20312 22508 20343
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 22664 20389 22692 20420
rect 22925 20417 22937 20451
rect 22971 20448 22983 20451
rect 23290 20448 23296 20460
rect 22971 20420 23296 20448
rect 22971 20417 22983 20420
rect 22925 20411 22983 20417
rect 23290 20408 23296 20420
rect 23348 20408 23354 20460
rect 26602 20448 26608 20460
rect 24136 20420 26608 20448
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20349 22707 20383
rect 22649 20343 22707 20349
rect 22787 20383 22845 20389
rect 22787 20349 22799 20383
rect 22833 20380 22845 20383
rect 23474 20380 23480 20392
rect 22833 20352 23480 20380
rect 22833 20349 22845 20352
rect 22787 20343 22845 20349
rect 23474 20340 23480 20352
rect 23532 20380 23538 20392
rect 24026 20380 24032 20392
rect 23532 20352 24032 20380
rect 23532 20340 23538 20352
rect 24026 20340 24032 20352
rect 24084 20340 24090 20392
rect 23934 20312 23940 20324
rect 22480 20284 23940 20312
rect 23934 20272 23940 20284
rect 23992 20272 23998 20324
rect 20530 20244 20536 20256
rect 19996 20216 20536 20244
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 22094 20204 22100 20256
rect 22152 20204 22158 20256
rect 22186 20204 22192 20256
rect 22244 20244 22250 20256
rect 22281 20247 22339 20253
rect 22281 20244 22293 20247
rect 22244 20216 22293 20244
rect 22244 20204 22250 20216
rect 22281 20213 22293 20216
rect 22327 20213 22339 20247
rect 22281 20207 22339 20213
rect 22554 20204 22560 20256
rect 22612 20244 22618 20256
rect 24136 20244 24164 20420
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 25332 20389 25360 20420
rect 26602 20408 26608 20420
rect 26660 20408 26666 20460
rect 25041 20383 25099 20389
rect 25041 20380 25053 20383
rect 24268 20352 25053 20380
rect 24268 20340 24274 20352
rect 25041 20349 25053 20352
rect 25087 20349 25099 20383
rect 25041 20343 25099 20349
rect 25189 20383 25247 20389
rect 25189 20349 25201 20383
rect 25235 20380 25247 20383
rect 25317 20383 25375 20389
rect 25235 20349 25268 20380
rect 25189 20343 25268 20349
rect 25317 20349 25329 20383
rect 25363 20349 25375 20383
rect 25317 20343 25375 20349
rect 22612 20216 24164 20244
rect 25240 20244 25268 20343
rect 25498 20340 25504 20392
rect 25556 20389 25562 20392
rect 25556 20380 25564 20389
rect 26053 20383 26111 20389
rect 25556 20352 25601 20380
rect 25556 20343 25564 20352
rect 26053 20349 26065 20383
rect 26099 20380 26111 20383
rect 27982 20380 27988 20392
rect 26099 20352 27988 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 25556 20340 25562 20343
rect 27982 20340 27988 20352
rect 28040 20340 28046 20392
rect 28261 20383 28319 20389
rect 28261 20349 28273 20383
rect 28307 20380 28319 20383
rect 28350 20380 28356 20392
rect 28307 20352 28356 20380
rect 28307 20349 28319 20352
rect 28261 20343 28319 20349
rect 28350 20340 28356 20352
rect 28408 20340 28414 20392
rect 25409 20315 25467 20321
rect 25409 20281 25421 20315
rect 25455 20312 25467 20315
rect 25682 20312 25688 20324
rect 25455 20284 25688 20312
rect 25455 20281 25467 20284
rect 25409 20275 25467 20281
rect 25682 20272 25688 20284
rect 25740 20272 25746 20324
rect 25866 20272 25872 20324
rect 25924 20312 25930 20324
rect 27430 20312 27436 20324
rect 25924 20284 27436 20312
rect 25924 20272 25930 20284
rect 27430 20272 27436 20284
rect 27488 20272 27494 20324
rect 26050 20244 26056 20256
rect 25240 20216 26056 20244
rect 22612 20204 22618 20216
rect 26050 20204 26056 20216
rect 26108 20204 26114 20256
rect 27706 20204 27712 20256
rect 27764 20244 27770 20256
rect 28074 20244 28080 20256
rect 27764 20216 28080 20244
rect 27764 20204 27770 20216
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 552 20154 31648 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 12096 20154
rect 12148 20102 12160 20154
rect 12212 20102 12224 20154
rect 12276 20102 12288 20154
rect 12340 20102 12352 20154
rect 12404 20102 19870 20154
rect 19922 20102 19934 20154
rect 19986 20102 19998 20154
rect 20050 20102 20062 20154
rect 20114 20102 20126 20154
rect 20178 20102 27644 20154
rect 27696 20102 27708 20154
rect 27760 20102 27772 20154
rect 27824 20102 27836 20154
rect 27888 20102 27900 20154
rect 27952 20102 31648 20154
rect 552 20080 31648 20102
rect 14826 20000 14832 20052
rect 14884 20040 14890 20052
rect 18230 20040 18236 20052
rect 14884 20012 18236 20040
rect 14884 20000 14890 20012
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 19061 20043 19119 20049
rect 19061 20040 19073 20043
rect 18564 20012 19073 20040
rect 18564 20000 18570 20012
rect 19061 20009 19073 20012
rect 19107 20040 19119 20043
rect 19242 20040 19248 20052
rect 19107 20012 19248 20040
rect 19107 20009 19119 20012
rect 19061 20003 19119 20009
rect 19242 20000 19248 20012
rect 19300 20000 19306 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22152 20012 26188 20040
rect 22152 20000 22158 20012
rect 16482 19972 16488 19984
rect 14936 19944 16488 19972
rect 14826 19864 14832 19916
rect 14884 19864 14890 19916
rect 14936 19913 14964 19944
rect 16482 19932 16488 19944
rect 16540 19932 16546 19984
rect 18322 19972 18328 19984
rect 17696 19944 18328 19972
rect 14921 19907 14979 19913
rect 14921 19873 14933 19907
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 15013 19907 15071 19913
rect 15013 19873 15025 19907
rect 15059 19873 15071 19907
rect 15013 19867 15071 19873
rect 15197 19907 15255 19913
rect 15197 19873 15209 19907
rect 15243 19904 15255 19907
rect 15378 19904 15384 19916
rect 15243 19876 15384 19904
rect 15243 19873 15255 19876
rect 15197 19867 15255 19873
rect 15028 19836 15056 19867
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 17696 19913 17724 19944
rect 18322 19932 18328 19944
rect 18380 19932 18386 19984
rect 19420 19975 19478 19981
rect 19420 19941 19432 19975
rect 19466 19972 19478 19975
rect 19610 19972 19616 19984
rect 19466 19944 19616 19972
rect 19466 19941 19478 19944
rect 19420 19935 19478 19941
rect 19610 19932 19616 19944
rect 19668 19932 19674 19984
rect 20254 19932 20260 19984
rect 20312 19972 20318 19984
rect 21545 19975 21603 19981
rect 20312 19944 21496 19972
rect 20312 19932 20318 19944
rect 17954 19913 17960 19916
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 17948 19867 17960 19913
rect 17954 19864 17960 19867
rect 18012 19864 18018 19916
rect 19150 19864 19156 19916
rect 19208 19864 19214 19916
rect 21468 19913 21496 19944
rect 21545 19941 21557 19975
rect 21591 19972 21603 19975
rect 22002 19972 22008 19984
rect 21591 19944 22008 19972
rect 21591 19941 21603 19944
rect 21545 19935 21603 19941
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 23109 19975 23167 19981
rect 23109 19941 23121 19975
rect 23155 19972 23167 19975
rect 23382 19972 23388 19984
rect 23155 19944 23388 19972
rect 23155 19941 23167 19944
rect 23109 19935 23167 19941
rect 23382 19932 23388 19944
rect 23440 19972 23446 19984
rect 25314 19972 25320 19984
rect 23440 19944 25320 19972
rect 23440 19932 23446 19944
rect 25314 19932 25320 19944
rect 25372 19932 25378 19984
rect 26160 19981 26188 20012
rect 26234 20000 26240 20052
rect 26292 20040 26298 20052
rect 26292 20012 27016 20040
rect 26292 20000 26298 20012
rect 26145 19975 26203 19981
rect 25700 19944 26004 19972
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 21269 19907 21327 19913
rect 21269 19904 21281 19907
rect 20855 19876 21281 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 21269 19873 21281 19876
rect 21315 19873 21327 19907
rect 21269 19867 21327 19873
rect 21453 19907 21511 19913
rect 21453 19873 21465 19907
rect 21499 19873 21511 19907
rect 21453 19867 21511 19873
rect 21634 19864 21640 19916
rect 21692 19864 21698 19916
rect 21726 19864 21732 19916
rect 21784 19913 21790 19916
rect 21784 19907 21813 19913
rect 21801 19873 21813 19907
rect 21784 19867 21813 19873
rect 21913 19907 21971 19913
rect 21913 19873 21925 19907
rect 21959 19904 21971 19907
rect 23658 19904 23664 19916
rect 21959 19876 23664 19904
rect 21959 19873 21971 19876
rect 21913 19867 21971 19873
rect 21784 19864 21790 19867
rect 15838 19836 15844 19848
rect 15028 19808 15844 19836
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 20993 19839 21051 19845
rect 20993 19836 21005 19839
rect 20180 19808 21005 19836
rect 14553 19703 14611 19709
rect 14553 19669 14565 19703
rect 14599 19700 14611 19703
rect 14642 19700 14648 19712
rect 14599 19672 14648 19700
rect 14599 19669 14611 19672
rect 14553 19663 14611 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 19794 19660 19800 19712
rect 19852 19700 19858 19712
rect 20180 19700 20208 19808
rect 20993 19805 21005 19808
rect 21039 19805 21051 19839
rect 20993 19799 21051 19805
rect 21082 19796 21088 19848
rect 21140 19836 21146 19848
rect 21928 19836 21956 19867
rect 23658 19864 23664 19876
rect 23716 19864 23722 19916
rect 23845 19907 23903 19913
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24118 19904 24124 19916
rect 23891 19876 24124 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24118 19864 24124 19876
rect 24176 19904 24182 19916
rect 24302 19904 24308 19916
rect 24176 19876 24308 19904
rect 24176 19864 24182 19876
rect 24302 19864 24308 19876
rect 24360 19864 24366 19916
rect 24946 19864 24952 19916
rect 25004 19864 25010 19916
rect 25700 19904 25728 19944
rect 25332 19876 25728 19904
rect 21140 19808 21956 19836
rect 21140 19796 21146 19808
rect 22278 19796 22284 19848
rect 22336 19796 22342 19848
rect 23750 19796 23756 19848
rect 23808 19796 23814 19848
rect 24210 19796 24216 19848
rect 24268 19796 24274 19848
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19805 24915 19839
rect 24857 19799 24915 19805
rect 20530 19728 20536 19780
rect 20588 19768 20594 19780
rect 24872 19768 24900 19799
rect 25332 19777 25360 19876
rect 25774 19864 25780 19916
rect 25832 19864 25838 19916
rect 25869 19907 25927 19913
rect 25869 19873 25881 19907
rect 25915 19873 25927 19907
rect 25976 19904 26004 19944
rect 26145 19941 26157 19975
rect 26191 19972 26203 19975
rect 26988 19972 27016 20012
rect 28902 19972 28908 19984
rect 26191 19944 26832 19972
rect 26191 19941 26203 19944
rect 26145 19935 26203 19941
rect 26421 19907 26479 19913
rect 26421 19904 26433 19907
rect 25976 19876 26433 19904
rect 25869 19867 25927 19873
rect 26421 19873 26433 19876
rect 26467 19873 26479 19907
rect 26421 19867 26479 19873
rect 25682 19796 25688 19848
rect 25740 19836 25746 19848
rect 25884 19836 25912 19867
rect 26602 19864 26608 19916
rect 26660 19864 26666 19916
rect 26804 19913 26832 19944
rect 26988 19944 28908 19972
rect 26988 19913 27016 19944
rect 28902 19932 28908 19944
rect 28960 19932 28966 19984
rect 26789 19907 26847 19913
rect 26789 19873 26801 19907
rect 26835 19873 26847 19907
rect 26789 19867 26847 19873
rect 26973 19907 27031 19913
rect 26973 19873 26985 19907
rect 27019 19873 27031 19907
rect 26973 19867 27031 19873
rect 27617 19907 27675 19913
rect 27617 19873 27629 19907
rect 27663 19904 27675 19907
rect 28166 19904 28172 19916
rect 27663 19876 28172 19904
rect 27663 19873 27675 19876
rect 27617 19867 27675 19873
rect 28166 19864 28172 19876
rect 28224 19864 28230 19916
rect 25740 19808 25912 19836
rect 25740 19796 25746 19808
rect 26234 19796 26240 19848
rect 26292 19796 26298 19848
rect 26697 19839 26755 19845
rect 26697 19836 26709 19839
rect 26528 19808 26709 19836
rect 20588 19740 24900 19768
rect 25317 19771 25375 19777
rect 20588 19728 20594 19740
rect 25317 19737 25329 19771
rect 25363 19737 25375 19771
rect 25317 19731 25375 19737
rect 19852 19672 20208 19700
rect 19852 19660 19858 19672
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 25593 19703 25651 19709
rect 25593 19669 25605 19703
rect 25639 19700 25651 19703
rect 25866 19700 25872 19712
rect 25639 19672 25872 19700
rect 25639 19669 25651 19672
rect 25593 19663 25651 19669
rect 25866 19660 25872 19672
rect 25924 19660 25930 19712
rect 26050 19660 26056 19712
rect 26108 19700 26114 19712
rect 26528 19700 26556 19808
rect 26697 19805 26709 19808
rect 26743 19805 26755 19839
rect 26697 19799 26755 19805
rect 27430 19796 27436 19848
rect 27488 19836 27494 19848
rect 27525 19839 27583 19845
rect 27525 19836 27537 19839
rect 27488 19808 27537 19836
rect 27488 19796 27494 19808
rect 27525 19805 27537 19808
rect 27571 19805 27583 19839
rect 27525 19799 27583 19805
rect 26108 19672 26556 19700
rect 26108 19660 26114 19672
rect 26694 19660 26700 19712
rect 26752 19700 26758 19712
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 26752 19672 27169 19700
rect 26752 19660 26758 19672
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 27157 19663 27215 19669
rect 27249 19703 27307 19709
rect 27249 19669 27261 19703
rect 27295 19700 27307 19703
rect 27338 19700 27344 19712
rect 27295 19672 27344 19700
rect 27295 19669 27307 19672
rect 27249 19663 27307 19669
rect 27338 19660 27344 19672
rect 27396 19660 27402 19712
rect 552 19610 31648 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 11436 19610
rect 11488 19558 11500 19610
rect 11552 19558 11564 19610
rect 11616 19558 11628 19610
rect 11680 19558 11692 19610
rect 11744 19558 19210 19610
rect 19262 19558 19274 19610
rect 19326 19558 19338 19610
rect 19390 19558 19402 19610
rect 19454 19558 19466 19610
rect 19518 19558 26984 19610
rect 27036 19558 27048 19610
rect 27100 19558 27112 19610
rect 27164 19558 27176 19610
rect 27228 19558 27240 19610
rect 27292 19558 31648 19610
rect 552 19536 31648 19558
rect 19245 19499 19303 19505
rect 19245 19465 19257 19499
rect 19291 19496 19303 19499
rect 19610 19496 19616 19508
rect 19291 19468 19616 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 21082 19496 21088 19508
rect 19720 19468 21088 19496
rect 16574 19428 16580 19440
rect 16224 19400 16580 19428
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 14642 19301 14648 19304
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13872 19264 14105 19292
rect 13872 19252 13878 19264
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 14231 19264 14381 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 14369 19261 14381 19264
rect 14415 19261 14427 19295
rect 14636 19292 14648 19301
rect 14603 19264 14648 19292
rect 14369 19255 14427 19261
rect 14636 19255 14648 19264
rect 14642 19252 14648 19255
rect 14700 19252 14706 19304
rect 15838 19252 15844 19304
rect 15896 19252 15902 19304
rect 16224 19301 16252 19400
rect 16574 19388 16580 19400
rect 16632 19388 16638 19440
rect 17402 19388 17408 19440
rect 17460 19428 17466 19440
rect 19720 19428 19748 19468
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 21729 19499 21787 19505
rect 21729 19465 21741 19499
rect 21775 19496 21787 19499
rect 22002 19496 22008 19508
rect 21775 19468 22008 19496
rect 21775 19465 21787 19468
rect 21729 19459 21787 19465
rect 22002 19456 22008 19468
rect 22060 19456 22066 19508
rect 22554 19456 22560 19508
rect 22612 19496 22618 19508
rect 23201 19499 23259 19505
rect 23201 19496 23213 19499
rect 22612 19468 23213 19496
rect 22612 19456 22618 19468
rect 23201 19465 23213 19468
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 26421 19499 26479 19505
rect 26421 19465 26433 19499
rect 26467 19496 26479 19499
rect 26510 19496 26516 19508
rect 26467 19468 26516 19496
rect 26467 19465 26479 19468
rect 26421 19459 26479 19465
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 28261 19499 28319 19505
rect 28261 19496 28273 19499
rect 28132 19468 28273 19496
rect 28132 19456 28138 19468
rect 28261 19465 28273 19468
rect 28307 19465 28319 19499
rect 28261 19459 28319 19465
rect 17460 19400 19748 19428
rect 17460 19388 17466 19400
rect 16209 19295 16267 19301
rect 16209 19292 16221 19295
rect 15948 19264 16221 19292
rect 15194 19184 15200 19236
rect 15252 19224 15258 19236
rect 15948 19224 15976 19264
rect 16209 19261 16221 19264
rect 16255 19261 16267 19295
rect 16209 19255 16267 19261
rect 16482 19252 16488 19304
rect 16540 19294 16546 19304
rect 16540 19266 16712 19294
rect 16540 19264 16574 19266
rect 16540 19252 16546 19264
rect 15252 19196 15976 19224
rect 16025 19227 16083 19233
rect 15252 19184 15258 19196
rect 16025 19193 16037 19227
rect 16071 19193 16083 19227
rect 16684 19224 16712 19266
rect 16758 19252 16764 19304
rect 16816 19252 16822 19304
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 16868 19224 16896 19255
rect 16942 19252 16948 19304
rect 17000 19252 17006 19304
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19261 17187 19295
rect 17129 19255 17187 19261
rect 16684 19196 16896 19224
rect 17144 19224 17172 19255
rect 17218 19252 17224 19304
rect 17276 19252 17282 19304
rect 17788 19292 17816 19400
rect 25222 19388 25228 19440
rect 25280 19428 25286 19440
rect 27430 19428 27436 19440
rect 25280 19400 27436 19428
rect 25280 19388 25286 19400
rect 27430 19388 27436 19400
rect 27488 19388 27494 19440
rect 19702 19360 19708 19372
rect 19444 19332 19708 19360
rect 17865 19295 17923 19301
rect 17865 19292 17877 19295
rect 17788 19264 17877 19292
rect 17865 19261 17877 19264
rect 17911 19261 17923 19295
rect 17865 19255 17923 19261
rect 17957 19295 18015 19301
rect 17957 19261 17969 19295
rect 18003 19261 18015 19295
rect 17957 19255 18015 19261
rect 17770 19224 17776 19236
rect 17144 19196 17776 19224
rect 16025 19187 16083 19193
rect 15654 19116 15660 19168
rect 15712 19156 15718 19168
rect 15749 19159 15807 19165
rect 15749 19156 15761 19159
rect 15712 19128 15761 19156
rect 15712 19116 15718 19128
rect 15749 19125 15761 19128
rect 15795 19156 15807 19159
rect 16040 19156 16068 19187
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 17972 19224 18000 19255
rect 18046 19252 18052 19304
rect 18104 19252 18110 19304
rect 19444 19301 19472 19332
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 20272 19332 20484 19360
rect 18233 19295 18291 19301
rect 18233 19261 18245 19295
rect 18279 19292 18291 19295
rect 19429 19295 19487 19301
rect 18279 19264 19380 19292
rect 18279 19261 18291 19264
rect 18233 19255 18291 19261
rect 17972 19196 18276 19224
rect 18248 19168 18276 19196
rect 15795 19128 16068 19156
rect 15795 19125 15807 19128
rect 15749 19119 15807 19125
rect 16482 19116 16488 19168
rect 16540 19116 16546 19168
rect 16574 19116 16580 19168
rect 16632 19156 16638 19168
rect 17313 19159 17371 19165
rect 17313 19156 17325 19159
rect 16632 19128 17325 19156
rect 16632 19116 16638 19128
rect 17313 19125 17325 19128
rect 17359 19125 17371 19159
rect 17313 19119 17371 19125
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19156 17647 19159
rect 17954 19156 17960 19168
rect 17635 19128 17960 19156
rect 17635 19125 17647 19128
rect 17589 19119 17647 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 18230 19116 18236 19168
rect 18288 19116 18294 19168
rect 19352 19156 19380 19264
rect 19429 19261 19441 19295
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19292 19671 19295
rect 19794 19292 19800 19304
rect 19659 19264 19800 19292
rect 19659 19261 19671 19264
rect 19613 19255 19671 19261
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 20272 19301 20300 19332
rect 20257 19295 20315 19301
rect 20257 19292 20269 19295
rect 20235 19264 20269 19292
rect 20257 19261 20269 19264
rect 20303 19261 20315 19295
rect 20257 19255 20315 19261
rect 20349 19295 20407 19301
rect 20349 19261 20361 19295
rect 20395 19261 20407 19295
rect 20456 19292 20484 19332
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 26694 19320 26700 19372
rect 26752 19320 26758 19372
rect 21450 19292 21456 19304
rect 20456 19264 21456 19292
rect 20349 19255 20407 19261
rect 20165 19227 20223 19233
rect 20165 19193 20177 19227
rect 20211 19224 20223 19227
rect 20364 19224 20392 19255
rect 21450 19252 21456 19264
rect 21508 19252 21514 19304
rect 21542 19252 21548 19304
rect 21600 19292 21606 19304
rect 21821 19295 21879 19301
rect 21821 19292 21833 19295
rect 21600 19264 21833 19292
rect 21600 19252 21606 19264
rect 21821 19261 21833 19264
rect 21867 19261 21879 19295
rect 21821 19255 21879 19261
rect 23477 19295 23535 19301
rect 23477 19261 23489 19295
rect 23523 19292 23535 19295
rect 23566 19292 23572 19304
rect 23523 19264 23572 19292
rect 23523 19261 23535 19264
rect 23477 19255 23535 19261
rect 23566 19252 23572 19264
rect 23624 19252 23630 19304
rect 23845 19295 23903 19301
rect 23845 19261 23857 19295
rect 23891 19292 23903 19295
rect 24394 19292 24400 19304
rect 23891 19264 24400 19292
rect 23891 19261 23903 19264
rect 23845 19255 23903 19261
rect 24394 19252 24400 19264
rect 24452 19252 24458 19304
rect 25314 19252 25320 19304
rect 25372 19252 25378 19304
rect 26326 19252 26332 19304
rect 26384 19252 26390 19304
rect 26970 19252 26976 19304
rect 27028 19252 27034 19304
rect 27157 19295 27215 19301
rect 27157 19261 27169 19295
rect 27203 19292 27215 19295
rect 27338 19292 27344 19304
rect 27203 19264 27344 19292
rect 27203 19261 27215 19264
rect 27157 19255 27215 19261
rect 27338 19252 27344 19264
rect 27396 19252 27402 19304
rect 27982 19252 27988 19304
rect 28040 19292 28046 19304
rect 28534 19292 28540 19304
rect 28040 19264 28540 19292
rect 28040 19252 28046 19264
rect 20622 19233 20628 19236
rect 20616 19224 20628 19233
rect 20211 19196 20392 19224
rect 20583 19196 20628 19224
rect 20211 19193 20223 19196
rect 20165 19187 20223 19193
rect 20616 19187 20628 19196
rect 20622 19184 20628 19187
rect 20680 19184 20686 19236
rect 22094 19233 22100 19236
rect 22088 19187 22100 19233
rect 22094 19184 22100 19187
rect 22152 19184 22158 19236
rect 23661 19227 23719 19233
rect 23661 19193 23673 19227
rect 23707 19224 23719 19227
rect 24090 19227 24148 19233
rect 24090 19224 24102 19227
rect 23707 19196 24102 19224
rect 23707 19193 23719 19196
rect 23661 19187 23719 19193
rect 24090 19193 24102 19196
rect 24136 19193 24148 19227
rect 24090 19187 24148 19193
rect 24486 19184 24492 19236
rect 24544 19224 24550 19236
rect 26053 19227 26111 19233
rect 26053 19224 26065 19227
rect 24544 19196 26065 19224
rect 24544 19184 24550 19196
rect 26053 19193 26065 19196
rect 26099 19193 26111 19227
rect 26053 19187 26111 19193
rect 26142 19184 26148 19236
rect 26200 19224 26206 19236
rect 28092 19233 28120 19264
rect 28534 19252 28540 19264
rect 28592 19252 28598 19304
rect 26421 19227 26479 19233
rect 26421 19224 26433 19227
rect 26200 19196 26433 19224
rect 26200 19184 26206 19196
rect 26421 19193 26433 19196
rect 26467 19193 26479 19227
rect 27065 19227 27123 19233
rect 27065 19224 27077 19227
rect 26421 19187 26479 19193
rect 26528 19196 27077 19224
rect 22370 19156 22376 19168
rect 19352 19128 22376 19156
rect 22370 19116 22376 19128
rect 22428 19156 22434 19168
rect 23290 19156 23296 19168
rect 22428 19128 23296 19156
rect 22428 19116 22434 19128
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 26528 19165 26556 19196
rect 27065 19193 27077 19196
rect 27111 19193 27123 19227
rect 27065 19187 27123 19193
rect 28077 19227 28135 19233
rect 28077 19193 28089 19227
rect 28123 19193 28135 19227
rect 28077 19187 28135 19193
rect 28258 19184 28264 19236
rect 28316 19233 28322 19236
rect 28316 19227 28335 19233
rect 28323 19193 28335 19227
rect 28316 19187 28335 19193
rect 28316 19184 28322 19187
rect 26513 19159 26571 19165
rect 26513 19125 26525 19159
rect 26559 19125 26571 19159
rect 26513 19119 26571 19125
rect 28442 19116 28448 19168
rect 28500 19116 28506 19168
rect 28626 19116 28632 19168
rect 28684 19156 28690 19168
rect 29362 19156 29368 19168
rect 28684 19128 29368 19156
rect 28684 19116 28690 19128
rect 29362 19116 29368 19128
rect 29420 19116 29426 19168
rect 552 19066 31648 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 12096 19066
rect 12148 19014 12160 19066
rect 12212 19014 12224 19066
rect 12276 19014 12288 19066
rect 12340 19014 12352 19066
rect 12404 19014 19870 19066
rect 19922 19014 19934 19066
rect 19986 19014 19998 19066
rect 20050 19014 20062 19066
rect 20114 19014 20126 19066
rect 20178 19014 27644 19066
rect 27696 19014 27708 19066
rect 27760 19014 27772 19066
rect 27824 19014 27836 19066
rect 27888 19014 27900 19066
rect 27952 19014 31648 19066
rect 552 18992 31648 19014
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 16540 18912 16574 18952
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 21266 18952 21272 18964
rect 16908 18924 21272 18952
rect 16908 18912 16914 18924
rect 21266 18912 21272 18924
rect 21324 18912 21330 18964
rect 21542 18912 21548 18964
rect 21600 18912 21606 18964
rect 22094 18912 22100 18964
rect 22152 18912 22158 18964
rect 23566 18912 23572 18964
rect 23624 18912 23630 18964
rect 23934 18952 23940 18964
rect 23768 18924 23940 18952
rect 16546 18884 16574 18912
rect 16730 18887 16788 18893
rect 16730 18884 16742 18887
rect 16546 18856 16742 18884
rect 16730 18853 16742 18856
rect 16776 18853 16788 18887
rect 16730 18847 16788 18853
rect 17862 18844 17868 18896
rect 17920 18884 17926 18896
rect 18049 18887 18107 18893
rect 18049 18884 18061 18887
rect 17920 18856 18061 18884
rect 17920 18844 17926 18856
rect 18049 18853 18061 18856
rect 18095 18853 18107 18887
rect 22278 18884 22284 18896
rect 18049 18847 18107 18853
rect 21560 18856 22284 18884
rect 21560 18828 21588 18856
rect 22278 18844 22284 18856
rect 22336 18884 22342 18896
rect 22336 18856 22416 18884
rect 22336 18844 22342 18856
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15565 18819 15623 18825
rect 15565 18816 15577 18819
rect 15252 18788 15577 18816
rect 15252 18776 15258 18788
rect 15565 18785 15577 18788
rect 15611 18785 15623 18819
rect 15565 18779 15623 18785
rect 15749 18819 15807 18825
rect 15749 18785 15761 18819
rect 15795 18816 15807 18819
rect 16298 18816 16304 18828
rect 15795 18788 16304 18816
rect 15795 18785 15807 18788
rect 15749 18779 15807 18785
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 16574 18816 16580 18828
rect 16531 18788 16580 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 19613 18819 19671 18825
rect 19613 18816 19625 18819
rect 18892 18788 19625 18816
rect 18892 18760 18920 18788
rect 19613 18785 19625 18788
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 21453 18817 21511 18823
rect 21453 18783 21465 18817
rect 21499 18816 21511 18817
rect 21542 18816 21548 18828
rect 21499 18788 21548 18816
rect 21499 18783 21511 18788
rect 21453 18777 21511 18783
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 21913 18819 21971 18825
rect 21913 18785 21925 18819
rect 21959 18816 21971 18819
rect 22186 18816 22192 18828
rect 21959 18788 22192 18816
rect 21959 18785 21971 18788
rect 21913 18779 21971 18785
rect 22186 18776 22192 18788
rect 22244 18776 22250 18828
rect 22388 18825 22416 18856
rect 22373 18819 22431 18825
rect 22373 18785 22385 18819
rect 22419 18785 22431 18819
rect 22373 18779 22431 18785
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 23658 18816 23664 18828
rect 23072 18788 23664 18816
rect 23072 18776 23078 18788
rect 23658 18776 23664 18788
rect 23716 18816 23722 18828
rect 23768 18825 23796 18924
rect 23934 18912 23940 18924
rect 23992 18912 23998 18964
rect 24394 18912 24400 18964
rect 24452 18912 24458 18964
rect 25869 18955 25927 18961
rect 25869 18921 25881 18955
rect 25915 18952 25927 18955
rect 26050 18952 26056 18964
rect 25915 18924 26056 18952
rect 25915 18921 25927 18924
rect 25869 18915 25927 18921
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 27801 18955 27859 18961
rect 27801 18952 27813 18955
rect 27172 18924 27813 18952
rect 23845 18887 23903 18893
rect 23845 18853 23857 18887
rect 23891 18884 23903 18887
rect 25222 18884 25228 18896
rect 23891 18856 25228 18884
rect 23891 18853 23903 18856
rect 23845 18847 23903 18853
rect 25222 18844 25228 18856
rect 25280 18844 25286 18896
rect 23753 18819 23811 18825
rect 23753 18816 23765 18819
rect 23716 18788 23765 18816
rect 23716 18776 23722 18788
rect 23753 18785 23765 18788
rect 23799 18785 23811 18819
rect 23937 18819 23995 18825
rect 23937 18816 23949 18819
rect 23753 18779 23811 18785
rect 23860 18788 23949 18816
rect 18874 18708 18880 18760
rect 18932 18708 18938 18760
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18748 21787 18751
rect 23290 18748 23296 18760
rect 21775 18720 23296 18748
rect 21775 18717 21787 18720
rect 21729 18711 21787 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 17770 18640 17776 18692
rect 17828 18680 17834 18692
rect 19794 18680 19800 18692
rect 17828 18652 19800 18680
rect 17828 18640 17834 18652
rect 19794 18640 19800 18652
rect 19852 18640 19858 18692
rect 21634 18640 21640 18692
rect 21692 18680 21698 18692
rect 23860 18680 23888 18788
rect 23937 18785 23949 18788
rect 23983 18785 23995 18819
rect 23937 18779 23995 18785
rect 24026 18776 24032 18828
rect 24084 18825 24090 18828
rect 24084 18819 24113 18825
rect 24101 18816 24113 18819
rect 24101 18788 24440 18816
rect 24101 18785 24113 18788
rect 24084 18779 24113 18785
rect 24084 18776 24090 18779
rect 24213 18751 24271 18757
rect 24213 18748 24225 18751
rect 23952 18720 24225 18748
rect 23952 18692 23980 18720
rect 24213 18717 24225 18720
rect 24259 18717 24271 18751
rect 24412 18748 24440 18788
rect 24486 18776 24492 18828
rect 24544 18816 24550 18828
rect 25041 18819 25099 18825
rect 25041 18816 25053 18819
rect 24544 18788 25053 18816
rect 24544 18776 24550 18788
rect 25041 18785 25053 18788
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 25130 18776 25136 18828
rect 25188 18816 25194 18828
rect 25961 18819 26019 18825
rect 25961 18816 25973 18819
rect 25188 18788 25973 18816
rect 25188 18776 25194 18788
rect 25961 18785 25973 18788
rect 26007 18785 26019 18819
rect 25961 18779 26019 18785
rect 26605 18819 26663 18825
rect 26605 18785 26617 18819
rect 26651 18816 26663 18819
rect 26878 18816 26884 18828
rect 26651 18788 26884 18816
rect 26651 18785 26663 18788
rect 26605 18779 26663 18785
rect 26878 18776 26884 18788
rect 26936 18776 26942 18828
rect 27172 18825 27200 18924
rect 27801 18921 27813 18924
rect 27847 18952 27859 18955
rect 27847 18924 29684 18952
rect 27847 18921 27859 18924
rect 27801 18915 27859 18921
rect 27433 18887 27491 18893
rect 27433 18884 27445 18887
rect 27356 18856 27445 18884
rect 27356 18825 27384 18856
rect 27433 18853 27445 18856
rect 27479 18853 27491 18887
rect 28261 18887 28319 18893
rect 28261 18884 28273 18887
rect 27433 18847 27491 18853
rect 27724 18856 28273 18884
rect 27724 18825 27752 18856
rect 28261 18853 28273 18856
rect 28307 18853 28319 18887
rect 28261 18847 28319 18853
rect 28534 18844 28540 18896
rect 28592 18884 28598 18896
rect 28592 18856 29132 18884
rect 28592 18844 28598 18856
rect 27157 18819 27215 18825
rect 27157 18785 27169 18819
rect 27203 18785 27215 18819
rect 27157 18779 27215 18785
rect 27341 18819 27399 18825
rect 27341 18785 27353 18819
rect 27387 18785 27399 18819
rect 27341 18779 27399 18785
rect 27709 18819 27767 18825
rect 27709 18785 27721 18819
rect 27755 18785 27767 18819
rect 27709 18779 27767 18785
rect 27985 18819 28043 18825
rect 27985 18785 27997 18819
rect 28031 18816 28043 18819
rect 28031 18788 28304 18816
rect 28031 18785 28043 18788
rect 27985 18779 28043 18785
rect 24762 18748 24768 18760
rect 24412 18720 24768 18748
rect 24213 18711 24271 18717
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 26510 18708 26516 18760
rect 26568 18708 26574 18760
rect 26970 18708 26976 18760
rect 27028 18708 27034 18760
rect 27430 18708 27436 18760
rect 27488 18748 27494 18760
rect 27617 18751 27675 18757
rect 27488 18720 27568 18748
rect 27488 18708 27494 18720
rect 21692 18652 23888 18680
rect 21692 18640 21698 18652
rect 15838 18572 15844 18624
rect 15896 18612 15902 18624
rect 15933 18615 15991 18621
rect 15933 18612 15945 18615
rect 15896 18584 15945 18612
rect 15896 18572 15902 18584
rect 15933 18581 15945 18584
rect 15979 18581 15991 18615
rect 15933 18575 15991 18581
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 17865 18615 17923 18621
rect 17865 18612 17877 18615
rect 17552 18584 17877 18612
rect 17552 18572 17558 18584
rect 17865 18581 17877 18584
rect 17911 18581 17923 18615
rect 17865 18575 17923 18581
rect 19521 18615 19579 18621
rect 19521 18581 19533 18615
rect 19567 18612 19579 18615
rect 19610 18612 19616 18624
rect 19567 18584 19616 18612
rect 19567 18581 19579 18584
rect 19521 18575 19579 18581
rect 19610 18572 19616 18584
rect 19668 18572 19674 18624
rect 23860 18612 23888 18652
rect 23934 18640 23940 18692
rect 23992 18640 23998 18692
rect 24026 18612 24032 18624
rect 23860 18584 24032 18612
rect 24026 18572 24032 18584
rect 24084 18612 24090 18624
rect 24854 18612 24860 18624
rect 24084 18584 24860 18612
rect 24084 18572 24090 18584
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 27341 18615 27399 18621
rect 27341 18581 27353 18615
rect 27387 18612 27399 18615
rect 27430 18612 27436 18624
rect 27387 18584 27436 18612
rect 27387 18581 27399 18584
rect 27341 18575 27399 18581
rect 27430 18572 27436 18584
rect 27488 18572 27494 18624
rect 27540 18612 27568 18720
rect 27617 18717 27629 18751
rect 27663 18748 27675 18751
rect 28000 18748 28028 18779
rect 28276 18760 28304 18788
rect 28442 18776 28448 18828
rect 28500 18816 28506 18828
rect 28997 18819 29055 18825
rect 28997 18816 29009 18819
rect 28500 18788 29009 18816
rect 28500 18776 28506 18788
rect 28997 18785 29009 18788
rect 29043 18785 29055 18819
rect 29104 18816 29132 18856
rect 29362 18844 29368 18896
rect 29420 18844 29426 18896
rect 29656 18893 29684 18924
rect 29641 18887 29699 18893
rect 29641 18853 29653 18887
rect 29687 18853 29699 18887
rect 29641 18847 29699 18853
rect 29825 18819 29883 18825
rect 29825 18816 29837 18819
rect 29104 18788 29837 18816
rect 28997 18779 29055 18785
rect 29825 18785 29837 18788
rect 29871 18816 29883 18819
rect 30374 18816 30380 18828
rect 29871 18788 30380 18816
rect 29871 18785 29883 18788
rect 29825 18779 29883 18785
rect 30374 18776 30380 18788
rect 30432 18776 30438 18828
rect 27663 18720 28028 18748
rect 27663 18717 27675 18720
rect 27617 18711 27675 18717
rect 28074 18708 28080 18760
rect 28132 18748 28138 18760
rect 28169 18751 28227 18757
rect 28169 18748 28181 18751
rect 28132 18720 28181 18748
rect 28132 18708 28138 18720
rect 28169 18717 28181 18720
rect 28215 18717 28227 18751
rect 28169 18711 28227 18717
rect 28184 18680 28212 18711
rect 28258 18708 28264 18760
rect 28316 18708 28322 18760
rect 28813 18751 28871 18757
rect 28813 18717 28825 18751
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 28718 18680 28724 18692
rect 28184 18652 28724 18680
rect 28718 18640 28724 18652
rect 28776 18680 28782 18692
rect 28828 18680 28856 18711
rect 30009 18683 30067 18689
rect 30009 18680 30021 18683
rect 28776 18652 28856 18680
rect 29380 18652 30021 18680
rect 28776 18640 28782 18652
rect 28626 18612 28632 18624
rect 27540 18584 28632 18612
rect 28626 18572 28632 18584
rect 28684 18572 28690 18624
rect 29380 18621 29408 18652
rect 30009 18649 30021 18652
rect 30055 18649 30067 18683
rect 30009 18643 30067 18649
rect 29365 18615 29423 18621
rect 29365 18581 29377 18615
rect 29411 18581 29423 18615
rect 29365 18575 29423 18581
rect 29546 18572 29552 18624
rect 29604 18572 29610 18624
rect 552 18522 31648 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 11436 18522
rect 11488 18470 11500 18522
rect 11552 18470 11564 18522
rect 11616 18470 11628 18522
rect 11680 18470 11692 18522
rect 11744 18470 19210 18522
rect 19262 18470 19274 18522
rect 19326 18470 19338 18522
rect 19390 18470 19402 18522
rect 19454 18470 19466 18522
rect 19518 18470 26984 18522
rect 27036 18470 27048 18522
rect 27100 18470 27112 18522
rect 27164 18470 27176 18522
rect 27228 18470 27240 18522
rect 27292 18470 31648 18522
rect 552 18448 31648 18470
rect 16298 18368 16304 18420
rect 16356 18408 16362 18420
rect 16761 18411 16819 18417
rect 16761 18408 16773 18411
rect 16356 18380 16773 18408
rect 16356 18368 16362 18380
rect 16761 18377 16773 18380
rect 16807 18377 16819 18411
rect 16761 18371 16819 18377
rect 26050 18368 26056 18420
rect 26108 18408 26114 18420
rect 27982 18408 27988 18420
rect 26108 18380 27988 18408
rect 26108 18368 26114 18380
rect 27982 18368 27988 18380
rect 28040 18368 28046 18420
rect 30374 18368 30380 18420
rect 30432 18368 30438 18420
rect 18966 18272 18972 18284
rect 18156 18244 18972 18272
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14553 18207 14611 18213
rect 14553 18204 14565 18207
rect 13872 18176 14565 18204
rect 13872 18164 13878 18176
rect 14553 18173 14565 18176
rect 14599 18173 14611 18207
rect 14553 18167 14611 18173
rect 14645 18207 14703 18213
rect 14645 18173 14657 18207
rect 14691 18204 14703 18207
rect 15381 18207 15439 18213
rect 15381 18204 15393 18207
rect 14691 18176 15393 18204
rect 14691 18173 14703 18176
rect 14645 18167 14703 18173
rect 15381 18173 15393 18176
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 17773 18207 17831 18213
rect 17773 18173 17785 18207
rect 17819 18204 17831 18207
rect 17862 18204 17868 18216
rect 17819 18176 17868 18204
rect 17819 18173 17831 18176
rect 17773 18167 17831 18173
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 18156 18213 18184 18244
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20530 18272 20536 18284
rect 20312 18244 20536 18272
rect 20312 18232 20318 18244
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18173 18199 18207
rect 18141 18167 18199 18173
rect 18230 18164 18236 18216
rect 18288 18164 18294 18216
rect 18322 18164 18328 18216
rect 18380 18164 18386 18216
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 15013 18139 15071 18145
rect 15013 18105 15025 18139
rect 15059 18105 15071 18139
rect 15013 18099 15071 18105
rect 14826 18028 14832 18080
rect 14884 18028 14890 18080
rect 15028 18068 15056 18099
rect 15194 18096 15200 18148
rect 15252 18096 15258 18148
rect 15470 18096 15476 18148
rect 15528 18136 15534 18148
rect 15626 18139 15684 18145
rect 15626 18136 15638 18139
rect 15528 18108 15638 18136
rect 15528 18096 15534 18108
rect 15626 18105 15638 18108
rect 15672 18105 15684 18139
rect 15626 18099 15684 18105
rect 16574 18096 16580 18148
rect 16632 18136 16638 18148
rect 16945 18139 17003 18145
rect 16945 18136 16957 18139
rect 16632 18108 16957 18136
rect 16632 18096 16638 18108
rect 16945 18105 16957 18108
rect 16991 18136 17003 18139
rect 17218 18136 17224 18148
rect 16991 18108 17224 18136
rect 16991 18105 17003 18108
rect 16945 18099 17003 18105
rect 17218 18096 17224 18108
rect 17276 18096 17282 18148
rect 18248 18136 18276 18164
rect 17788 18108 18276 18136
rect 18524 18136 18552 18167
rect 18874 18164 18880 18216
rect 18932 18164 18938 18216
rect 20364 18213 20392 18244
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 20622 18232 20628 18284
rect 20680 18232 20686 18284
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20772 18244 20821 18272
rect 20772 18232 20778 18244
rect 20809 18241 20821 18244
rect 20855 18272 20867 18275
rect 21818 18272 21824 18284
rect 20855 18244 21824 18272
rect 20855 18241 20867 18244
rect 20809 18235 20867 18241
rect 21818 18232 21824 18244
rect 21876 18272 21882 18284
rect 22002 18272 22008 18284
rect 21876 18244 22008 18272
rect 21876 18232 21882 18244
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 20349 18207 20407 18213
rect 20349 18173 20361 18207
rect 20395 18173 20407 18207
rect 20640 18204 20668 18232
rect 21634 18204 21640 18216
rect 20349 18167 20407 18173
rect 20548 18176 21640 18204
rect 19794 18136 19800 18148
rect 18524 18108 19800 18136
rect 15286 18068 15292 18080
rect 15028 18040 15292 18068
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 17788 18068 17816 18108
rect 19794 18096 19800 18108
rect 19852 18096 19858 18148
rect 20548 18145 20576 18176
rect 21634 18164 21640 18176
rect 21692 18164 21698 18216
rect 24486 18164 24492 18216
rect 24544 18204 24550 18216
rect 27065 18207 27123 18213
rect 27065 18204 27077 18207
rect 24544 18176 27077 18204
rect 24544 18164 24550 18176
rect 27065 18173 27077 18176
rect 27111 18173 27123 18207
rect 27065 18167 27123 18173
rect 27157 18207 27215 18213
rect 27157 18173 27169 18207
rect 27203 18204 27215 18207
rect 27341 18207 27399 18213
rect 27341 18204 27353 18207
rect 27203 18176 27353 18204
rect 27203 18173 27215 18176
rect 27157 18167 27215 18173
rect 27341 18173 27353 18176
rect 27387 18173 27399 18207
rect 27341 18167 27399 18173
rect 20441 18139 20499 18145
rect 20441 18105 20453 18139
rect 20487 18105 20499 18139
rect 20441 18099 20499 18105
rect 20533 18139 20591 18145
rect 20533 18105 20545 18139
rect 20579 18105 20591 18139
rect 20533 18099 20591 18105
rect 20671 18139 20729 18145
rect 20671 18105 20683 18139
rect 20717 18136 20729 18139
rect 21726 18136 21732 18148
rect 20717 18108 21732 18136
rect 20717 18105 20729 18108
rect 20671 18099 20729 18105
rect 16448 18040 17816 18068
rect 17865 18071 17923 18077
rect 16448 18028 16454 18040
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 18046 18068 18052 18080
rect 17911 18040 18052 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 19702 18028 19708 18080
rect 19760 18068 19766 18080
rect 20165 18071 20223 18077
rect 20165 18068 20177 18071
rect 19760 18040 20177 18068
rect 19760 18028 19766 18040
rect 20165 18037 20177 18040
rect 20211 18037 20223 18071
rect 20456 18068 20484 18099
rect 21726 18096 21732 18108
rect 21784 18096 21790 18148
rect 20806 18068 20812 18080
rect 20456 18040 20812 18068
rect 20165 18031 20223 18037
rect 20806 18028 20812 18040
rect 20864 18028 20870 18080
rect 27080 18068 27108 18167
rect 27430 18164 27436 18216
rect 27488 18204 27494 18216
rect 27597 18207 27655 18213
rect 27597 18204 27609 18207
rect 27488 18176 27609 18204
rect 27488 18164 27494 18176
rect 27597 18173 27609 18176
rect 27643 18173 27655 18207
rect 27597 18167 27655 18173
rect 28994 18164 29000 18216
rect 29052 18164 29058 18216
rect 29264 18207 29322 18213
rect 29264 18173 29276 18207
rect 29310 18204 29322 18207
rect 29546 18204 29552 18216
rect 29310 18176 29552 18204
rect 29310 18173 29322 18176
rect 29264 18167 29322 18173
rect 29546 18164 29552 18176
rect 29604 18164 29610 18216
rect 27982 18068 27988 18080
rect 27080 18040 27988 18068
rect 27982 18028 27988 18040
rect 28040 18028 28046 18080
rect 28718 18028 28724 18080
rect 28776 18028 28782 18080
rect 552 17978 31648 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 12096 17978
rect 12148 17926 12160 17978
rect 12212 17926 12224 17978
rect 12276 17926 12288 17978
rect 12340 17926 12352 17978
rect 12404 17926 19870 17978
rect 19922 17926 19934 17978
rect 19986 17926 19998 17978
rect 20050 17926 20062 17978
rect 20114 17926 20126 17978
rect 20178 17926 27644 17978
rect 27696 17926 27708 17978
rect 27760 17926 27772 17978
rect 27824 17926 27836 17978
rect 27888 17926 27900 17978
rect 27952 17926 31648 17978
rect 552 17904 31648 17926
rect 15197 17867 15255 17873
rect 15197 17833 15209 17867
rect 15243 17864 15255 17867
rect 15286 17864 15292 17876
rect 15243 17836 15292 17864
rect 15243 17833 15255 17836
rect 15197 17827 15255 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 17313 17867 17371 17873
rect 17313 17864 17325 17867
rect 17000 17836 17325 17864
rect 17000 17824 17006 17836
rect 17313 17833 17325 17836
rect 17359 17833 17371 17867
rect 17313 17827 17371 17833
rect 19610 17824 19616 17876
rect 19668 17824 19674 17876
rect 20717 17867 20775 17873
rect 20717 17833 20729 17867
rect 20763 17864 20775 17867
rect 20806 17864 20812 17876
rect 20763 17836 20812 17864
rect 20763 17833 20775 17836
rect 20717 17827 20775 17833
rect 20806 17824 20812 17836
rect 20864 17824 20870 17876
rect 21910 17864 21916 17876
rect 21560 17836 21916 17864
rect 15746 17796 15752 17808
rect 14752 17768 15752 17796
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14752 17737 14780 17768
rect 15746 17756 15752 17768
rect 15804 17796 15810 17808
rect 16390 17796 16396 17808
rect 15804 17768 16396 17796
rect 15804 17756 15810 17768
rect 16390 17756 16396 17768
rect 16448 17756 16454 17808
rect 17494 17756 17500 17808
rect 17552 17796 17558 17808
rect 17862 17796 17868 17808
rect 17552 17768 17868 17796
rect 17552 17756 17558 17768
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 19628 17796 19656 17824
rect 21560 17805 21588 17836
rect 21910 17824 21916 17836
rect 21968 17864 21974 17876
rect 26510 17864 26516 17876
rect 21968 17836 26516 17864
rect 21968 17824 21974 17836
rect 26510 17824 26516 17836
rect 26568 17824 26574 17876
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 29181 17867 29239 17873
rect 29181 17864 29193 17867
rect 29052 17836 29193 17864
rect 29052 17824 29058 17836
rect 29181 17833 29193 17836
rect 29227 17833 29239 17867
rect 29181 17827 29239 17833
rect 19352 17768 19656 17796
rect 21545 17799 21603 17805
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 13964 17700 14657 17728
rect 13964 17688 13970 17700
rect 14645 17697 14657 17700
rect 14691 17697 14703 17731
rect 14645 17691 14703 17697
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 14826 17688 14832 17740
rect 14884 17688 14890 17740
rect 15013 17731 15071 17737
rect 15013 17697 15025 17731
rect 15059 17728 15071 17731
rect 15378 17728 15384 17740
rect 15059 17700 15384 17728
rect 15059 17697 15071 17700
rect 15013 17691 15071 17697
rect 15378 17688 15384 17700
rect 15436 17728 15442 17740
rect 16022 17728 16028 17740
rect 15436 17700 16028 17728
rect 15436 17688 15442 17700
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 16574 17688 16580 17740
rect 16632 17688 16638 17740
rect 17586 17688 17592 17740
rect 17644 17728 17650 17740
rect 18046 17737 18052 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 17644 17700 17693 17728
rect 17644 17688 17650 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 18040 17728 18052 17737
rect 18007 17700 18052 17728
rect 17681 17691 17739 17697
rect 18040 17691 18052 17700
rect 18046 17688 18052 17691
rect 18104 17688 18110 17740
rect 19352 17737 19380 17768
rect 21545 17765 21557 17799
rect 21591 17765 21603 17799
rect 21545 17759 21603 17765
rect 21634 17756 21640 17808
rect 21692 17796 21698 17808
rect 22465 17799 22523 17805
rect 22465 17796 22477 17799
rect 21692 17768 22477 17796
rect 21692 17756 21698 17768
rect 22465 17765 22477 17768
rect 22511 17765 22523 17799
rect 22465 17759 22523 17765
rect 22557 17799 22615 17805
rect 22557 17765 22569 17799
rect 22603 17796 22615 17799
rect 23750 17796 23756 17808
rect 22603 17768 23756 17796
rect 22603 17765 22615 17768
rect 22557 17759 22615 17765
rect 23750 17756 23756 17768
rect 23808 17756 23814 17808
rect 24765 17799 24823 17805
rect 24765 17765 24777 17799
rect 24811 17796 24823 17799
rect 25774 17796 25780 17808
rect 24811 17768 25780 17796
rect 24811 17765 24823 17768
rect 24765 17759 24823 17765
rect 25774 17756 25780 17768
rect 25832 17756 25838 17808
rect 19610 17737 19616 17740
rect 19337 17731 19395 17737
rect 19337 17697 19349 17731
rect 19383 17697 19395 17731
rect 19337 17691 19395 17697
rect 19604 17691 19616 17737
rect 19610 17688 19616 17691
rect 19668 17688 19674 17740
rect 20530 17688 20536 17740
rect 20588 17728 20594 17740
rect 21358 17728 21364 17740
rect 20588 17700 21364 17728
rect 20588 17688 20594 17700
rect 21358 17688 21364 17700
rect 21416 17728 21422 17740
rect 21453 17731 21511 17737
rect 21453 17728 21465 17731
rect 21416 17700 21465 17728
rect 21416 17688 21422 17700
rect 21453 17697 21465 17700
rect 21499 17697 21511 17731
rect 21453 17691 21511 17697
rect 21726 17688 21732 17740
rect 21784 17737 21790 17740
rect 21784 17731 21813 17737
rect 21801 17697 21813 17731
rect 21784 17691 21813 17697
rect 21784 17688 21790 17691
rect 22002 17688 22008 17740
rect 22060 17728 22066 17740
rect 22189 17731 22247 17737
rect 22189 17728 22201 17731
rect 22060 17700 22201 17728
rect 22060 17688 22066 17700
rect 22189 17697 22201 17700
rect 22235 17697 22247 17731
rect 22189 17691 22247 17697
rect 22347 17731 22405 17737
rect 22347 17697 22359 17731
rect 22393 17697 22405 17731
rect 22347 17691 22405 17697
rect 22649 17731 22707 17737
rect 22649 17697 22661 17731
rect 22695 17728 22707 17731
rect 23014 17728 23020 17740
rect 22695 17700 23020 17728
rect 22695 17697 22707 17700
rect 22649 17691 22707 17697
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15344 17632 15761 17660
rect 15344 17620 15350 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 17770 17620 17776 17672
rect 17828 17620 17834 17672
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21913 17663 21971 17669
rect 21913 17660 21925 17663
rect 21324 17632 21925 17660
rect 21324 17620 21330 17632
rect 21913 17629 21925 17632
rect 21959 17660 21971 17663
rect 22094 17660 22100 17672
rect 21959 17632 22100 17660
rect 21959 17629 21971 17632
rect 21913 17623 21971 17629
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 22362 17660 22390 17691
rect 23014 17688 23020 17700
rect 23072 17688 23078 17740
rect 23106 17688 23112 17740
rect 23164 17688 23170 17740
rect 23216 17700 23428 17728
rect 22554 17660 22560 17672
rect 22362 17632 22560 17660
rect 22554 17620 22560 17632
rect 22612 17660 22618 17672
rect 23216 17660 23244 17700
rect 22612 17632 23244 17660
rect 22612 17620 22618 17632
rect 23290 17620 23296 17672
rect 23348 17620 23354 17672
rect 23400 17660 23428 17700
rect 24486 17688 24492 17740
rect 24544 17688 24550 17740
rect 24670 17688 24676 17740
rect 24728 17688 24734 17740
rect 25225 17731 25283 17737
rect 25225 17697 25237 17731
rect 25271 17697 25283 17731
rect 25225 17691 25283 17697
rect 24394 17660 24400 17672
rect 23400 17632 24400 17660
rect 24394 17620 24400 17632
rect 24452 17660 24458 17672
rect 24762 17660 24768 17672
rect 24452 17632 24768 17660
rect 24452 17620 24458 17632
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25133 17663 25191 17669
rect 25133 17660 25145 17663
rect 24872 17632 25145 17660
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 24872 17592 24900 17632
rect 25133 17629 25145 17632
rect 25179 17629 25191 17663
rect 25233 17660 25261 17691
rect 25682 17688 25688 17740
rect 25740 17728 25746 17740
rect 25899 17731 25957 17737
rect 25899 17728 25911 17731
rect 25740 17700 25911 17728
rect 25740 17688 25746 17700
rect 25899 17697 25911 17700
rect 25945 17697 25957 17731
rect 25899 17691 25957 17697
rect 26050 17688 26056 17740
rect 26108 17688 26114 17740
rect 27982 17688 27988 17740
rect 28040 17728 28046 17740
rect 29089 17731 29147 17737
rect 29089 17728 29101 17731
rect 28040 17700 29101 17728
rect 28040 17688 28046 17700
rect 29089 17697 29101 17700
rect 29135 17697 29147 17731
rect 29089 17691 29147 17697
rect 28718 17660 28724 17672
rect 25233 17632 28724 17660
rect 25133 17623 25191 17629
rect 28718 17620 28724 17632
rect 28776 17620 28782 17672
rect 23072 17564 24900 17592
rect 23072 17552 23078 17564
rect 25498 17552 25504 17604
rect 25556 17592 25562 17604
rect 25685 17595 25743 17601
rect 25685 17592 25697 17595
rect 25556 17564 25697 17592
rect 25556 17552 25562 17564
rect 25685 17561 25697 17564
rect 25731 17561 25743 17595
rect 25685 17555 25743 17561
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 14240 17496 14381 17524
rect 14240 17484 14246 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 14369 17487 14427 17493
rect 19058 17484 19064 17536
rect 19116 17524 19122 17536
rect 19153 17527 19211 17533
rect 19153 17524 19165 17527
rect 19116 17496 19165 17524
rect 19116 17484 19122 17496
rect 19153 17493 19165 17496
rect 19199 17493 19211 17527
rect 19153 17487 19211 17493
rect 21266 17484 21272 17536
rect 21324 17484 21330 17536
rect 21818 17484 21824 17536
rect 21876 17524 21882 17536
rect 22833 17527 22891 17533
rect 22833 17524 22845 17527
rect 21876 17496 22845 17524
rect 21876 17484 21882 17496
rect 22833 17493 22845 17496
rect 22879 17493 22891 17527
rect 22833 17487 22891 17493
rect 22922 17484 22928 17536
rect 22980 17484 22986 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 24268 17496 24409 17524
rect 24268 17484 24274 17496
rect 24397 17493 24409 17496
rect 24443 17493 24455 17527
rect 24397 17487 24455 17493
rect 25593 17527 25651 17533
rect 25593 17493 25605 17527
rect 25639 17524 25651 17527
rect 26234 17524 26240 17536
rect 25639 17496 26240 17524
rect 25639 17493 25651 17496
rect 25593 17487 25651 17493
rect 26234 17484 26240 17496
rect 26292 17484 26298 17536
rect 552 17434 31648 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 11436 17434
rect 11488 17382 11500 17434
rect 11552 17382 11564 17434
rect 11616 17382 11628 17434
rect 11680 17382 11692 17434
rect 11744 17382 19210 17434
rect 19262 17382 19274 17434
rect 19326 17382 19338 17434
rect 19390 17382 19402 17434
rect 19454 17382 19466 17434
rect 19518 17382 26984 17434
rect 27036 17382 27048 17434
rect 27100 17382 27112 17434
rect 27164 17382 27176 17434
rect 27228 17382 27240 17434
rect 27292 17382 31648 17434
rect 552 17360 31648 17382
rect 15286 17280 15292 17332
rect 15344 17280 15350 17332
rect 15381 17323 15439 17329
rect 15381 17289 15393 17323
rect 15427 17320 15439 17323
rect 15470 17320 15476 17332
rect 15427 17292 15476 17320
rect 15427 17289 15439 17292
rect 15381 17283 15439 17289
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 17770 17280 17776 17332
rect 17828 17320 17834 17332
rect 17957 17323 18015 17329
rect 17957 17320 17969 17323
rect 17828 17292 17969 17320
rect 17828 17280 17834 17292
rect 17957 17289 17969 17292
rect 18003 17289 18015 17323
rect 17957 17283 18015 17289
rect 19429 17323 19487 17329
rect 19429 17289 19441 17323
rect 19475 17320 19487 17323
rect 19610 17320 19616 17332
rect 19475 17292 19616 17320
rect 19475 17289 19487 17292
rect 19429 17283 19487 17289
rect 19610 17280 19616 17292
rect 19668 17280 19674 17332
rect 20714 17320 20720 17332
rect 20088 17292 20720 17320
rect 17681 17255 17739 17261
rect 17681 17221 17693 17255
rect 17727 17252 17739 17255
rect 18322 17252 18328 17264
rect 17727 17224 18328 17252
rect 17727 17221 17739 17224
rect 17681 17215 17739 17221
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 20088 17184 20116 17292
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 21821 17323 21879 17329
rect 21821 17289 21833 17323
rect 21867 17320 21879 17323
rect 21910 17320 21916 17332
rect 21867 17292 21916 17320
rect 21867 17289 21879 17292
rect 21821 17283 21879 17289
rect 21910 17280 21916 17292
rect 21968 17280 21974 17332
rect 22830 17280 22836 17332
rect 22888 17320 22894 17332
rect 23569 17323 23627 17329
rect 23569 17320 23581 17323
rect 22888 17292 23581 17320
rect 22888 17280 22894 17292
rect 23569 17289 23581 17292
rect 23615 17320 23627 17323
rect 24670 17320 24676 17332
rect 23615 17292 24676 17320
rect 23615 17289 23627 17292
rect 23569 17283 23627 17289
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 26237 17323 26295 17329
rect 26237 17289 26249 17323
rect 26283 17320 26295 17323
rect 26326 17320 26332 17332
rect 26283 17292 26332 17320
rect 26283 17289 26295 17292
rect 26237 17283 26295 17289
rect 26326 17280 26332 17292
rect 26384 17280 26390 17332
rect 26602 17280 26608 17332
rect 26660 17320 26666 17332
rect 26973 17323 27031 17329
rect 26660 17292 26924 17320
rect 26660 17280 26666 17292
rect 24026 17212 24032 17264
rect 24084 17212 24090 17264
rect 24302 17212 24308 17264
rect 24360 17252 24366 17264
rect 24360 17224 24532 17252
rect 24360 17212 24366 17224
rect 15672 17156 20116 17184
rect 20257 17187 20315 17193
rect 13630 17076 13636 17128
rect 13688 17076 13694 17128
rect 14182 17125 14188 17128
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17116 13783 17119
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13771 17088 13921 17116
rect 13771 17085 13783 17088
rect 13725 17079 13783 17085
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 14176 17116 14188 17125
rect 14143 17088 14188 17116
rect 13909 17079 13967 17085
rect 14176 17079 14188 17088
rect 14182 17076 14188 17079
rect 14240 17076 14246 17128
rect 15672 17125 15700 17156
rect 20257 17153 20269 17187
rect 20303 17184 20315 17187
rect 20441 17187 20499 17193
rect 20441 17184 20453 17187
rect 20303 17156 20453 17184
rect 20303 17153 20315 17156
rect 20257 17147 20315 17153
rect 20441 17153 20453 17156
rect 20487 17153 20499 17187
rect 24044 17184 24072 17212
rect 24504 17193 24532 17224
rect 25884 17224 26832 17252
rect 24489 17187 24547 17193
rect 24044 17156 24165 17184
rect 20441 17147 20499 17153
rect 15657 17119 15715 17125
rect 15657 17085 15669 17119
rect 15703 17085 15715 17119
rect 15657 17079 15715 17085
rect 15746 17076 15752 17128
rect 15804 17076 15810 17128
rect 15838 17076 15844 17128
rect 15896 17076 15902 17128
rect 16022 17076 16028 17128
rect 16080 17076 16086 17128
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 17586 17116 17592 17128
rect 17359 17088 17592 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18874 17116 18880 17128
rect 18095 17088 18880 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18874 17076 18880 17088
rect 18932 17076 18938 17128
rect 19613 17119 19671 17125
rect 19613 17085 19625 17119
rect 19659 17116 19671 17119
rect 19702 17116 19708 17128
rect 19659 17088 19708 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 19702 17076 19708 17088
rect 19760 17076 19766 17128
rect 19794 17076 19800 17128
rect 19852 17076 19858 17128
rect 20349 17119 20407 17125
rect 20349 17085 20361 17119
rect 20395 17116 20407 17119
rect 21542 17116 21548 17128
rect 20395 17088 21548 17116
rect 20395 17085 20407 17088
rect 20349 17079 20407 17085
rect 21542 17076 21548 17088
rect 21600 17116 21606 17128
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21600 17088 21925 17116
rect 21600 17076 21606 17088
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 22005 17119 22063 17125
rect 22005 17085 22017 17119
rect 22051 17116 22063 17119
rect 22189 17119 22247 17125
rect 22189 17116 22201 17119
rect 22051 17088 22201 17116
rect 22051 17085 22063 17088
rect 22005 17079 22063 17085
rect 22189 17085 22201 17088
rect 22235 17085 22247 17119
rect 22189 17079 22247 17085
rect 22456 17119 22514 17125
rect 22456 17085 22468 17119
rect 22502 17116 22514 17119
rect 22922 17116 22928 17128
rect 22502 17088 22928 17116
rect 22502 17085 22514 17088
rect 22456 17079 22514 17085
rect 22922 17076 22928 17088
rect 22980 17076 22986 17128
rect 23658 17076 23664 17128
rect 23716 17116 23722 17128
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23716 17088 24041 17116
rect 23716 17076 23722 17088
rect 24029 17085 24041 17088
rect 24075 17085 24087 17119
rect 24137 17118 24165 17156
rect 24489 17153 24501 17187
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 24578 17144 24584 17196
rect 24636 17144 24642 17196
rect 25590 17184 25596 17196
rect 24964 17156 25596 17184
rect 24394 17125 24400 17128
rect 24213 17119 24271 17125
rect 24213 17118 24225 17119
rect 24137 17090 24225 17118
rect 24029 17079 24087 17085
rect 24213 17085 24225 17090
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 24351 17119 24400 17125
rect 24351 17085 24363 17119
rect 24397 17085 24400 17119
rect 24351 17079 24400 17085
rect 24394 17076 24400 17079
rect 24452 17076 24458 17128
rect 24854 17076 24860 17128
rect 24912 17076 24918 17128
rect 24964 17125 24992 17156
rect 25590 17144 25596 17156
rect 25648 17184 25654 17196
rect 25884 17193 25912 17224
rect 25869 17187 25927 17193
rect 25869 17184 25881 17187
rect 25648 17156 25881 17184
rect 25648 17144 25654 17156
rect 25869 17153 25881 17156
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 26068 17156 26740 17184
rect 24949 17119 25007 17125
rect 24949 17085 24961 17119
rect 24995 17085 25007 17119
rect 24949 17079 25007 17085
rect 25038 17076 25044 17128
rect 25096 17076 25102 17128
rect 25498 17076 25504 17128
rect 25556 17076 25562 17128
rect 25685 17119 25743 17125
rect 25685 17085 25697 17119
rect 25731 17085 25743 17119
rect 25685 17079 25743 17085
rect 25777 17119 25835 17125
rect 25777 17085 25789 17119
rect 25823 17116 25835 17119
rect 25958 17116 25964 17128
rect 25823 17088 25964 17116
rect 25823 17085 25835 17088
rect 25777 17079 25835 17085
rect 17497 17051 17555 17057
rect 17497 17017 17509 17051
rect 17543 17048 17555 17051
rect 19058 17048 19064 17060
rect 17543 17020 19064 17048
rect 17543 17017 17555 17020
rect 17497 17011 17555 17017
rect 19058 17008 19064 17020
rect 19116 17008 19122 17060
rect 19610 16940 19616 16992
rect 19668 16980 19674 16992
rect 19812 16980 19840 17076
rect 20530 17008 20536 17060
rect 20588 17048 20594 17060
rect 24762 17057 24768 17060
rect 20686 17051 20744 17057
rect 20686 17048 20698 17051
rect 20588 17020 20698 17048
rect 20588 17008 20594 17020
rect 20686 17017 20698 17020
rect 20732 17017 20744 17051
rect 24122 17051 24180 17057
rect 24122 17048 24134 17051
rect 20686 17011 20744 17017
rect 24116 17017 24134 17048
rect 24168 17017 24180 17051
rect 24116 17011 24180 17017
rect 24739 17051 24768 17057
rect 24739 17017 24751 17051
rect 24739 17011 24768 17017
rect 19668 16952 19840 16980
rect 19668 16940 19674 16952
rect 23658 16940 23664 16992
rect 23716 16980 23722 16992
rect 23845 16983 23903 16989
rect 23845 16980 23857 16983
rect 23716 16952 23857 16980
rect 23716 16940 23722 16952
rect 23845 16949 23857 16952
rect 23891 16949 23903 16983
rect 24116 16980 24144 17011
rect 24762 17008 24768 17011
rect 24820 17008 24826 17060
rect 25700 17048 25728 17079
rect 25958 17076 25964 17088
rect 26016 17076 26022 17128
rect 26068 17125 26096 17156
rect 26053 17119 26111 17125
rect 26053 17085 26065 17119
rect 26099 17085 26111 17119
rect 26053 17079 26111 17085
rect 26234 17076 26240 17128
rect 26292 17116 26298 17128
rect 26329 17119 26387 17125
rect 26329 17116 26341 17119
rect 26292 17088 26341 17116
rect 26292 17076 26298 17088
rect 26329 17085 26341 17088
rect 26375 17085 26387 17119
rect 26329 17079 26387 17085
rect 26418 17076 26424 17128
rect 26476 17116 26482 17128
rect 26476 17088 26521 17116
rect 26476 17076 26482 17088
rect 26712 17057 26740 17156
rect 26804 17125 26832 17224
rect 26794 17119 26852 17125
rect 26794 17085 26806 17119
rect 26840 17085 26852 17119
rect 26896 17116 26924 17292
rect 26973 17289 26985 17323
rect 27019 17320 27031 17323
rect 27522 17320 27528 17332
rect 27019 17292 27528 17320
rect 27019 17289 27031 17292
rect 26973 17283 27031 17289
rect 27522 17280 27528 17292
rect 27580 17280 27586 17332
rect 27246 17116 27252 17128
rect 26896 17088 27252 17116
rect 26794 17079 26852 17085
rect 27246 17076 27252 17088
rect 27304 17076 27310 17128
rect 26605 17051 26663 17057
rect 26605 17048 26617 17051
rect 25148 17020 26617 17048
rect 25148 16992 25176 17020
rect 26605 17017 26617 17020
rect 26651 17017 26663 17051
rect 26605 17011 26663 17017
rect 26697 17051 26755 17057
rect 26697 17017 26709 17051
rect 26743 17048 26755 17051
rect 27157 17051 27215 17057
rect 27157 17048 27169 17051
rect 26743 17020 27169 17048
rect 26743 17017 26755 17020
rect 26697 17011 26755 17017
rect 27157 17017 27169 17020
rect 27203 17017 27215 17051
rect 27157 17011 27215 17017
rect 25130 16980 25136 16992
rect 24116 16952 25136 16980
rect 23845 16943 23903 16949
rect 25130 16940 25136 16952
rect 25188 16940 25194 16992
rect 25225 16983 25283 16989
rect 25225 16949 25237 16983
rect 25271 16980 25283 16983
rect 25866 16980 25872 16992
rect 25271 16952 25872 16980
rect 25271 16949 25283 16952
rect 25225 16943 25283 16949
rect 25866 16940 25872 16952
rect 25924 16940 25930 16992
rect 25958 16940 25964 16992
rect 26016 16980 26022 16992
rect 26418 16980 26424 16992
rect 26016 16952 26424 16980
rect 26016 16940 26022 16952
rect 26418 16940 26424 16952
rect 26476 16940 26482 16992
rect 552 16890 31648 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 12096 16890
rect 12148 16838 12160 16890
rect 12212 16838 12224 16890
rect 12276 16838 12288 16890
rect 12340 16838 12352 16890
rect 12404 16838 19870 16890
rect 19922 16838 19934 16890
rect 19986 16838 19998 16890
rect 20050 16838 20062 16890
rect 20114 16838 20126 16890
rect 20178 16838 27644 16890
rect 27696 16838 27708 16890
rect 27760 16838 27772 16890
rect 27824 16838 27836 16890
rect 27888 16838 27900 16890
rect 27952 16838 31648 16890
rect 552 16816 31648 16838
rect 17313 16779 17371 16785
rect 17313 16745 17325 16779
rect 17359 16776 17371 16779
rect 18322 16776 18328 16788
rect 17359 16748 18328 16776
rect 17359 16745 17371 16748
rect 17313 16739 17371 16745
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 20530 16736 20536 16788
rect 20588 16736 20594 16788
rect 23014 16776 23020 16788
rect 21560 16748 23020 16776
rect 16666 16708 16672 16720
rect 16408 16680 16672 16708
rect 15286 16600 15292 16652
rect 15344 16600 15350 16652
rect 15470 16649 15476 16652
rect 15443 16643 15476 16649
rect 15443 16609 15455 16643
rect 15443 16603 15476 16609
rect 15470 16600 15476 16603
rect 15528 16600 15534 16652
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 16408 16649 16436 16680
rect 16666 16668 16672 16680
rect 16724 16708 16730 16720
rect 17034 16708 17040 16720
rect 16724 16680 17040 16708
rect 16724 16668 16730 16680
rect 17034 16668 17040 16680
rect 17092 16668 17098 16720
rect 17957 16711 18015 16717
rect 17957 16677 17969 16711
rect 18003 16708 18015 16711
rect 18230 16708 18236 16720
rect 18003 16680 18236 16708
rect 18003 16677 18015 16680
rect 17957 16671 18015 16677
rect 18230 16668 18236 16680
rect 18288 16708 18294 16720
rect 21560 16717 21588 16748
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 23106 16736 23112 16788
rect 23164 16736 23170 16788
rect 23474 16736 23480 16788
rect 23532 16776 23538 16788
rect 25038 16776 25044 16788
rect 23532 16748 25044 16776
rect 23532 16736 23538 16748
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 25590 16736 25596 16788
rect 25648 16736 25654 16788
rect 27246 16736 27252 16788
rect 27304 16776 27310 16788
rect 27304 16748 27660 16776
rect 27304 16736 27310 16748
rect 21545 16711 21603 16717
rect 18288 16680 18644 16708
rect 18288 16668 18294 16680
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15712 16612 16129 16640
rect 15712 16600 15718 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16393 16643 16451 16649
rect 16393 16609 16405 16643
rect 16439 16609 16451 16643
rect 16393 16603 16451 16609
rect 16482 16600 16488 16652
rect 16540 16600 16546 16652
rect 17126 16600 17132 16652
rect 17184 16600 17190 16652
rect 17402 16600 17408 16652
rect 17460 16600 17466 16652
rect 18506 16600 18512 16652
rect 18564 16600 18570 16652
rect 18616 16649 18644 16680
rect 21545 16677 21557 16711
rect 21591 16677 21603 16711
rect 21545 16671 21603 16677
rect 21634 16668 21640 16720
rect 21692 16668 21698 16720
rect 21726 16668 21732 16720
rect 21784 16717 21790 16720
rect 21784 16711 21833 16717
rect 21784 16677 21787 16711
rect 21821 16677 21833 16711
rect 21784 16671 21833 16677
rect 21784 16668 21790 16671
rect 22554 16668 22560 16720
rect 22612 16717 22618 16720
rect 22612 16711 22661 16717
rect 22612 16677 22615 16711
rect 22649 16677 22661 16711
rect 22612 16671 22661 16677
rect 22612 16668 22618 16671
rect 22830 16668 22836 16720
rect 22888 16668 22894 16720
rect 23290 16668 23296 16720
rect 23348 16708 23354 16720
rect 23348 16680 26004 16708
rect 23348 16668 23354 16680
rect 18602 16643 18660 16649
rect 18602 16609 18614 16643
rect 18648 16609 18660 16643
rect 18602 16603 18660 16609
rect 18874 16600 18880 16652
rect 18932 16640 18938 16652
rect 19702 16640 19708 16652
rect 18932 16612 19708 16640
rect 18932 16600 18938 16612
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 20717 16643 20775 16649
rect 20717 16609 20729 16643
rect 20763 16640 20775 16643
rect 21266 16640 21272 16652
rect 20763 16612 21272 16640
rect 20763 16609 20775 16612
rect 20717 16603 20775 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 21453 16643 21511 16649
rect 21453 16640 21465 16643
rect 21416 16612 21465 16640
rect 21416 16600 21422 16612
rect 21453 16609 21465 16612
rect 21499 16609 21511 16643
rect 21453 16603 21511 16609
rect 15657 16507 15715 16513
rect 15657 16473 15669 16507
rect 15703 16504 15715 16507
rect 16114 16504 16120 16516
rect 15703 16476 16120 16504
rect 15703 16473 15715 16476
rect 15657 16467 15715 16473
rect 16114 16464 16120 16476
rect 16172 16464 16178 16516
rect 18325 16507 18383 16513
rect 18325 16473 18337 16507
rect 18371 16504 18383 16507
rect 18524 16504 18552 16600
rect 19610 16532 19616 16584
rect 19668 16572 19674 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 19668 16544 20913 16572
rect 19668 16532 19674 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 21652 16572 21680 16668
rect 21913 16643 21971 16649
rect 21913 16609 21925 16643
rect 21959 16640 21971 16643
rect 22462 16640 22468 16652
rect 21959 16612 22468 16640
rect 21959 16609 21971 16612
rect 21913 16603 21971 16609
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 22741 16643 22799 16649
rect 22741 16609 22753 16643
rect 22787 16609 22799 16643
rect 22741 16603 22799 16609
rect 22925 16643 22983 16649
rect 22925 16609 22937 16643
rect 22971 16640 22983 16643
rect 23474 16640 23480 16652
rect 22971 16612 23480 16640
rect 22971 16609 22983 16612
rect 22925 16603 22983 16609
rect 22756 16572 22784 16603
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 23584 16649 23612 16680
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 23658 16600 23664 16652
rect 23716 16600 23722 16652
rect 24210 16600 24216 16652
rect 24268 16600 24274 16652
rect 24480 16643 24538 16649
rect 24480 16609 24492 16643
rect 24526 16640 24538 16643
rect 25685 16643 25743 16649
rect 25685 16640 25697 16643
rect 24526 16612 25697 16640
rect 24526 16609 24538 16612
rect 24480 16603 24538 16609
rect 25685 16609 25697 16612
rect 25731 16609 25743 16643
rect 25685 16603 25743 16609
rect 25866 16600 25872 16652
rect 25924 16600 25930 16652
rect 25976 16649 26004 16680
rect 26786 16668 26792 16720
rect 26844 16708 26850 16720
rect 26844 16680 27568 16708
rect 26844 16668 26850 16680
rect 25961 16643 26019 16649
rect 25961 16609 25973 16643
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 26878 16600 26884 16652
rect 26936 16600 26942 16652
rect 27249 16643 27307 16649
rect 27249 16609 27261 16643
rect 27295 16640 27307 16643
rect 27338 16640 27344 16652
rect 27295 16612 27344 16640
rect 27295 16609 27307 16612
rect 27249 16603 27307 16609
rect 27338 16600 27344 16612
rect 27396 16600 27402 16652
rect 27430 16600 27436 16652
rect 27488 16600 27494 16652
rect 27540 16649 27568 16680
rect 27632 16649 27660 16748
rect 27525 16643 27583 16649
rect 27525 16609 27537 16643
rect 27571 16609 27583 16643
rect 27525 16603 27583 16609
rect 27617 16643 27675 16649
rect 27617 16609 27629 16643
rect 27663 16609 27675 16643
rect 27617 16603 27675 16609
rect 27982 16600 27988 16652
rect 28040 16640 28046 16652
rect 28994 16640 29000 16652
rect 28040 16612 29000 16640
rect 28040 16600 28046 16612
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 21652 16544 22784 16572
rect 20901 16535 20959 16541
rect 18371 16476 18552 16504
rect 18877 16507 18935 16513
rect 18371 16473 18383 16476
rect 18325 16467 18383 16473
rect 18877 16473 18889 16507
rect 18923 16504 18935 16507
rect 18966 16504 18972 16516
rect 18923 16476 18972 16504
rect 18923 16473 18935 16476
rect 18877 16467 18935 16473
rect 18966 16464 18972 16476
rect 19024 16464 19030 16516
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 16209 16439 16267 16445
rect 16209 16436 16221 16439
rect 15436 16408 16221 16436
rect 15436 16396 15442 16408
rect 16209 16405 16221 16408
rect 16255 16405 16267 16439
rect 16209 16399 16267 16405
rect 16666 16396 16672 16448
rect 16724 16396 16730 16448
rect 16942 16396 16948 16448
rect 17000 16396 17006 16448
rect 17310 16396 17316 16448
rect 17368 16436 17374 16448
rect 17862 16436 17868 16448
rect 17368 16408 17868 16436
rect 17368 16396 17374 16408
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 18417 16439 18475 16445
rect 18417 16405 18429 16439
rect 18463 16436 18475 16439
rect 18598 16436 18604 16448
rect 18463 16408 18604 16436
rect 18463 16405 18475 16408
rect 18417 16399 18475 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 21269 16439 21327 16445
rect 21269 16436 21281 16439
rect 20956 16408 21281 16436
rect 20956 16396 20962 16408
rect 21269 16405 21281 16408
rect 21315 16405 21327 16439
rect 21269 16399 21327 16405
rect 23845 16439 23903 16445
rect 23845 16405 23857 16439
rect 23891 16436 23903 16439
rect 23934 16436 23940 16448
rect 23891 16408 23940 16436
rect 23891 16405 23903 16408
rect 23845 16399 23903 16405
rect 23934 16396 23940 16408
rect 23992 16396 23998 16448
rect 26418 16396 26424 16448
rect 26476 16436 26482 16448
rect 26973 16439 27031 16445
rect 26973 16436 26985 16439
rect 26476 16408 26985 16436
rect 26476 16396 26482 16408
rect 26973 16405 26985 16408
rect 27019 16405 27031 16439
rect 26973 16399 27031 16405
rect 27893 16439 27951 16445
rect 27893 16405 27905 16439
rect 27939 16436 27951 16439
rect 27982 16436 27988 16448
rect 27939 16408 27988 16436
rect 27939 16405 27951 16408
rect 27893 16399 27951 16405
rect 27982 16396 27988 16408
rect 28040 16396 28046 16448
rect 28077 16439 28135 16445
rect 28077 16405 28089 16439
rect 28123 16436 28135 16439
rect 28718 16436 28724 16448
rect 28123 16408 28724 16436
rect 28123 16405 28135 16408
rect 28077 16399 28135 16405
rect 28718 16396 28724 16408
rect 28776 16396 28782 16448
rect 552 16346 31648 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 11436 16346
rect 11488 16294 11500 16346
rect 11552 16294 11564 16346
rect 11616 16294 11628 16346
rect 11680 16294 11692 16346
rect 11744 16294 19210 16346
rect 19262 16294 19274 16346
rect 19326 16294 19338 16346
rect 19390 16294 19402 16346
rect 19454 16294 19466 16346
rect 19518 16294 26984 16346
rect 27036 16294 27048 16346
rect 27100 16294 27112 16346
rect 27164 16294 27176 16346
rect 27228 16294 27240 16346
rect 27292 16294 31648 16346
rect 552 16272 31648 16294
rect 16761 16235 16819 16241
rect 16761 16201 16773 16235
rect 16807 16232 16819 16235
rect 17126 16232 17132 16244
rect 16807 16204 17132 16232
rect 16807 16201 16819 16204
rect 16761 16195 16819 16201
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 17402 16192 17408 16244
rect 17460 16192 17466 16244
rect 17770 16232 17776 16244
rect 17512 16204 17776 16232
rect 16942 16164 16948 16176
rect 15304 16136 16948 16164
rect 15304 15960 15332 16136
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 16666 16096 16672 16108
rect 15764 16068 16672 16096
rect 15378 15988 15384 16040
rect 15436 15988 15442 16040
rect 15473 16031 15531 16037
rect 15473 15997 15485 16031
rect 15519 16028 15531 16031
rect 15654 16028 15660 16040
rect 15519 16000 15660 16028
rect 15519 15997 15531 16000
rect 15473 15991 15531 15997
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 15764 16037 15792 16068
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 17512 16096 17540 16204
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 19337 16235 19395 16241
rect 19337 16232 19349 16235
rect 18380 16204 19349 16232
rect 18380 16192 18386 16204
rect 19337 16201 19349 16204
rect 19383 16201 19395 16235
rect 19337 16195 19395 16201
rect 19518 16192 19524 16244
rect 19576 16232 19582 16244
rect 20346 16232 20352 16244
rect 19576 16204 20352 16232
rect 19576 16192 19582 16204
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 25225 16235 25283 16241
rect 25225 16232 25237 16235
rect 25188 16204 25237 16232
rect 25188 16192 25194 16204
rect 25225 16201 25237 16204
rect 25271 16201 25283 16235
rect 25225 16195 25283 16201
rect 27249 16235 27307 16241
rect 27249 16201 27261 16235
rect 27295 16232 27307 16235
rect 27430 16232 27436 16244
rect 27295 16204 27436 16232
rect 27295 16201 27307 16204
rect 27249 16195 27307 16201
rect 27430 16192 27436 16204
rect 27488 16192 27494 16244
rect 18506 16164 18512 16176
rect 17144 16068 17540 16096
rect 17604 16136 18512 16164
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15838 15988 15844 16040
rect 15896 15988 15902 16040
rect 15934 16031 15992 16037
rect 15934 15997 15946 16031
rect 15980 15997 15992 16031
rect 15934 15991 15992 15997
rect 15565 15963 15623 15969
rect 15565 15960 15577 15963
rect 15304 15932 15577 15960
rect 15565 15929 15577 15932
rect 15611 15929 15623 15963
rect 15565 15923 15623 15929
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15948 15892 15976 15991
rect 16114 15988 16120 16040
rect 16172 15988 16178 16040
rect 16390 16037 16396 16040
rect 16347 16031 16396 16037
rect 16347 15997 16359 16031
rect 16393 15997 16396 16031
rect 16347 15991 16396 15997
rect 16390 15988 16396 15991
rect 16448 15988 16454 16040
rect 16482 15988 16488 16040
rect 16540 16028 16546 16040
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 16540 16000 16957 16028
rect 16540 15988 16546 16000
rect 16945 15997 16957 16000
rect 16991 15997 17003 16031
rect 16945 15991 17003 15997
rect 17034 15988 17040 16040
rect 17092 15988 17098 16040
rect 17144 16037 17172 16068
rect 17129 16031 17187 16037
rect 17129 15997 17141 16031
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 17310 15988 17316 16040
rect 17368 15988 17374 16040
rect 17604 16037 17632 16136
rect 18506 16124 18512 16136
rect 18564 16164 18570 16176
rect 18564 16136 19104 16164
rect 18564 16124 18570 16136
rect 17770 16056 17776 16108
rect 17828 16096 17834 16108
rect 17865 16099 17923 16105
rect 17865 16096 17877 16099
rect 17828 16068 17877 16096
rect 17828 16056 17834 16068
rect 17865 16065 17877 16068
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16096 18475 16099
rect 18463 16068 18828 16096
rect 18463 16065 18475 16068
rect 18417 16059 18475 16065
rect 17589 16031 17647 16037
rect 17589 15997 17601 16031
rect 17635 15997 17647 16031
rect 17589 15991 17647 15997
rect 17681 16031 17739 16037
rect 17681 15997 17693 16031
rect 17727 16028 17739 16031
rect 17727 16000 17816 16028
rect 17727 15997 17739 16000
rect 17681 15991 17739 15997
rect 16206 15920 16212 15972
rect 16264 15920 16270 15972
rect 15243 15864 15976 15892
rect 16485 15895 16543 15901
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 16485 15861 16497 15895
rect 16531 15892 16543 15895
rect 17586 15892 17592 15904
rect 16531 15864 17592 15892
rect 16531 15861 16543 15864
rect 16485 15855 16543 15861
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 17788 15892 17816 16000
rect 17954 15988 17960 16040
rect 18012 15988 18018 16040
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18064 15960 18092 15991
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 18196 16000 18241 16028
rect 18196 15988 18202 16000
rect 18598 15988 18604 16040
rect 18656 16028 18662 16040
rect 18800 16037 18828 16068
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18656 16000 18705 16028
rect 18656 15988 18662 16000
rect 18693 15997 18705 16000
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 18786 16031 18844 16037
rect 18786 15997 18798 16031
rect 18832 15997 18844 16031
rect 18786 15991 18844 15997
rect 18966 15988 18972 16040
rect 19024 15988 19030 16040
rect 19076 16028 19104 16136
rect 26510 16124 26516 16176
rect 26568 16164 26574 16176
rect 26694 16164 26700 16176
rect 26568 16136 26700 16164
rect 26568 16124 26574 16136
rect 26694 16124 26700 16136
rect 26752 16164 26758 16176
rect 27065 16167 27123 16173
rect 27065 16164 27077 16167
rect 26752 16136 27077 16164
rect 26752 16124 26758 16136
rect 27065 16133 27077 16136
rect 27111 16133 27123 16167
rect 27065 16127 27123 16133
rect 20438 16096 20444 16108
rect 19444 16068 20444 16096
rect 19158 16031 19216 16037
rect 19158 16028 19170 16031
rect 19076 16000 19170 16028
rect 19158 15997 19170 16000
rect 19204 15997 19216 16031
rect 19158 15991 19216 15997
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19444 16037 19472 16068
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16096 20775 16099
rect 21174 16096 21180 16108
rect 20763 16068 21180 16096
rect 20763 16065 20775 16068
rect 20717 16059 20775 16065
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 28813 16099 28871 16105
rect 28813 16065 28825 16099
rect 28859 16096 28871 16099
rect 29089 16099 29147 16105
rect 29089 16096 29101 16099
rect 28859 16068 29101 16096
rect 28859 16065 28871 16068
rect 28813 16059 28871 16065
rect 29089 16065 29101 16068
rect 29135 16065 29147 16099
rect 29089 16059 29147 16065
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 19392 16000 19441 16028
rect 19392 15988 19398 16000
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 19610 15988 19616 16040
rect 19668 15988 19674 16040
rect 20898 15988 20904 16040
rect 20956 15988 20962 16040
rect 21542 15988 21548 16040
rect 21600 16028 21606 16040
rect 23477 16031 23535 16037
rect 23477 16028 23489 16031
rect 21600 16000 23489 16028
rect 21600 15988 21606 16000
rect 23477 15997 23489 16000
rect 23523 15997 23535 16031
rect 23477 15991 23535 15997
rect 23569 16031 23627 16037
rect 23569 15997 23581 16031
rect 23615 16028 23627 16031
rect 23845 16031 23903 16037
rect 23845 16028 23857 16031
rect 23615 16000 23857 16028
rect 23615 15997 23627 16000
rect 23569 15991 23627 15997
rect 23845 15997 23857 16000
rect 23891 15997 23903 16031
rect 23845 15991 23903 15997
rect 23934 15988 23940 16040
rect 23992 16028 23998 16040
rect 24101 16031 24159 16037
rect 24101 16028 24113 16031
rect 23992 16000 24113 16028
rect 23992 15988 23998 16000
rect 24101 15997 24113 16000
rect 24147 15997 24159 16031
rect 24101 15991 24159 15997
rect 26697 16031 26755 16037
rect 26697 15997 26709 16031
rect 26743 16028 26755 16031
rect 26786 16028 26792 16040
rect 26743 16000 26792 16028
rect 26743 15997 26755 16000
rect 26697 15991 26755 15997
rect 26786 15988 26792 16000
rect 26844 16028 26850 16040
rect 27157 16031 27215 16037
rect 27157 16028 27169 16031
rect 26844 16000 27169 16028
rect 26844 15988 26850 16000
rect 27157 15997 27169 16000
rect 27203 15997 27215 16031
rect 27157 15991 27215 15997
rect 27338 15988 27344 16040
rect 27396 15988 27402 16040
rect 27982 15988 27988 16040
rect 28040 16028 28046 16040
rect 28546 16031 28604 16037
rect 28546 16028 28558 16031
rect 28040 16000 28558 16028
rect 28040 15988 28046 16000
rect 28546 15997 28558 16000
rect 28592 15997 28604 16031
rect 28546 15991 28604 15997
rect 28994 15988 29000 16040
rect 29052 15988 29058 16040
rect 18414 15960 18420 15972
rect 18064 15932 18420 15960
rect 18414 15920 18420 15932
rect 18472 15920 18478 15972
rect 19058 15920 19064 15972
rect 19116 15920 19122 15972
rect 26878 15920 26884 15972
rect 26936 15920 26942 15972
rect 19076 15892 19104 15920
rect 17788 15864 19104 15892
rect 21082 15852 21088 15904
rect 21140 15852 21146 15904
rect 21266 15852 21272 15904
rect 21324 15892 21330 15904
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 21324 15864 21465 15892
rect 21324 15852 21330 15864
rect 21453 15861 21465 15864
rect 21499 15861 21511 15895
rect 21453 15855 21511 15861
rect 26234 15852 26240 15904
rect 26292 15892 26298 15904
rect 26513 15895 26571 15901
rect 26513 15892 26525 15895
rect 26292 15864 26525 15892
rect 26292 15852 26298 15864
rect 26513 15861 26525 15864
rect 26559 15861 26571 15895
rect 26513 15855 26571 15861
rect 26789 15895 26847 15901
rect 26789 15861 26801 15895
rect 26835 15892 26847 15895
rect 27356 15892 27384 15988
rect 27433 15895 27491 15901
rect 27433 15892 27445 15895
rect 26835 15864 27445 15892
rect 26835 15861 26847 15864
rect 26789 15855 26847 15861
rect 27433 15861 27445 15864
rect 27479 15861 27491 15895
rect 27433 15855 27491 15861
rect 552 15802 31648 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 12096 15802
rect 12148 15750 12160 15802
rect 12212 15750 12224 15802
rect 12276 15750 12288 15802
rect 12340 15750 12352 15802
rect 12404 15750 19870 15802
rect 19922 15750 19934 15802
rect 19986 15750 19998 15802
rect 20050 15750 20062 15802
rect 20114 15750 20126 15802
rect 20178 15750 27644 15802
rect 27696 15750 27708 15802
rect 27760 15750 27772 15802
rect 27824 15750 27836 15802
rect 27888 15750 27900 15802
rect 27952 15750 31648 15802
rect 552 15728 31648 15750
rect 15657 15691 15715 15697
rect 15657 15657 15669 15691
rect 15703 15688 15715 15691
rect 15838 15688 15844 15700
rect 15703 15660 15844 15688
rect 15703 15657 15715 15660
rect 15657 15651 15715 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16393 15691 16451 15697
rect 16393 15657 16405 15691
rect 16439 15688 16451 15691
rect 16482 15688 16488 15700
rect 16439 15660 16488 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 17770 15648 17776 15700
rect 17828 15648 17834 15700
rect 22649 15691 22707 15697
rect 22649 15657 22661 15691
rect 22695 15688 22707 15691
rect 23014 15688 23020 15700
rect 22695 15660 23020 15688
rect 22695 15657 22707 15660
rect 22649 15651 22707 15657
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 27249 15691 27307 15697
rect 27249 15657 27261 15691
rect 27295 15657 27307 15691
rect 27249 15651 27307 15657
rect 15197 15623 15255 15629
rect 15197 15589 15209 15623
rect 15243 15620 15255 15623
rect 15470 15620 15476 15632
rect 15243 15592 15476 15620
rect 15243 15589 15255 15592
rect 15197 15583 15255 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 20257 15623 20315 15629
rect 20257 15620 20269 15623
rect 19444 15592 20269 15620
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15552 16543 15555
rect 16850 15552 16856 15564
rect 16531 15524 16856 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 17865 15555 17923 15561
rect 17865 15521 17877 15555
rect 17911 15552 17923 15555
rect 18046 15552 18052 15564
rect 17911 15524 18052 15552
rect 17911 15521 17923 15524
rect 17865 15515 17923 15521
rect 18046 15512 18052 15524
rect 18104 15512 18110 15564
rect 19444 15561 19472 15592
rect 20257 15589 20269 15592
rect 20303 15589 20315 15623
rect 20257 15583 20315 15589
rect 21082 15580 21088 15632
rect 21140 15620 21146 15632
rect 21514 15623 21572 15629
rect 21514 15620 21526 15623
rect 21140 15592 21526 15620
rect 21140 15580 21146 15592
rect 21514 15589 21526 15592
rect 21560 15589 21572 15623
rect 21514 15583 21572 15589
rect 27065 15623 27123 15629
rect 27065 15589 27077 15623
rect 27111 15589 27123 15623
rect 27264 15620 27292 15651
rect 28454 15623 28512 15629
rect 28454 15620 28466 15623
rect 27264 15592 28466 15620
rect 27065 15583 27123 15589
rect 28454 15589 28466 15592
rect 28500 15589 28512 15623
rect 28454 15583 28512 15589
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 19702 15512 19708 15564
rect 19760 15552 19766 15564
rect 19889 15555 19947 15561
rect 19889 15552 19901 15555
rect 19760 15524 19901 15552
rect 19760 15512 19766 15524
rect 19889 15521 19901 15524
rect 19935 15521 19947 15555
rect 19889 15515 19947 15521
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 26418 15512 26424 15564
rect 26476 15512 26482 15564
rect 26605 15555 26663 15561
rect 26605 15521 26617 15555
rect 26651 15521 26663 15555
rect 27080 15552 27108 15583
rect 27338 15552 27344 15564
rect 27080 15524 27344 15552
rect 26605 15515 26663 15521
rect 19518 15444 19524 15496
rect 19576 15444 19582 15496
rect 20898 15444 20904 15496
rect 20956 15444 20962 15496
rect 26620 15484 26648 15515
rect 27338 15512 27344 15524
rect 27396 15512 27402 15564
rect 28718 15512 28724 15564
rect 28776 15512 28782 15564
rect 27430 15484 27436 15496
rect 26620 15456 27436 15484
rect 27430 15444 27436 15456
rect 27488 15444 27494 15496
rect 15286 15376 15292 15428
rect 15344 15416 15350 15428
rect 15473 15419 15531 15425
rect 15473 15416 15485 15419
rect 15344 15388 15485 15416
rect 15344 15376 15350 15388
rect 15473 15385 15485 15388
rect 15519 15385 15531 15419
rect 15473 15379 15531 15385
rect 19610 15376 19616 15428
rect 19668 15416 19674 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 19668 15388 19993 15416
rect 19668 15376 19674 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 26697 15419 26755 15425
rect 26697 15385 26709 15419
rect 26743 15385 26755 15419
rect 26697 15379 26755 15385
rect 19702 15308 19708 15360
rect 19760 15308 19766 15360
rect 26602 15308 26608 15360
rect 26660 15348 26666 15360
rect 26712 15348 26740 15379
rect 26878 15376 26884 15428
rect 26936 15416 26942 15428
rect 27341 15419 27399 15425
rect 27341 15416 27353 15419
rect 26936 15388 27353 15416
rect 26936 15376 26942 15388
rect 27341 15385 27353 15388
rect 27387 15385 27399 15419
rect 27341 15379 27399 15385
rect 26660 15320 26740 15348
rect 26660 15308 26666 15320
rect 26786 15308 26792 15360
rect 26844 15348 26850 15360
rect 27065 15351 27123 15357
rect 27065 15348 27077 15351
rect 26844 15320 27077 15348
rect 26844 15308 26850 15320
rect 27065 15317 27077 15320
rect 27111 15348 27123 15351
rect 27522 15348 27528 15360
rect 27111 15320 27528 15348
rect 27111 15317 27123 15320
rect 27065 15311 27123 15317
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 552 15258 31648 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 11436 15258
rect 11488 15206 11500 15258
rect 11552 15206 11564 15258
rect 11616 15206 11628 15258
rect 11680 15206 11692 15258
rect 11744 15206 19210 15258
rect 19262 15206 19274 15258
rect 19326 15206 19338 15258
rect 19390 15206 19402 15258
rect 19454 15206 19466 15258
rect 19518 15206 26984 15258
rect 27036 15206 27048 15258
rect 27100 15206 27112 15258
rect 27164 15206 27176 15258
rect 27228 15206 27240 15258
rect 27292 15206 31648 15258
rect 552 15184 31648 15206
rect 16942 15104 16948 15156
rect 17000 15104 17006 15156
rect 20898 15104 20904 15156
rect 20956 15144 20962 15156
rect 20993 15147 21051 15153
rect 20993 15144 21005 15147
rect 20956 15116 21005 15144
rect 20956 15104 20962 15116
rect 20993 15113 21005 15116
rect 21039 15113 21051 15147
rect 23290 15144 23296 15156
rect 20993 15107 21051 15113
rect 21652 15116 23296 15144
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 17865 15079 17923 15085
rect 17865 15076 17877 15079
rect 17276 15048 17877 15076
rect 17276 15036 17282 15048
rect 17865 15045 17877 15048
rect 17911 15076 17923 15079
rect 17911 15048 19380 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 16482 14968 16488 15020
rect 16540 14968 16546 15020
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 18248 14980 19257 15008
rect 18248 14952 18276 14980
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 13688 14912 14933 14940
rect 13688 14900 13694 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 14921 14903 14979 14909
rect 15933 14943 15991 14949
rect 15933 14909 15945 14943
rect 15979 14940 15991 14943
rect 16114 14940 16120 14952
rect 15979 14912 16120 14940
rect 15979 14909 15991 14912
rect 15933 14903 15991 14909
rect 14936 14872 14964 14903
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 16206 14900 16212 14952
rect 16264 14940 16270 14952
rect 16393 14943 16451 14949
rect 16393 14940 16405 14943
rect 16264 14912 16405 14940
rect 16264 14900 16270 14912
rect 16393 14909 16405 14912
rect 16439 14909 16451 14943
rect 16393 14903 16451 14909
rect 16666 14900 16672 14952
rect 16724 14900 16730 14952
rect 16761 14943 16819 14949
rect 16761 14909 16773 14943
rect 16807 14940 16819 14943
rect 17770 14940 17776 14952
rect 16807 14912 17776 14940
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 17770 14900 17776 14912
rect 17828 14900 17834 14952
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 18230 14940 18236 14952
rect 18095 14912 18236 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 18966 14940 18972 14952
rect 18380 14912 18972 14940
rect 18380 14900 18386 14912
rect 18966 14900 18972 14912
rect 19024 14900 19030 14952
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14909 19119 14943
rect 19061 14903 19119 14909
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14940 19211 14943
rect 19352 14940 19380 15048
rect 19610 14968 19616 15020
rect 19668 14968 19674 15020
rect 21652 15017 21680 15116
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 23477 15147 23535 15153
rect 23477 15113 23489 15147
rect 23523 15144 23535 15147
rect 23750 15144 23756 15156
rect 23523 15116 23756 15144
rect 23523 15113 23535 15116
rect 23477 15107 23535 15113
rect 23750 15104 23756 15116
rect 23808 15104 23814 15156
rect 26602 15144 26608 15156
rect 25240 15116 26608 15144
rect 21637 15011 21695 15017
rect 21637 14977 21649 15011
rect 21683 14977 21695 15011
rect 21637 14971 21695 14977
rect 19199 14912 19380 14940
rect 19199 14909 19211 14912
rect 19153 14903 19211 14909
rect 16574 14872 16580 14884
rect 14936 14844 16580 14872
rect 16574 14832 16580 14844
rect 16632 14832 16638 14884
rect 18138 14832 18144 14884
rect 18196 14872 18202 14884
rect 19076 14872 19104 14903
rect 19702 14900 19708 14952
rect 19760 14940 19766 14952
rect 19869 14943 19927 14949
rect 19869 14940 19881 14943
rect 19760 14912 19881 14940
rect 19760 14900 19766 14912
rect 19869 14909 19881 14912
rect 19915 14909 19927 14943
rect 19869 14903 19927 14909
rect 21818 14900 21824 14952
rect 21876 14900 21882 14952
rect 22094 14900 22100 14952
rect 22152 14900 22158 14952
rect 24949 14943 25007 14949
rect 24949 14909 24961 14943
rect 24995 14940 25007 14943
rect 25038 14940 25044 14952
rect 24995 14912 25044 14940
rect 24995 14909 25007 14912
rect 24949 14903 25007 14909
rect 25038 14900 25044 14912
rect 25096 14900 25102 14952
rect 25240 14949 25268 15116
rect 26602 15104 26608 15116
rect 26660 15104 26666 15156
rect 26694 15104 26700 15156
rect 26752 15144 26758 15156
rect 27065 15147 27123 15153
rect 27065 15144 27077 15147
rect 26752 15116 27077 15144
rect 26752 15104 26758 15116
rect 27065 15113 27077 15116
rect 27111 15113 27123 15147
rect 27065 15107 27123 15113
rect 27249 15147 27307 15153
rect 27249 15113 27261 15147
rect 27295 15144 27307 15147
rect 27338 15144 27344 15156
rect 27295 15116 27344 15144
rect 27295 15113 27307 15116
rect 27249 15107 27307 15113
rect 27338 15104 27344 15116
rect 27396 15104 27402 15156
rect 25332 14980 25820 15008
rect 25332 14949 25360 14980
rect 25133 14943 25191 14949
rect 25133 14909 25145 14943
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 25225 14943 25283 14949
rect 25225 14909 25237 14943
rect 25271 14909 25283 14943
rect 25225 14903 25283 14909
rect 25317 14943 25375 14949
rect 25317 14909 25329 14943
rect 25363 14909 25375 14943
rect 25317 14903 25375 14909
rect 20898 14872 20904 14884
rect 18196 14844 20904 14872
rect 18196 14832 18202 14844
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 22005 14875 22063 14881
rect 22005 14841 22017 14875
rect 22051 14872 22063 14875
rect 22342 14875 22400 14881
rect 22342 14872 22354 14875
rect 22051 14844 22354 14872
rect 22051 14841 22063 14844
rect 22005 14835 22063 14841
rect 22342 14841 22354 14844
rect 22388 14841 22400 14875
rect 22342 14835 22400 14841
rect 14182 14764 14188 14816
rect 14240 14804 14246 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14240 14776 14841 14804
rect 14240 14764 14246 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15436 14776 15853 14804
rect 15436 14764 15442 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 15841 14767 15899 14773
rect 18233 14807 18291 14813
rect 18233 14773 18245 14807
rect 18279 14804 18291 14807
rect 18322 14804 18328 14816
rect 18279 14776 18328 14804
rect 18279 14773 18291 14776
rect 18233 14767 18291 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 18414 14764 18420 14816
rect 18472 14764 18478 14816
rect 18785 14807 18843 14813
rect 18785 14773 18797 14807
rect 18831 14804 18843 14807
rect 18966 14804 18972 14816
rect 18831 14776 18972 14804
rect 18831 14773 18843 14776
rect 18785 14767 18843 14773
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 25148 14804 25176 14903
rect 25682 14900 25688 14952
rect 25740 14900 25746 14952
rect 25792 14940 25820 14980
rect 25792 14912 26372 14940
rect 25593 14875 25651 14881
rect 25593 14841 25605 14875
rect 25639 14872 25651 14875
rect 25930 14875 25988 14881
rect 25930 14872 25942 14875
rect 25639 14844 25942 14872
rect 25639 14841 25651 14844
rect 25593 14835 25651 14841
rect 25930 14841 25942 14844
rect 25976 14841 25988 14875
rect 26344 14872 26372 14912
rect 26418 14900 26424 14952
rect 26476 14940 26482 14952
rect 27157 14943 27215 14949
rect 27157 14940 27169 14943
rect 26476 14912 27169 14940
rect 26476 14900 26482 14912
rect 27157 14909 27169 14912
rect 27203 14909 27215 14943
rect 27157 14903 27215 14909
rect 27341 14943 27399 14949
rect 27341 14909 27353 14943
rect 27387 14940 27399 14943
rect 27430 14940 27436 14952
rect 27387 14912 27436 14940
rect 27387 14909 27399 14912
rect 27341 14903 27399 14909
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 26694 14872 26700 14884
rect 26344 14844 26700 14872
rect 25930 14835 25988 14841
rect 26694 14832 26700 14844
rect 26752 14832 26758 14884
rect 26142 14804 26148 14816
rect 25148 14776 26148 14804
rect 26142 14764 26148 14776
rect 26200 14764 26206 14816
rect 552 14714 31648 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 12096 14714
rect 12148 14662 12160 14714
rect 12212 14662 12224 14714
rect 12276 14662 12288 14714
rect 12340 14662 12352 14714
rect 12404 14662 19870 14714
rect 19922 14662 19934 14714
rect 19986 14662 19998 14714
rect 20050 14662 20062 14714
rect 20114 14662 20126 14714
rect 20178 14662 27644 14714
rect 27696 14662 27708 14714
rect 27760 14662 27772 14714
rect 27824 14662 27836 14714
rect 27888 14662 27900 14714
rect 27952 14662 31648 14714
rect 552 14640 31648 14662
rect 15089 14603 15147 14609
rect 15089 14600 15101 14603
rect 14384 14572 15101 14600
rect 14384 14405 14412 14572
rect 15089 14569 15101 14572
rect 15135 14600 15147 14603
rect 15562 14600 15568 14612
rect 15135 14572 15568 14600
rect 15135 14569 15147 14572
rect 15089 14563 15147 14569
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 16114 14560 16120 14612
rect 16172 14560 16178 14612
rect 16666 14560 16672 14612
rect 16724 14600 16730 14612
rect 17313 14603 17371 14609
rect 17313 14600 17325 14603
rect 16724 14572 17325 14600
rect 16724 14560 16730 14572
rect 17313 14569 17325 14572
rect 17359 14569 17371 14603
rect 17313 14563 17371 14569
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 17865 14603 17923 14609
rect 17865 14600 17877 14603
rect 17828 14572 17877 14600
rect 17828 14560 17834 14572
rect 17865 14569 17877 14572
rect 17911 14569 17923 14603
rect 17865 14563 17923 14569
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 22152 14572 22293 14600
rect 22152 14560 22158 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 25117 14603 25175 14609
rect 25117 14569 25129 14603
rect 25163 14600 25175 14603
rect 25163 14572 25636 14600
rect 25163 14569 25175 14572
rect 25117 14563 25175 14569
rect 15289 14535 15347 14541
rect 15289 14501 15301 14535
rect 15335 14532 15347 14535
rect 15470 14532 15476 14544
rect 15335 14504 15476 14532
rect 15335 14501 15347 14504
rect 15289 14495 15347 14501
rect 15470 14492 15476 14504
rect 15528 14532 15534 14544
rect 15528 14504 17080 14532
rect 15528 14492 15534 14504
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14464 14519 14467
rect 15378 14464 15384 14476
rect 14507 14436 15384 14464
rect 14507 14433 14519 14436
rect 14461 14427 14519 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14464 15623 14467
rect 16482 14464 16488 14476
rect 15611 14436 16488 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16850 14424 16856 14476
rect 16908 14424 16914 14476
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 14369 14359 14427 14365
rect 15028 14368 15485 14396
rect 15028 14272 15056 14368
rect 15473 14365 15485 14368
rect 15519 14365 15531 14399
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 15473 14359 15531 14365
rect 16546 14368 16773 14396
rect 15286 14328 15292 14340
rect 15120 14300 15292 14328
rect 13998 14220 14004 14272
rect 14056 14260 14062 14272
rect 14185 14263 14243 14269
rect 14185 14260 14197 14263
rect 14056 14232 14197 14260
rect 14056 14220 14062 14232
rect 14185 14229 14197 14232
rect 14231 14229 14243 14263
rect 14185 14223 14243 14229
rect 14921 14263 14979 14269
rect 14921 14229 14933 14263
rect 14967 14260 14979 14263
rect 15010 14260 15016 14272
rect 14967 14232 15016 14260
rect 14967 14229 14979 14232
rect 14921 14223 14979 14229
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 15120 14269 15148 14300
rect 15286 14288 15292 14300
rect 15344 14328 15350 14340
rect 16546 14328 16574 14368
rect 16761 14365 16773 14368
rect 16807 14396 16819 14399
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16807 14368 16957 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 15344 14300 16574 14328
rect 15344 14288 15350 14300
rect 15105 14263 15163 14269
rect 15105 14229 15117 14263
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 15841 14263 15899 14269
rect 15841 14229 15853 14263
rect 15887 14260 15899 14263
rect 16390 14260 16396 14272
rect 15887 14232 16396 14260
rect 15887 14229 15899 14232
rect 15841 14223 15899 14229
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 17052 14269 17080 14504
rect 18138 14492 18144 14544
rect 18196 14532 18202 14544
rect 18325 14535 18383 14541
rect 18325 14532 18337 14535
rect 18196 14504 18337 14532
rect 18196 14492 18202 14504
rect 18325 14501 18337 14504
rect 18371 14501 18383 14535
rect 18325 14495 18383 14501
rect 24673 14535 24731 14541
rect 24673 14501 24685 14535
rect 24719 14532 24731 14535
rect 24946 14532 24952 14544
rect 24719 14504 24952 14532
rect 24719 14501 24731 14504
rect 24673 14495 24731 14501
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 25317 14535 25375 14541
rect 25317 14501 25329 14535
rect 25363 14532 25375 14535
rect 25406 14532 25412 14544
rect 25363 14504 25412 14532
rect 25363 14501 25375 14504
rect 25317 14495 25375 14501
rect 25406 14492 25412 14504
rect 25464 14492 25470 14544
rect 25608 14532 25636 14572
rect 25682 14560 25688 14612
rect 25740 14600 25746 14612
rect 25869 14603 25927 14609
rect 25869 14600 25881 14603
rect 25740 14572 25881 14600
rect 25740 14560 25746 14572
rect 25869 14569 25881 14572
rect 25915 14569 25927 14603
rect 25869 14563 25927 14569
rect 26142 14560 26148 14612
rect 26200 14560 26206 14612
rect 25608 14504 26280 14532
rect 26252 14476 26280 14504
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17494 14464 17500 14476
rect 17175 14436 17500 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 18046 14424 18052 14476
rect 18104 14424 18110 14476
rect 19702 14424 19708 14476
rect 19760 14473 19766 14476
rect 19760 14427 19772 14473
rect 20257 14467 20315 14473
rect 20257 14433 20269 14467
rect 20303 14464 20315 14467
rect 21542 14464 21548 14476
rect 20303 14436 21548 14464
rect 20303 14433 20315 14436
rect 20257 14427 20315 14433
rect 19760 14424 19766 14427
rect 21542 14424 21548 14436
rect 21600 14464 21606 14476
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 21600 14436 22385 14464
rect 21600 14424 21606 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 23937 14467 23995 14473
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24026 14464 24032 14476
rect 23983 14436 24032 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24026 14424 24032 14436
rect 24084 14424 24090 14476
rect 24121 14467 24179 14473
rect 24121 14433 24133 14467
rect 24167 14464 24179 14467
rect 24210 14464 24216 14476
rect 24167 14436 24216 14464
rect 24167 14433 24179 14436
rect 24121 14427 24179 14433
rect 24210 14424 24216 14436
rect 24268 14464 24274 14476
rect 24305 14467 24363 14473
rect 24305 14464 24317 14467
rect 24268 14436 24317 14464
rect 24268 14424 24274 14436
rect 24305 14433 24317 14436
rect 24351 14464 24363 14467
rect 24762 14464 24768 14476
rect 24351 14436 24768 14464
rect 24351 14433 24363 14436
rect 24305 14427 24363 14433
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 25958 14424 25964 14476
rect 26016 14424 26022 14476
rect 26234 14424 26240 14476
rect 26292 14424 26298 14476
rect 18230 14356 18236 14408
rect 18288 14396 18294 14408
rect 19981 14399 20039 14405
rect 18288 14368 18644 14396
rect 18288 14356 18294 14368
rect 18616 14337 18644 14368
rect 19981 14365 19993 14399
rect 20027 14396 20039 14399
rect 20165 14399 20223 14405
rect 20165 14396 20177 14399
rect 20027 14368 20177 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 20165 14365 20177 14368
rect 20211 14365 20223 14399
rect 25038 14396 25044 14408
rect 20165 14359 20223 14365
rect 24688 14368 25044 14396
rect 18601 14331 18659 14337
rect 18601 14297 18613 14331
rect 18647 14297 18659 14331
rect 18601 14291 18659 14297
rect 23566 14288 23572 14340
rect 23624 14328 23630 14340
rect 23624 14300 24164 14328
rect 23624 14288 23630 14300
rect 17037 14263 17095 14269
rect 17037 14229 17049 14263
rect 17083 14229 17095 14263
rect 17037 14223 17095 14229
rect 18230 14220 18236 14272
rect 18288 14220 18294 14272
rect 23474 14220 23480 14272
rect 23532 14260 23538 14272
rect 24029 14263 24087 14269
rect 24029 14260 24041 14263
rect 23532 14232 24041 14260
rect 23532 14220 23538 14232
rect 24029 14229 24041 14232
rect 24075 14229 24087 14263
rect 24136 14260 24164 14300
rect 24688 14269 24716 14368
rect 25038 14356 25044 14368
rect 25096 14396 25102 14408
rect 26326 14396 26332 14408
rect 25096 14368 26332 14396
rect 25096 14356 25102 14368
rect 26326 14356 26332 14368
rect 26384 14396 26390 14408
rect 26786 14396 26792 14408
rect 26384 14368 26792 14396
rect 26384 14356 26390 14368
rect 26786 14356 26792 14368
rect 26844 14356 26850 14408
rect 24762 14288 24768 14340
rect 24820 14328 24826 14340
rect 24949 14331 25007 14337
rect 24949 14328 24961 14331
rect 24820 14300 24961 14328
rect 24820 14288 24826 14300
rect 24949 14297 24961 14300
rect 24995 14297 25007 14331
rect 24949 14291 25007 14297
rect 24673 14263 24731 14269
rect 24673 14260 24685 14263
rect 24136 14232 24685 14260
rect 24029 14223 24087 14229
rect 24673 14229 24685 14232
rect 24719 14229 24731 14263
rect 24673 14223 24731 14229
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 25133 14263 25191 14269
rect 25133 14229 25145 14263
rect 25179 14260 25191 14263
rect 25222 14260 25228 14272
rect 25179 14232 25228 14260
rect 25179 14229 25191 14232
rect 25133 14223 25191 14229
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 552 14170 31648 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 11436 14170
rect 11488 14118 11500 14170
rect 11552 14118 11564 14170
rect 11616 14118 11628 14170
rect 11680 14118 11692 14170
rect 11744 14118 19210 14170
rect 19262 14118 19274 14170
rect 19326 14118 19338 14170
rect 19390 14118 19402 14170
rect 19454 14118 19466 14170
rect 19518 14118 26984 14170
rect 27036 14118 27048 14170
rect 27100 14118 27112 14170
rect 27164 14118 27176 14170
rect 27228 14118 27240 14170
rect 27292 14118 31648 14170
rect 552 14096 31648 14118
rect 15286 14016 15292 14068
rect 15344 14016 15350 14068
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14056 19211 14059
rect 19702 14056 19708 14068
rect 19199 14028 19708 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 19702 14016 19708 14028
rect 19760 14016 19766 14068
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 23566 14056 23572 14068
rect 23523 14028 23572 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 23566 14016 23572 14028
rect 23624 14016 23630 14068
rect 24026 14016 24032 14068
rect 24084 14056 24090 14068
rect 24084 14028 24808 14056
rect 24084 14016 24090 14028
rect 15470 13880 15476 13932
rect 15528 13880 15534 13932
rect 17512 13920 17540 14016
rect 18966 13948 18972 14000
rect 19024 13948 19030 14000
rect 24780 13988 24808 14028
rect 24946 14016 24952 14068
rect 25004 14056 25010 14068
rect 25317 14059 25375 14065
rect 25317 14056 25329 14059
rect 25004 14028 25329 14056
rect 25004 14016 25010 14028
rect 25317 14025 25329 14028
rect 25363 14025 25375 14059
rect 25317 14019 25375 14025
rect 25225 13991 25283 13997
rect 25225 13988 25237 13991
rect 24780 13960 25237 13988
rect 25225 13957 25237 13960
rect 25271 13957 25283 13991
rect 25225 13951 25283 13957
rect 25682 13948 25688 14000
rect 25740 13988 25746 14000
rect 25740 13960 27476 13988
rect 25740 13948 25746 13960
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17512 13892 18153 13920
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 18472 13892 18705 13920
rect 18472 13880 18478 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13920 23167 13923
rect 23845 13923 23903 13929
rect 23845 13920 23857 13923
rect 23155 13892 23857 13920
rect 23155 13889 23167 13892
rect 23109 13883 23167 13889
rect 23845 13889 23857 13892
rect 23891 13889 23903 13923
rect 25958 13920 25964 13932
rect 23845 13883 23903 13889
rect 25424 13892 25964 13920
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 13725 13855 13783 13861
rect 13725 13821 13737 13855
rect 13771 13852 13783 13855
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13771 13824 13921 13852
rect 13771 13821 13783 13824
rect 13725 13815 13783 13821
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 13909 13815 13967 13821
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14165 13855 14223 13861
rect 14165 13852 14177 13855
rect 14056 13824 14177 13852
rect 14056 13812 14062 13824
rect 14165 13821 14177 13824
rect 14211 13821 14223 13855
rect 14165 13815 14223 13821
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13852 16175 13855
rect 16666 13852 16672 13864
rect 16163 13824 16672 13852
rect 16163 13821 16175 13824
rect 16117 13815 16175 13821
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 23201 13855 23259 13861
rect 23201 13821 23213 13855
rect 23247 13852 23259 13855
rect 24486 13852 24492 13864
rect 23247 13824 24492 13852
rect 23247 13821 23259 13824
rect 23201 13815 23259 13821
rect 24486 13812 24492 13824
rect 24544 13852 24550 13864
rect 25424 13852 25452 13892
rect 25958 13880 25964 13892
rect 26016 13920 26022 13932
rect 27448 13929 27476 13960
rect 27433 13923 27491 13929
rect 26016 13892 26096 13920
rect 26016 13880 26022 13892
rect 24544 13824 25452 13852
rect 24544 13812 24550 13824
rect 25498 13812 25504 13864
rect 25556 13812 25562 13864
rect 25774 13812 25780 13864
rect 25832 13852 25838 13864
rect 26068 13861 26096 13892
rect 27433 13889 27445 13923
rect 27479 13920 27491 13923
rect 27982 13920 27988 13932
rect 27479 13892 27988 13920
rect 27479 13889 27491 13892
rect 27433 13883 27491 13889
rect 27982 13880 27988 13892
rect 28040 13880 28046 13932
rect 26053 13855 26111 13861
rect 25832 13824 25912 13852
rect 25832 13812 25838 13824
rect 16390 13793 16396 13796
rect 16384 13784 16396 13793
rect 16351 13756 16396 13784
rect 16384 13747 16396 13756
rect 16390 13744 16396 13747
rect 16448 13744 16454 13796
rect 23290 13744 23296 13796
rect 23348 13744 23354 13796
rect 23474 13744 23480 13796
rect 23532 13793 23538 13796
rect 23532 13787 23551 13793
rect 23539 13753 23551 13787
rect 24090 13787 24148 13793
rect 24090 13784 24102 13787
rect 23532 13747 23551 13753
rect 23676 13756 24102 13784
rect 23532 13744 23538 13747
rect 16022 13676 16028 13728
rect 16080 13676 16086 13728
rect 17586 13676 17592 13728
rect 17644 13676 17650 13728
rect 23676 13725 23704 13756
rect 24090 13753 24102 13756
rect 24136 13753 24148 13787
rect 24090 13747 24148 13753
rect 25222 13744 25228 13796
rect 25280 13784 25286 13796
rect 25682 13784 25688 13796
rect 25280 13756 25688 13784
rect 25280 13744 25286 13756
rect 25682 13744 25688 13756
rect 25740 13744 25746 13796
rect 25884 13784 25912 13824
rect 26053 13821 26065 13855
rect 26099 13852 26111 13855
rect 26697 13855 26755 13861
rect 26697 13852 26709 13855
rect 26099 13824 26709 13852
rect 26099 13821 26111 13824
rect 26053 13815 26111 13821
rect 26697 13821 26709 13824
rect 26743 13821 26755 13855
rect 26697 13815 26755 13821
rect 26142 13784 26148 13796
rect 25884 13756 26148 13784
rect 26142 13744 26148 13756
rect 26200 13744 26206 13796
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 26881 13787 26939 13793
rect 26881 13784 26893 13787
rect 26292 13756 26893 13784
rect 26292 13744 26298 13756
rect 26881 13753 26893 13756
rect 26927 13753 26939 13787
rect 26881 13747 26939 13753
rect 23661 13719 23719 13725
rect 23661 13685 23673 13719
rect 23707 13685 23719 13719
rect 23661 13679 23719 13685
rect 25866 13676 25872 13728
rect 25924 13716 25930 13728
rect 25961 13719 26019 13725
rect 25961 13716 25973 13719
rect 25924 13688 25973 13716
rect 25924 13676 25930 13688
rect 25961 13685 25973 13688
rect 26007 13685 26019 13719
rect 25961 13679 26019 13685
rect 26418 13676 26424 13728
rect 26476 13716 26482 13728
rect 26605 13719 26663 13725
rect 26605 13716 26617 13719
rect 26476 13688 26617 13716
rect 26476 13676 26482 13688
rect 26605 13685 26617 13688
rect 26651 13685 26663 13719
rect 26605 13679 26663 13685
rect 552 13626 31648 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 12096 13626
rect 12148 13574 12160 13626
rect 12212 13574 12224 13626
rect 12276 13574 12288 13626
rect 12340 13574 12352 13626
rect 12404 13574 19870 13626
rect 19922 13574 19934 13626
rect 19986 13574 19998 13626
rect 20050 13574 20062 13626
rect 20114 13574 20126 13626
rect 20178 13574 27644 13626
rect 27696 13574 27708 13626
rect 27760 13574 27772 13626
rect 27824 13574 27836 13626
rect 27888 13574 27900 13626
rect 27952 13574 31648 13626
rect 552 13552 31648 13574
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 15344 13484 15761 13512
rect 15344 13472 15350 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16540 13484 16957 13512
rect 16540 13472 16546 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 16945 13475 17003 13481
rect 18417 13515 18475 13521
rect 18417 13481 18429 13515
rect 18463 13512 18475 13515
rect 18506 13512 18512 13524
rect 18463 13484 18512 13512
rect 18463 13481 18475 13484
rect 18417 13475 18475 13481
rect 15933 13447 15991 13453
rect 15933 13413 15945 13447
rect 15979 13444 15991 13447
rect 16022 13444 16028 13456
rect 15979 13416 16028 13444
rect 15979 13413 15991 13416
rect 15933 13407 15991 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 14182 13336 14188 13388
rect 14240 13336 14246 13388
rect 14452 13379 14510 13385
rect 14452 13345 14464 13379
rect 14498 13376 14510 13379
rect 14918 13376 14924 13388
rect 14498 13348 14924 13376
rect 14498 13345 14510 13348
rect 14452 13339 14510 13345
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15620 13348 15669 13376
rect 15620 13336 15626 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13376 17095 13379
rect 17586 13376 17592 13388
rect 17083 13348 17592 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13376 17923 13379
rect 18432 13376 18460 13475
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23845 13515 23903 13521
rect 23845 13512 23857 13515
rect 23348 13484 23857 13512
rect 23348 13472 23354 13484
rect 23845 13481 23857 13484
rect 23891 13481 23903 13515
rect 23845 13475 23903 13481
rect 24305 13515 24363 13521
rect 24305 13481 24317 13515
rect 24351 13512 24363 13515
rect 25498 13512 25504 13524
rect 24351 13484 25504 13512
rect 24351 13481 24363 13484
rect 24305 13475 24363 13481
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 27801 13515 27859 13521
rect 27801 13481 27813 13515
rect 27847 13512 27859 13515
rect 27982 13512 27988 13524
rect 27847 13484 27988 13512
rect 27847 13481 27859 13484
rect 27801 13475 27859 13481
rect 27982 13472 27988 13484
rect 28040 13472 28046 13524
rect 24026 13404 24032 13456
rect 24084 13404 24090 13456
rect 24210 13404 24216 13456
rect 24268 13404 24274 13456
rect 24854 13404 24860 13456
rect 24912 13444 24918 13456
rect 25418 13447 25476 13453
rect 25418 13444 25430 13447
rect 24912 13416 25430 13444
rect 24912 13404 24918 13416
rect 25418 13413 25430 13416
rect 25464 13413 25476 13447
rect 25418 13407 25476 13413
rect 17911 13348 18460 13376
rect 18509 13379 18567 13385
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 18509 13345 18521 13379
rect 18555 13376 18567 13379
rect 18969 13379 19027 13385
rect 18969 13376 18981 13379
rect 18555 13348 18981 13376
rect 18555 13345 18567 13348
rect 18509 13339 18567 13345
rect 18969 13345 18981 13348
rect 19015 13345 19027 13379
rect 18969 13339 19027 13345
rect 25774 13336 25780 13388
rect 25832 13336 25838 13388
rect 25961 13379 26019 13385
rect 25961 13345 25973 13379
rect 26007 13376 26019 13379
rect 26234 13376 26240 13388
rect 26007 13348 26240 13376
rect 26007 13345 26019 13348
rect 25961 13339 26019 13345
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 26418 13336 26424 13388
rect 26476 13336 26482 13388
rect 26510 13336 26516 13388
rect 26568 13376 26574 13388
rect 26677 13379 26735 13385
rect 26677 13376 26689 13379
rect 26568 13348 26689 13376
rect 26568 13336 26574 13348
rect 26677 13345 26689 13348
rect 26723 13345 26735 13379
rect 26677 13339 26735 13345
rect 16669 13311 16727 13317
rect 16669 13308 16681 13311
rect 16546 13280 16681 13308
rect 15470 13200 15476 13252
rect 15528 13240 15534 13252
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 15528 13212 15577 13240
rect 15528 13200 15534 13212
rect 15565 13209 15577 13212
rect 15611 13209 15623 13243
rect 15565 13203 15623 13209
rect 15933 13243 15991 13249
rect 15933 13209 15945 13243
rect 15979 13240 15991 13243
rect 16546 13240 16574 13280
rect 16669 13277 16681 13280
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18414 13308 18420 13320
rect 18003 13280 18420 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 25685 13311 25743 13317
rect 25685 13277 25697 13311
rect 25731 13308 25743 13311
rect 25866 13308 25872 13320
rect 25731 13280 25872 13308
rect 25731 13277 25743 13280
rect 25685 13271 25743 13277
rect 15979 13212 16574 13240
rect 18233 13243 18291 13249
rect 15979 13209 15991 13212
rect 15933 13203 15991 13209
rect 18233 13209 18245 13243
rect 18279 13240 18291 13243
rect 18506 13240 18512 13252
rect 18279 13212 18512 13240
rect 18279 13209 18291 13212
rect 18233 13203 18291 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 19536 13240 19564 13271
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 19024 13212 19564 13240
rect 19024 13200 19030 13212
rect 16114 13132 16120 13184
rect 16172 13132 16178 13184
rect 25774 13132 25780 13184
rect 25832 13172 25838 13184
rect 25869 13175 25927 13181
rect 25869 13172 25881 13175
rect 25832 13144 25881 13172
rect 25832 13132 25838 13144
rect 25869 13141 25881 13144
rect 25915 13141 25927 13175
rect 25869 13135 25927 13141
rect 552 13082 31648 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 11436 13082
rect 11488 13030 11500 13082
rect 11552 13030 11564 13082
rect 11616 13030 11628 13082
rect 11680 13030 11692 13082
rect 11744 13030 19210 13082
rect 19262 13030 19274 13082
rect 19326 13030 19338 13082
rect 19390 13030 19402 13082
rect 19454 13030 19466 13082
rect 19518 13030 26984 13082
rect 27036 13030 27048 13082
rect 27100 13030 27112 13082
rect 27164 13030 27176 13082
rect 27228 13030 27240 13082
rect 27292 13030 31648 13082
rect 552 13008 31648 13030
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 14976 12940 15117 12968
rect 14976 12928 14982 12940
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 15105 12931 15163 12937
rect 16666 12928 16672 12980
rect 16724 12928 16730 12980
rect 26237 12971 26295 12977
rect 26237 12937 26249 12971
rect 26283 12968 26295 12971
rect 26510 12968 26516 12980
rect 26283 12940 26516 12968
rect 26283 12937 26295 12940
rect 26237 12931 26295 12937
rect 26510 12928 26516 12940
rect 26568 12928 26574 12980
rect 18049 12903 18107 12909
rect 18049 12900 18061 12903
rect 17972 12872 18061 12900
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16850 12832 16856 12844
rect 16531 12804 16856 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 17972 12841 18000 12872
rect 18049 12869 18061 12872
rect 18095 12869 18107 12903
rect 26326 12900 26332 12912
rect 18049 12863 18107 12869
rect 25608 12872 26332 12900
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12801 18015 12835
rect 17957 12795 18015 12801
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 15010 12764 15016 12776
rect 14967 12736 15016 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 15105 12767 15163 12773
rect 15105 12733 15117 12767
rect 15151 12764 15163 12767
rect 16114 12764 16120 12776
rect 15151 12736 16120 12764
rect 15151 12733 15163 12736
rect 15105 12727 15163 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16347 12736 16528 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16500 12708 16528 12736
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 16632 12736 16773 12764
rect 16632 12724 16638 12736
rect 16761 12733 16773 12736
rect 16807 12733 16819 12767
rect 16761 12727 16819 12733
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 17267 12736 17325 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 16482 12656 16488 12708
rect 16540 12696 16546 12708
rect 17052 12696 17080 12727
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 17552 12736 18337 12764
rect 17552 12724 17558 12736
rect 18325 12733 18337 12736
rect 18371 12764 18383 12767
rect 18414 12764 18420 12776
rect 18371 12736 18420 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18874 12724 18880 12776
rect 18932 12724 18938 12776
rect 25608 12773 25636 12872
rect 26326 12860 26332 12872
rect 26384 12860 26390 12912
rect 25682 12792 25688 12844
rect 25740 12832 25746 12844
rect 25740 12804 25912 12832
rect 25740 12792 25746 12804
rect 25593 12767 25651 12773
rect 25593 12733 25605 12767
rect 25639 12733 25651 12767
rect 25593 12727 25651 12733
rect 25774 12724 25780 12776
rect 25832 12724 25838 12776
rect 25884 12773 25912 12804
rect 25869 12767 25927 12773
rect 25869 12733 25881 12767
rect 25915 12733 25927 12767
rect 25869 12727 25927 12733
rect 25961 12767 26019 12773
rect 25961 12733 25973 12767
rect 26007 12733 26019 12767
rect 25961 12727 26019 12733
rect 16540 12668 17080 12696
rect 16540 12656 16546 12668
rect 18046 12656 18052 12708
rect 18104 12656 18110 12708
rect 25222 12656 25228 12708
rect 25280 12696 25286 12708
rect 25976 12696 26004 12727
rect 25280 12668 26004 12696
rect 25280 12656 25286 12668
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15620 12600 16129 12628
rect 15620 12588 15626 12600
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 16117 12591 16175 12597
rect 17126 12588 17132 12640
rect 17184 12588 17190 12640
rect 18230 12588 18236 12640
rect 18288 12588 18294 12640
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 18785 12631 18843 12637
rect 18785 12628 18797 12631
rect 18380 12600 18797 12628
rect 18380 12588 18386 12600
rect 18785 12597 18797 12600
rect 18831 12597 18843 12631
rect 18785 12591 18843 12597
rect 552 12538 31648 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 12096 12538
rect 12148 12486 12160 12538
rect 12212 12486 12224 12538
rect 12276 12486 12288 12538
rect 12340 12486 12352 12538
rect 12404 12486 19870 12538
rect 19922 12486 19934 12538
rect 19986 12486 19998 12538
rect 20050 12486 20062 12538
rect 20114 12486 20126 12538
rect 20178 12486 27644 12538
rect 27696 12486 27708 12538
rect 27760 12486 27772 12538
rect 27824 12486 27836 12538
rect 27888 12486 27900 12538
rect 27952 12486 31648 12538
rect 552 12464 31648 12486
rect 16482 12424 16488 12436
rect 15764 12396 16488 12424
rect 15764 12297 15792 12396
rect 16482 12384 16488 12396
rect 16540 12424 16546 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 16540 12396 17049 12424
rect 16540 12384 16546 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 17037 12387 17095 12393
rect 17205 12427 17263 12433
rect 17205 12393 17217 12427
rect 17251 12424 17263 12427
rect 17494 12424 17500 12436
rect 17251 12396 17500 12424
rect 17251 12393 17263 12396
rect 17205 12387 17263 12393
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 18104 12396 18153 12424
rect 18104 12384 18110 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18141 12387 18199 12393
rect 18506 12365 18512 12368
rect 17405 12359 17463 12365
rect 17405 12325 17417 12359
rect 17451 12325 17463 12359
rect 18500 12356 18512 12365
rect 18467 12328 18512 12356
rect 17405 12319 17463 12325
rect 18500 12319 18512 12328
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 15979 12260 16313 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 16850 12248 16856 12300
rect 16908 12248 16914 12300
rect 17420 12288 17448 12319
rect 18506 12316 18512 12319
rect 18564 12316 18570 12368
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 17420 12260 17601 12288
rect 17589 12257 17601 12260
rect 17635 12288 17647 12291
rect 17954 12288 17960 12300
rect 17635 12260 17960 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 18322 12288 18328 12300
rect 18279 12260 18328 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 15746 12044 15752 12096
rect 15804 12044 15810 12096
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 18230 12084 18236 12096
rect 17267 12056 18236 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 18230 12044 18236 12056
rect 18288 12084 18294 12096
rect 18966 12084 18972 12096
rect 18288 12056 18972 12084
rect 18288 12044 18294 12056
rect 18966 12044 18972 12056
rect 19024 12084 19030 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19024 12056 19625 12084
rect 19024 12044 19030 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 552 11994 31648 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 11436 11994
rect 11488 11942 11500 11994
rect 11552 11942 11564 11994
rect 11616 11942 11628 11994
rect 11680 11942 11692 11994
rect 11744 11942 19210 11994
rect 19262 11942 19274 11994
rect 19326 11942 19338 11994
rect 19390 11942 19402 11994
rect 19454 11942 19466 11994
rect 19518 11942 26984 11994
rect 27036 11942 27048 11994
rect 27100 11942 27112 11994
rect 27164 11942 27176 11994
rect 27228 11942 27240 11994
rect 27292 11942 31648 11994
rect 552 11920 31648 11942
rect 16574 11880 16580 11892
rect 14936 11852 16580 11880
rect 14936 11685 14964 11852
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18233 11883 18291 11889
rect 18233 11880 18245 11883
rect 18012 11852 18245 11880
rect 18012 11840 18018 11852
rect 18233 11849 18245 11852
rect 18279 11849 18291 11883
rect 18233 11843 18291 11849
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 15059 11648 15209 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15197 11645 15209 11648
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 16850 11636 16856 11688
rect 16908 11636 16914 11688
rect 17126 11685 17132 11688
rect 17120 11676 17132 11685
rect 17087 11648 17132 11676
rect 17120 11639 17132 11648
rect 17126 11636 17132 11639
rect 17184 11636 17190 11688
rect 15464 11611 15522 11617
rect 15464 11577 15476 11611
rect 15510 11608 15522 11611
rect 15654 11608 15660 11620
rect 15510 11580 15660 11608
rect 15510 11577 15522 11580
rect 15464 11571 15522 11577
rect 15654 11568 15660 11580
rect 15712 11568 15718 11620
rect 16577 11543 16635 11549
rect 16577 11509 16589 11543
rect 16623 11540 16635 11543
rect 16758 11540 16764 11552
rect 16623 11512 16764 11540
rect 16623 11509 16635 11512
rect 16577 11503 16635 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 552 11450 31648 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 12096 11450
rect 12148 11398 12160 11450
rect 12212 11398 12224 11450
rect 12276 11398 12288 11450
rect 12340 11398 12352 11450
rect 12404 11398 19870 11450
rect 19922 11398 19934 11450
rect 19986 11398 19998 11450
rect 20050 11398 20062 11450
rect 20114 11398 20126 11450
rect 20178 11398 27644 11450
rect 27696 11398 27708 11450
rect 27760 11398 27772 11450
rect 27824 11398 27836 11450
rect 27888 11398 27900 11450
rect 27952 11398 31648 11450
rect 552 11376 31648 11398
rect 15654 11296 15660 11348
rect 15712 11296 15718 11348
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 17037 11339 17095 11345
rect 17037 11336 17049 11339
rect 16908 11308 17049 11336
rect 16908 11296 16914 11308
rect 17037 11305 17049 11308
rect 17083 11305 17095 11339
rect 17037 11299 17095 11305
rect 15562 11160 15568 11212
rect 15620 11160 15626 11212
rect 15746 11160 15752 11212
rect 15804 11160 15810 11212
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 18874 11200 18880 11212
rect 17175 11172 18880 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 18874 11160 18880 11172
rect 18932 11160 18938 11212
rect 552 10906 31648 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 11436 10906
rect 11488 10854 11500 10906
rect 11552 10854 11564 10906
rect 11616 10854 11628 10906
rect 11680 10854 11692 10906
rect 11744 10854 19210 10906
rect 19262 10854 19274 10906
rect 19326 10854 19338 10906
rect 19390 10854 19402 10906
rect 19454 10854 19466 10906
rect 19518 10854 26984 10906
rect 27036 10854 27048 10906
rect 27100 10854 27112 10906
rect 27164 10854 27176 10906
rect 27228 10854 27240 10906
rect 27292 10854 31648 10906
rect 552 10832 31648 10854
rect 552 10362 31648 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 12096 10362
rect 12148 10310 12160 10362
rect 12212 10310 12224 10362
rect 12276 10310 12288 10362
rect 12340 10310 12352 10362
rect 12404 10310 19870 10362
rect 19922 10310 19934 10362
rect 19986 10310 19998 10362
rect 20050 10310 20062 10362
rect 20114 10310 20126 10362
rect 20178 10310 27644 10362
rect 27696 10310 27708 10362
rect 27760 10310 27772 10362
rect 27824 10310 27836 10362
rect 27888 10310 27900 10362
rect 27952 10310 31648 10362
rect 552 10288 31648 10310
rect 552 9818 31648 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 11436 9818
rect 11488 9766 11500 9818
rect 11552 9766 11564 9818
rect 11616 9766 11628 9818
rect 11680 9766 11692 9818
rect 11744 9766 19210 9818
rect 19262 9766 19274 9818
rect 19326 9766 19338 9818
rect 19390 9766 19402 9818
rect 19454 9766 19466 9818
rect 19518 9766 26984 9818
rect 27036 9766 27048 9818
rect 27100 9766 27112 9818
rect 27164 9766 27176 9818
rect 27228 9766 27240 9818
rect 27292 9766 31648 9818
rect 552 9744 31648 9766
rect 552 9274 31648 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 12096 9274
rect 12148 9222 12160 9274
rect 12212 9222 12224 9274
rect 12276 9222 12288 9274
rect 12340 9222 12352 9274
rect 12404 9222 19870 9274
rect 19922 9222 19934 9274
rect 19986 9222 19998 9274
rect 20050 9222 20062 9274
rect 20114 9222 20126 9274
rect 20178 9222 27644 9274
rect 27696 9222 27708 9274
rect 27760 9222 27772 9274
rect 27824 9222 27836 9274
rect 27888 9222 27900 9274
rect 27952 9222 31648 9274
rect 552 9200 31648 9222
rect 552 8730 31648 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 11436 8730
rect 11488 8678 11500 8730
rect 11552 8678 11564 8730
rect 11616 8678 11628 8730
rect 11680 8678 11692 8730
rect 11744 8678 19210 8730
rect 19262 8678 19274 8730
rect 19326 8678 19338 8730
rect 19390 8678 19402 8730
rect 19454 8678 19466 8730
rect 19518 8678 26984 8730
rect 27036 8678 27048 8730
rect 27100 8678 27112 8730
rect 27164 8678 27176 8730
rect 27228 8678 27240 8730
rect 27292 8678 31648 8730
rect 552 8656 31648 8678
rect 552 8186 31648 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 12096 8186
rect 12148 8134 12160 8186
rect 12212 8134 12224 8186
rect 12276 8134 12288 8186
rect 12340 8134 12352 8186
rect 12404 8134 19870 8186
rect 19922 8134 19934 8186
rect 19986 8134 19998 8186
rect 20050 8134 20062 8186
rect 20114 8134 20126 8186
rect 20178 8134 27644 8186
rect 27696 8134 27708 8186
rect 27760 8134 27772 8186
rect 27824 8134 27836 8186
rect 27888 8134 27900 8186
rect 27952 8134 31648 8186
rect 552 8112 31648 8134
rect 552 7642 31648 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 11436 7642
rect 11488 7590 11500 7642
rect 11552 7590 11564 7642
rect 11616 7590 11628 7642
rect 11680 7590 11692 7642
rect 11744 7590 19210 7642
rect 19262 7590 19274 7642
rect 19326 7590 19338 7642
rect 19390 7590 19402 7642
rect 19454 7590 19466 7642
rect 19518 7590 26984 7642
rect 27036 7590 27048 7642
rect 27100 7590 27112 7642
rect 27164 7590 27176 7642
rect 27228 7590 27240 7642
rect 27292 7590 31648 7642
rect 552 7568 31648 7590
rect 552 7098 31648 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 12096 7098
rect 12148 7046 12160 7098
rect 12212 7046 12224 7098
rect 12276 7046 12288 7098
rect 12340 7046 12352 7098
rect 12404 7046 19870 7098
rect 19922 7046 19934 7098
rect 19986 7046 19998 7098
rect 20050 7046 20062 7098
rect 20114 7046 20126 7098
rect 20178 7046 27644 7098
rect 27696 7046 27708 7098
rect 27760 7046 27772 7098
rect 27824 7046 27836 7098
rect 27888 7046 27900 7098
rect 27952 7046 31648 7098
rect 552 7024 31648 7046
rect 552 6554 31648 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 11436 6554
rect 11488 6502 11500 6554
rect 11552 6502 11564 6554
rect 11616 6502 11628 6554
rect 11680 6502 11692 6554
rect 11744 6502 19210 6554
rect 19262 6502 19274 6554
rect 19326 6502 19338 6554
rect 19390 6502 19402 6554
rect 19454 6502 19466 6554
rect 19518 6502 26984 6554
rect 27036 6502 27048 6554
rect 27100 6502 27112 6554
rect 27164 6502 27176 6554
rect 27228 6502 27240 6554
rect 27292 6502 31648 6554
rect 552 6480 31648 6502
rect 552 6010 31648 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 12096 6010
rect 12148 5958 12160 6010
rect 12212 5958 12224 6010
rect 12276 5958 12288 6010
rect 12340 5958 12352 6010
rect 12404 5958 19870 6010
rect 19922 5958 19934 6010
rect 19986 5958 19998 6010
rect 20050 5958 20062 6010
rect 20114 5958 20126 6010
rect 20178 5958 27644 6010
rect 27696 5958 27708 6010
rect 27760 5958 27772 6010
rect 27824 5958 27836 6010
rect 27888 5958 27900 6010
rect 27952 5958 31648 6010
rect 552 5936 31648 5958
rect 552 5466 31648 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 11436 5466
rect 11488 5414 11500 5466
rect 11552 5414 11564 5466
rect 11616 5414 11628 5466
rect 11680 5414 11692 5466
rect 11744 5414 19210 5466
rect 19262 5414 19274 5466
rect 19326 5414 19338 5466
rect 19390 5414 19402 5466
rect 19454 5414 19466 5466
rect 19518 5414 26984 5466
rect 27036 5414 27048 5466
rect 27100 5414 27112 5466
rect 27164 5414 27176 5466
rect 27228 5414 27240 5466
rect 27292 5414 31648 5466
rect 552 5392 31648 5414
rect 552 4922 31648 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 12096 4922
rect 12148 4870 12160 4922
rect 12212 4870 12224 4922
rect 12276 4870 12288 4922
rect 12340 4870 12352 4922
rect 12404 4870 19870 4922
rect 19922 4870 19934 4922
rect 19986 4870 19998 4922
rect 20050 4870 20062 4922
rect 20114 4870 20126 4922
rect 20178 4870 27644 4922
rect 27696 4870 27708 4922
rect 27760 4870 27772 4922
rect 27824 4870 27836 4922
rect 27888 4870 27900 4922
rect 27952 4870 31648 4922
rect 552 4848 31648 4870
rect 552 4378 31648 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 11436 4378
rect 11488 4326 11500 4378
rect 11552 4326 11564 4378
rect 11616 4326 11628 4378
rect 11680 4326 11692 4378
rect 11744 4326 19210 4378
rect 19262 4326 19274 4378
rect 19326 4326 19338 4378
rect 19390 4326 19402 4378
rect 19454 4326 19466 4378
rect 19518 4326 26984 4378
rect 27036 4326 27048 4378
rect 27100 4326 27112 4378
rect 27164 4326 27176 4378
rect 27228 4326 27240 4378
rect 27292 4326 31648 4378
rect 552 4304 31648 4326
rect 552 3834 31648 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 12096 3834
rect 12148 3782 12160 3834
rect 12212 3782 12224 3834
rect 12276 3782 12288 3834
rect 12340 3782 12352 3834
rect 12404 3782 19870 3834
rect 19922 3782 19934 3834
rect 19986 3782 19998 3834
rect 20050 3782 20062 3834
rect 20114 3782 20126 3834
rect 20178 3782 27644 3834
rect 27696 3782 27708 3834
rect 27760 3782 27772 3834
rect 27824 3782 27836 3834
rect 27888 3782 27900 3834
rect 27952 3782 31648 3834
rect 552 3760 31648 3782
rect 552 3290 31648 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 11436 3290
rect 11488 3238 11500 3290
rect 11552 3238 11564 3290
rect 11616 3238 11628 3290
rect 11680 3238 11692 3290
rect 11744 3238 19210 3290
rect 19262 3238 19274 3290
rect 19326 3238 19338 3290
rect 19390 3238 19402 3290
rect 19454 3238 19466 3290
rect 19518 3238 26984 3290
rect 27036 3238 27048 3290
rect 27100 3238 27112 3290
rect 27164 3238 27176 3290
rect 27228 3238 27240 3290
rect 27292 3238 31648 3290
rect 552 3216 31648 3238
rect 552 2746 31648 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 12096 2746
rect 12148 2694 12160 2746
rect 12212 2694 12224 2746
rect 12276 2694 12288 2746
rect 12340 2694 12352 2746
rect 12404 2694 19870 2746
rect 19922 2694 19934 2746
rect 19986 2694 19998 2746
rect 20050 2694 20062 2746
rect 20114 2694 20126 2746
rect 20178 2694 27644 2746
rect 27696 2694 27708 2746
rect 27760 2694 27772 2746
rect 27824 2694 27836 2746
rect 27888 2694 27900 2746
rect 27952 2694 31648 2746
rect 552 2672 31648 2694
rect 552 2202 31648 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 11436 2202
rect 11488 2150 11500 2202
rect 11552 2150 11564 2202
rect 11616 2150 11628 2202
rect 11680 2150 11692 2202
rect 11744 2150 19210 2202
rect 19262 2150 19274 2202
rect 19326 2150 19338 2202
rect 19390 2150 19402 2202
rect 19454 2150 19466 2202
rect 19518 2150 26984 2202
rect 27036 2150 27048 2202
rect 27100 2150 27112 2202
rect 27164 2150 27176 2202
rect 27228 2150 27240 2202
rect 27292 2150 31648 2202
rect 552 2128 31648 2150
rect 552 1658 31648 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 12096 1658
rect 12148 1606 12160 1658
rect 12212 1606 12224 1658
rect 12276 1606 12288 1658
rect 12340 1606 12352 1658
rect 12404 1606 19870 1658
rect 19922 1606 19934 1658
rect 19986 1606 19998 1658
rect 20050 1606 20062 1658
rect 20114 1606 20126 1658
rect 20178 1606 27644 1658
rect 27696 1606 27708 1658
rect 27760 1606 27772 1658
rect 27824 1606 27836 1658
rect 27888 1606 27900 1658
rect 27952 1606 31648 1658
rect 552 1584 31648 1606
rect 552 1114 31648 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 11436 1114
rect 11488 1062 11500 1114
rect 11552 1062 11564 1114
rect 11616 1062 11628 1114
rect 11680 1062 11692 1114
rect 11744 1062 19210 1114
rect 19262 1062 19274 1114
rect 19326 1062 19338 1114
rect 19390 1062 19402 1114
rect 19454 1062 19466 1114
rect 19518 1062 26984 1114
rect 27036 1062 27048 1114
rect 27100 1062 27112 1114
rect 27164 1062 27176 1114
rect 27228 1062 27240 1114
rect 27292 1062 31648 1114
rect 552 1040 31648 1062
rect 552 570 31648 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 12096 570
rect 12148 518 12160 570
rect 12212 518 12224 570
rect 12276 518 12288 570
rect 12340 518 12352 570
rect 12404 518 19870 570
rect 19922 518 19934 570
rect 19986 518 19998 570
rect 20050 518 20062 570
rect 20114 518 20126 570
rect 20178 518 27644 570
rect 27696 518 27708 570
rect 27760 518 27772 570
rect 27824 518 27836 570
rect 27888 518 27900 570
rect 27952 518 31648 570
rect 552 496 31648 518
<< via1 >>
rect 3662 44582 3714 44634
rect 3726 44582 3778 44634
rect 3790 44582 3842 44634
rect 3854 44582 3906 44634
rect 3918 44582 3970 44634
rect 11436 44582 11488 44634
rect 11500 44582 11552 44634
rect 11564 44582 11616 44634
rect 11628 44582 11680 44634
rect 11692 44582 11744 44634
rect 19210 44582 19262 44634
rect 19274 44582 19326 44634
rect 19338 44582 19390 44634
rect 19402 44582 19454 44634
rect 19466 44582 19518 44634
rect 26984 44582 27036 44634
rect 27048 44582 27100 44634
rect 27112 44582 27164 44634
rect 27176 44582 27228 44634
rect 27240 44582 27292 44634
rect 7196 44523 7248 44532
rect 7196 44489 7205 44523
rect 7205 44489 7239 44523
rect 7239 44489 7248 44523
rect 7196 44480 7248 44489
rect 7656 44523 7708 44532
rect 7656 44489 7665 44523
rect 7665 44489 7699 44523
rect 7699 44489 7708 44523
rect 7656 44480 7708 44489
rect 8300 44480 8352 44532
rect 8760 44523 8812 44532
rect 8760 44489 8769 44523
rect 8769 44489 8803 44523
rect 8803 44489 8812 44523
rect 8760 44480 8812 44489
rect 9312 44523 9364 44532
rect 9312 44489 9321 44523
rect 9321 44489 9355 44523
rect 9355 44489 9364 44523
rect 9312 44480 9364 44489
rect 11796 44480 11848 44532
rect 12808 44523 12860 44532
rect 12808 44489 12817 44523
rect 12817 44489 12851 44523
rect 12851 44489 12860 44523
rect 12808 44480 12860 44489
rect 13084 44523 13136 44532
rect 13084 44489 13093 44523
rect 13093 44489 13127 44523
rect 13127 44489 13136 44523
rect 13084 44480 13136 44489
rect 27436 44480 27488 44532
rect 25228 44412 25280 44464
rect 11888 44344 11940 44396
rect 8208 44276 8260 44328
rect 11060 44208 11112 44260
rect 13728 44319 13780 44328
rect 13728 44285 13737 44319
rect 13737 44285 13771 44319
rect 13771 44285 13780 44319
rect 13728 44276 13780 44285
rect 13820 44319 13872 44328
rect 13820 44285 13829 44319
rect 13829 44285 13863 44319
rect 13863 44285 13872 44319
rect 13820 44276 13872 44285
rect 14004 44319 14056 44328
rect 14004 44285 14013 44319
rect 14013 44285 14047 44319
rect 14047 44285 14056 44319
rect 14004 44276 14056 44285
rect 15844 44276 15896 44328
rect 16488 44276 16540 44328
rect 21640 44319 21692 44328
rect 21640 44285 21649 44319
rect 21649 44285 21683 44319
rect 21683 44285 21692 44319
rect 21640 44276 21692 44285
rect 24032 44319 24084 44328
rect 24032 44285 24041 44319
rect 24041 44285 24075 44319
rect 24075 44285 24084 44319
rect 24032 44276 24084 44285
rect 24400 44319 24452 44328
rect 24400 44285 24409 44319
rect 24409 44285 24443 44319
rect 24443 44285 24452 44319
rect 24400 44276 24452 44285
rect 24952 44319 25004 44328
rect 24952 44285 24961 44319
rect 24961 44285 24995 44319
rect 24995 44285 25004 44319
rect 24952 44276 25004 44285
rect 25504 44319 25556 44328
rect 25504 44285 25513 44319
rect 25513 44285 25547 44319
rect 25547 44285 25556 44319
rect 25504 44276 25556 44285
rect 26516 44344 26568 44396
rect 26056 44319 26108 44328
rect 26056 44285 26065 44319
rect 26065 44285 26099 44319
rect 26099 44285 26108 44319
rect 26056 44276 26108 44285
rect 29000 44387 29052 44396
rect 29000 44353 29009 44387
rect 29009 44353 29043 44387
rect 29043 44353 29052 44387
rect 29000 44344 29052 44353
rect 28172 44319 28224 44328
rect 28172 44285 28181 44319
rect 28181 44285 28215 44319
rect 28215 44285 28224 44319
rect 28172 44276 28224 44285
rect 29276 44319 29328 44328
rect 29276 44285 29285 44319
rect 29285 44285 29319 44319
rect 29319 44285 29328 44319
rect 29276 44276 29328 44285
rect 8300 44140 8352 44192
rect 12440 44140 12492 44192
rect 12532 44183 12584 44192
rect 12532 44149 12541 44183
rect 12541 44149 12575 44183
rect 12575 44149 12584 44183
rect 12532 44140 12584 44149
rect 13544 44183 13596 44192
rect 13544 44149 13553 44183
rect 13553 44149 13587 44183
rect 13587 44149 13596 44183
rect 13544 44140 13596 44149
rect 14280 44140 14332 44192
rect 15752 44140 15804 44192
rect 16764 44140 16816 44192
rect 19248 44140 19300 44192
rect 21824 44183 21876 44192
rect 21824 44149 21833 44183
rect 21833 44149 21867 44183
rect 21867 44149 21876 44183
rect 21824 44140 21876 44149
rect 22008 44140 22060 44192
rect 24584 44183 24636 44192
rect 24584 44149 24593 44183
rect 24593 44149 24627 44183
rect 24627 44149 24636 44183
rect 24584 44140 24636 44149
rect 25136 44183 25188 44192
rect 25136 44149 25145 44183
rect 25145 44149 25179 44183
rect 25179 44149 25188 44183
rect 25136 44140 25188 44149
rect 25688 44183 25740 44192
rect 25688 44149 25697 44183
rect 25697 44149 25731 44183
rect 25731 44149 25740 44183
rect 25688 44140 25740 44149
rect 26240 44183 26292 44192
rect 26240 44149 26249 44183
rect 26249 44149 26283 44183
rect 26283 44149 26292 44183
rect 26240 44140 26292 44149
rect 27436 44208 27488 44260
rect 28080 44183 28132 44192
rect 28080 44149 28089 44183
rect 28089 44149 28123 44183
rect 28123 44149 28132 44183
rect 28080 44140 28132 44149
rect 29000 44140 29052 44192
rect 4322 44038 4374 44090
rect 4386 44038 4438 44090
rect 4450 44038 4502 44090
rect 4514 44038 4566 44090
rect 4578 44038 4630 44090
rect 12096 44038 12148 44090
rect 12160 44038 12212 44090
rect 12224 44038 12276 44090
rect 12288 44038 12340 44090
rect 12352 44038 12404 44090
rect 19870 44038 19922 44090
rect 19934 44038 19986 44090
rect 19998 44038 20050 44090
rect 20062 44038 20114 44090
rect 20126 44038 20178 44090
rect 27644 44038 27696 44090
rect 27708 44038 27760 44090
rect 27772 44038 27824 44090
rect 27836 44038 27888 44090
rect 27900 44038 27952 44090
rect 6552 43979 6604 43988
rect 6552 43945 6561 43979
rect 6561 43945 6595 43979
rect 6595 43945 6604 43979
rect 6552 43936 6604 43945
rect 6920 43979 6972 43988
rect 6920 43945 6929 43979
rect 6929 43945 6963 43979
rect 6963 43945 6972 43979
rect 6920 43936 6972 43945
rect 8208 43936 8260 43988
rect 8208 43800 8260 43852
rect 8300 43843 8352 43852
rect 8300 43809 8309 43843
rect 8309 43809 8343 43843
rect 8343 43809 8352 43843
rect 8300 43800 8352 43809
rect 8852 43800 8904 43852
rect 10692 43979 10744 43988
rect 10692 43945 10701 43979
rect 10701 43945 10735 43979
rect 10735 43945 10744 43979
rect 10692 43936 10744 43945
rect 13268 43979 13320 43988
rect 13268 43945 13277 43979
rect 13277 43945 13311 43979
rect 13311 43945 13320 43979
rect 13268 43936 13320 43945
rect 13820 43936 13872 43988
rect 18144 43979 18196 43988
rect 18144 43945 18153 43979
rect 18153 43945 18187 43979
rect 18187 43945 18196 43979
rect 18144 43936 18196 43945
rect 16580 43868 16632 43920
rect 21824 43868 21876 43920
rect 25136 43911 25188 43920
rect 25136 43877 25154 43911
rect 25154 43877 25188 43911
rect 25136 43868 25188 43877
rect 26240 43868 26292 43920
rect 11244 43800 11296 43852
rect 12348 43843 12400 43852
rect 12348 43809 12357 43843
rect 12357 43809 12391 43843
rect 12391 43809 12400 43843
rect 12348 43800 12400 43809
rect 14004 43800 14056 43852
rect 14280 43843 14332 43852
rect 14280 43809 14289 43843
rect 14289 43809 14323 43843
rect 14323 43809 14332 43843
rect 14280 43800 14332 43809
rect 16120 43800 16172 43852
rect 16764 43843 16816 43852
rect 16764 43809 16773 43843
rect 16773 43809 16807 43843
rect 16807 43809 16816 43843
rect 16764 43800 16816 43809
rect 19248 43843 19300 43852
rect 19248 43809 19257 43843
rect 19257 43809 19291 43843
rect 19291 43809 19300 43843
rect 19248 43800 19300 43809
rect 22928 43800 22980 43852
rect 23388 43800 23440 43852
rect 29000 43843 29052 43852
rect 29000 43809 29018 43843
rect 29018 43809 29052 43843
rect 29000 43800 29052 43809
rect 14188 43775 14240 43784
rect 14188 43741 14197 43775
rect 14197 43741 14231 43775
rect 14231 43741 14240 43775
rect 14188 43732 14240 43741
rect 15292 43732 15344 43784
rect 17040 43775 17092 43784
rect 17040 43741 17049 43775
rect 17049 43741 17083 43775
rect 17083 43741 17092 43775
rect 17040 43732 17092 43741
rect 19708 43732 19760 43784
rect 15844 43664 15896 43716
rect 9772 43639 9824 43648
rect 9772 43605 9781 43639
rect 9781 43605 9815 43639
rect 9815 43605 9824 43639
rect 9772 43596 9824 43605
rect 10968 43639 11020 43648
rect 10968 43605 10977 43639
rect 10977 43605 11011 43639
rect 11011 43605 11020 43639
rect 10968 43596 11020 43605
rect 13820 43596 13872 43648
rect 19616 43596 19668 43648
rect 21456 43596 21508 43648
rect 22376 43596 22428 43648
rect 25412 43775 25464 43784
rect 25412 43741 25421 43775
rect 25421 43741 25455 43775
rect 25455 43741 25464 43775
rect 25412 43732 25464 43741
rect 23204 43596 23256 43648
rect 24400 43596 24452 43648
rect 27528 43596 27580 43648
rect 3662 43494 3714 43546
rect 3726 43494 3778 43546
rect 3790 43494 3842 43546
rect 3854 43494 3906 43546
rect 3918 43494 3970 43546
rect 11436 43494 11488 43546
rect 11500 43494 11552 43546
rect 11564 43494 11616 43546
rect 11628 43494 11680 43546
rect 11692 43494 11744 43546
rect 19210 43494 19262 43546
rect 19274 43494 19326 43546
rect 19338 43494 19390 43546
rect 19402 43494 19454 43546
rect 19466 43494 19518 43546
rect 26984 43494 27036 43546
rect 27048 43494 27100 43546
rect 27112 43494 27164 43546
rect 27176 43494 27228 43546
rect 27240 43494 27292 43546
rect 8852 43435 8904 43444
rect 8852 43401 8861 43435
rect 8861 43401 8895 43435
rect 8895 43401 8904 43435
rect 8852 43392 8904 43401
rect 11336 43392 11388 43444
rect 14372 43392 14424 43444
rect 15292 43435 15344 43444
rect 15292 43401 15301 43435
rect 15301 43401 15335 43435
rect 15335 43401 15344 43435
rect 15292 43392 15344 43401
rect 9772 43324 9824 43376
rect 14188 43324 14240 43376
rect 17132 43324 17184 43376
rect 23480 43392 23532 43444
rect 9404 43188 9456 43240
rect 10324 43188 10376 43240
rect 10968 43188 11020 43240
rect 11980 43231 12032 43240
rect 11980 43197 11989 43231
rect 11989 43197 12023 43231
rect 12023 43197 12032 43231
rect 11980 43188 12032 43197
rect 13544 43188 13596 43240
rect 14004 43188 14056 43240
rect 14188 43188 14240 43240
rect 15016 43231 15068 43240
rect 15016 43197 15025 43231
rect 15025 43197 15059 43231
rect 15059 43197 15068 43231
rect 15016 43188 15068 43197
rect 15660 43231 15712 43240
rect 15660 43197 15669 43231
rect 15669 43197 15703 43231
rect 15703 43197 15712 43231
rect 15660 43188 15712 43197
rect 11060 43120 11112 43172
rect 11888 43052 11940 43104
rect 14188 43052 14240 43104
rect 15568 43052 15620 43104
rect 15844 43188 15896 43240
rect 16028 43231 16080 43240
rect 16028 43197 16037 43231
rect 16037 43197 16071 43231
rect 16071 43197 16080 43231
rect 16028 43188 16080 43197
rect 16304 43231 16356 43240
rect 16304 43197 16313 43231
rect 16313 43197 16347 43231
rect 16347 43197 16356 43231
rect 16304 43188 16356 43197
rect 16488 43256 16540 43308
rect 16580 43188 16632 43240
rect 17132 43188 17184 43240
rect 17408 43231 17460 43240
rect 17408 43197 17417 43231
rect 17417 43197 17451 43231
rect 17451 43197 17460 43231
rect 17408 43188 17460 43197
rect 17500 43188 17552 43240
rect 17776 43188 17828 43240
rect 19524 43256 19576 43308
rect 18144 43163 18196 43172
rect 18144 43129 18153 43163
rect 18153 43129 18187 43163
rect 18187 43129 18196 43163
rect 18144 43120 18196 43129
rect 16396 43052 16448 43104
rect 16580 43095 16632 43104
rect 16580 43061 16589 43095
rect 16589 43061 16623 43095
rect 16623 43061 16632 43095
rect 16580 43052 16632 43061
rect 16764 43052 16816 43104
rect 17224 43095 17276 43104
rect 17224 43061 17233 43095
rect 17233 43061 17267 43095
rect 17267 43061 17276 43095
rect 17224 43052 17276 43061
rect 17592 43095 17644 43104
rect 17592 43061 17601 43095
rect 17601 43061 17635 43095
rect 17635 43061 17644 43095
rect 17592 43052 17644 43061
rect 17776 43095 17828 43104
rect 17776 43061 17785 43095
rect 17785 43061 17819 43095
rect 17819 43061 17828 43095
rect 17776 43052 17828 43061
rect 17960 43052 18012 43104
rect 18880 43188 18932 43240
rect 19616 43231 19668 43240
rect 19616 43197 19625 43231
rect 19625 43197 19659 43231
rect 19659 43197 19668 43231
rect 19616 43188 19668 43197
rect 19800 43188 19852 43240
rect 19156 43120 19208 43172
rect 19616 43052 19668 43104
rect 22376 43188 22428 43240
rect 24584 43188 24636 43240
rect 25412 43188 25464 43240
rect 27528 43188 27580 43240
rect 21640 43120 21692 43172
rect 22008 43163 22060 43172
rect 22008 43129 22042 43163
rect 22042 43129 22060 43163
rect 22008 43120 22060 43129
rect 23296 43163 23348 43172
rect 23296 43129 23305 43163
rect 23305 43129 23339 43163
rect 23339 43129 23348 43163
rect 23296 43120 23348 43129
rect 25688 43120 25740 43172
rect 28080 43120 28132 43172
rect 20260 43052 20312 43104
rect 20352 43095 20404 43104
rect 20352 43061 20361 43095
rect 20361 43061 20395 43095
rect 20395 43061 20404 43095
rect 20352 43052 20404 43061
rect 21088 43095 21140 43104
rect 21088 43061 21097 43095
rect 21097 43061 21131 43095
rect 21131 43061 21140 43095
rect 21088 43052 21140 43061
rect 21272 43052 21324 43104
rect 23020 43052 23072 43104
rect 23572 43095 23624 43104
rect 23572 43061 23581 43095
rect 23581 43061 23615 43095
rect 23615 43061 23624 43095
rect 23572 43052 23624 43061
rect 24124 43052 24176 43104
rect 25320 43095 25372 43104
rect 25320 43061 25329 43095
rect 25329 43061 25363 43095
rect 25363 43061 25372 43095
rect 25320 43052 25372 43061
rect 26792 43095 26844 43104
rect 26792 43061 26801 43095
rect 26801 43061 26835 43095
rect 26835 43061 26844 43095
rect 26792 43052 26844 43061
rect 4322 42950 4374 43002
rect 4386 42950 4438 43002
rect 4450 42950 4502 43002
rect 4514 42950 4566 43002
rect 4578 42950 4630 43002
rect 12096 42950 12148 43002
rect 12160 42950 12212 43002
rect 12224 42950 12276 43002
rect 12288 42950 12340 43002
rect 12352 42950 12404 43002
rect 19870 42950 19922 43002
rect 19934 42950 19986 43002
rect 19998 42950 20050 43002
rect 20062 42950 20114 43002
rect 20126 42950 20178 43002
rect 27644 42950 27696 43002
rect 27708 42950 27760 43002
rect 27772 42950 27824 43002
rect 27836 42950 27888 43002
rect 27900 42950 27952 43002
rect 11980 42848 12032 42900
rect 14004 42848 14056 42900
rect 15016 42848 15068 42900
rect 15476 42848 15528 42900
rect 16304 42848 16356 42900
rect 9404 42755 9456 42764
rect 9404 42721 9413 42755
rect 9413 42721 9447 42755
rect 9447 42721 9456 42755
rect 9404 42712 9456 42721
rect 9680 42755 9732 42764
rect 9680 42721 9714 42755
rect 9714 42721 9732 42755
rect 9680 42712 9732 42721
rect 11060 42712 11112 42764
rect 12532 42755 12584 42764
rect 12532 42721 12541 42755
rect 12541 42721 12575 42755
rect 12575 42721 12584 42755
rect 12532 42712 12584 42721
rect 13544 42712 13596 42764
rect 14648 42712 14700 42764
rect 16212 42712 16264 42764
rect 16672 42848 16724 42900
rect 19708 42891 19760 42900
rect 19708 42857 19717 42891
rect 19717 42857 19751 42891
rect 19751 42857 19760 42891
rect 19708 42848 19760 42857
rect 23296 42848 23348 42900
rect 17132 42780 17184 42832
rect 11336 42644 11388 42696
rect 14280 42687 14332 42696
rect 14280 42653 14289 42687
rect 14289 42653 14323 42687
rect 14323 42653 14332 42687
rect 14280 42644 14332 42653
rect 15016 42644 15068 42696
rect 16304 42644 16356 42696
rect 16948 42712 17000 42764
rect 18144 42780 18196 42832
rect 20536 42780 20588 42832
rect 17408 42755 17460 42764
rect 17408 42721 17417 42755
rect 17417 42721 17451 42755
rect 17451 42721 17460 42755
rect 17408 42712 17460 42721
rect 17960 42755 18012 42764
rect 17960 42721 17969 42755
rect 17969 42721 18003 42755
rect 18003 42721 18012 42755
rect 17960 42712 18012 42721
rect 19524 42712 19576 42764
rect 16028 42576 16080 42628
rect 19616 42576 19668 42628
rect 10968 42551 11020 42560
rect 10968 42517 10977 42551
rect 10977 42517 11011 42551
rect 11011 42517 11020 42551
rect 10968 42508 11020 42517
rect 17500 42508 17552 42560
rect 18972 42508 19024 42560
rect 19156 42508 19208 42560
rect 20076 42755 20128 42764
rect 20076 42721 20085 42755
rect 20085 42721 20119 42755
rect 20119 42721 20128 42755
rect 20076 42712 20128 42721
rect 20260 42712 20312 42764
rect 20352 42755 20404 42764
rect 20352 42721 20361 42755
rect 20361 42721 20395 42755
rect 20395 42721 20404 42755
rect 20352 42712 20404 42721
rect 21272 42755 21324 42764
rect 21272 42721 21281 42755
rect 21281 42721 21315 42755
rect 21315 42721 21324 42755
rect 21272 42712 21324 42721
rect 21364 42712 21416 42764
rect 22928 42755 22980 42764
rect 22928 42721 22937 42755
rect 22937 42721 22971 42755
rect 22971 42721 22980 42755
rect 22928 42712 22980 42721
rect 23020 42755 23072 42764
rect 23020 42721 23029 42755
rect 23029 42721 23063 42755
rect 23063 42721 23072 42755
rect 23020 42712 23072 42721
rect 23296 42755 23348 42764
rect 23296 42721 23305 42755
rect 23305 42721 23339 42755
rect 23339 42721 23348 42755
rect 23296 42712 23348 42721
rect 23480 42712 23532 42764
rect 23756 42712 23808 42764
rect 24492 42848 24544 42900
rect 23940 42755 23992 42764
rect 23940 42721 23949 42755
rect 23949 42721 23983 42755
rect 23983 42721 23992 42755
rect 23940 42712 23992 42721
rect 24032 42712 24084 42764
rect 25228 42780 25280 42832
rect 24492 42755 24544 42764
rect 24492 42721 24501 42755
rect 24501 42721 24535 42755
rect 24535 42721 24544 42755
rect 24492 42712 24544 42721
rect 24584 42755 24636 42764
rect 24584 42721 24593 42755
rect 24593 42721 24627 42755
rect 24627 42721 24636 42755
rect 24584 42712 24636 42721
rect 27528 42712 27580 42764
rect 25320 42644 25372 42696
rect 22652 42576 22704 42628
rect 23940 42576 23992 42628
rect 24216 42576 24268 42628
rect 29276 42576 29328 42628
rect 22284 42508 22336 42560
rect 23388 42508 23440 42560
rect 29368 42508 29420 42560
rect 3662 42406 3714 42458
rect 3726 42406 3778 42458
rect 3790 42406 3842 42458
rect 3854 42406 3906 42458
rect 3918 42406 3970 42458
rect 11436 42406 11488 42458
rect 11500 42406 11552 42458
rect 11564 42406 11616 42458
rect 11628 42406 11680 42458
rect 11692 42406 11744 42458
rect 19210 42406 19262 42458
rect 19274 42406 19326 42458
rect 19338 42406 19390 42458
rect 19402 42406 19454 42458
rect 19466 42406 19518 42458
rect 26984 42406 27036 42458
rect 27048 42406 27100 42458
rect 27112 42406 27164 42458
rect 27176 42406 27228 42458
rect 27240 42406 27292 42458
rect 13544 42347 13596 42356
rect 13544 42313 13553 42347
rect 13553 42313 13587 42347
rect 13587 42313 13596 42347
rect 13544 42304 13596 42313
rect 14280 42304 14332 42356
rect 15016 42347 15068 42356
rect 15016 42313 15025 42347
rect 15025 42313 15059 42347
rect 15059 42313 15068 42347
rect 15016 42304 15068 42313
rect 17040 42304 17092 42356
rect 17316 42347 17368 42356
rect 17316 42313 17325 42347
rect 17325 42313 17359 42347
rect 17359 42313 17368 42347
rect 17316 42304 17368 42313
rect 13728 42143 13780 42152
rect 13728 42109 13737 42143
rect 13737 42109 13771 42143
rect 13771 42109 13780 42143
rect 13728 42100 13780 42109
rect 14004 42143 14056 42152
rect 14004 42109 14013 42143
rect 14013 42109 14047 42143
rect 14047 42109 14056 42143
rect 14004 42100 14056 42109
rect 14188 42143 14240 42152
rect 14188 42109 14197 42143
rect 14197 42109 14231 42143
rect 14231 42109 14240 42143
rect 14188 42100 14240 42109
rect 14648 42143 14700 42152
rect 14648 42109 14657 42143
rect 14657 42109 14691 42143
rect 14691 42109 14700 42143
rect 14648 42100 14700 42109
rect 15476 42236 15528 42288
rect 16396 42236 16448 42288
rect 15660 42168 15712 42220
rect 15476 42143 15528 42152
rect 15476 42109 15485 42143
rect 15485 42109 15519 42143
rect 15519 42109 15528 42143
rect 15476 42100 15528 42109
rect 15752 42143 15804 42152
rect 15752 42109 15761 42143
rect 15761 42109 15795 42143
rect 15795 42109 15804 42143
rect 15752 42100 15804 42109
rect 16856 42168 16908 42220
rect 15200 41964 15252 42016
rect 15752 41964 15804 42016
rect 16764 42143 16816 42152
rect 16764 42109 16773 42143
rect 16773 42109 16807 42143
rect 16807 42109 16816 42143
rect 16764 42100 16816 42109
rect 16948 42143 17000 42152
rect 16948 42109 16957 42143
rect 16957 42109 16991 42143
rect 16991 42109 17000 42143
rect 16948 42100 17000 42109
rect 17224 42032 17276 42084
rect 18696 42304 18748 42356
rect 19432 42304 19484 42356
rect 19616 42304 19668 42356
rect 21364 42304 21416 42356
rect 23296 42304 23348 42356
rect 18972 42236 19024 42288
rect 20076 42236 20128 42288
rect 18512 42143 18564 42152
rect 18512 42109 18530 42143
rect 18530 42109 18564 42143
rect 18512 42100 18564 42109
rect 18696 42143 18748 42152
rect 18696 42109 18705 42143
rect 18705 42109 18739 42143
rect 18739 42109 18748 42143
rect 18696 42100 18748 42109
rect 18144 41964 18196 42016
rect 18328 41964 18380 42016
rect 19064 42143 19116 42152
rect 19064 42109 19073 42143
rect 19073 42109 19107 42143
rect 19107 42109 19116 42143
rect 19064 42100 19116 42109
rect 19156 42100 19208 42152
rect 19340 42075 19392 42084
rect 19340 42041 19349 42075
rect 19349 42041 19383 42075
rect 19383 42041 19392 42075
rect 19340 42032 19392 42041
rect 19524 42100 19576 42152
rect 19708 42100 19760 42152
rect 20260 42143 20312 42152
rect 20260 42109 20269 42143
rect 20269 42109 20303 42143
rect 20303 42109 20312 42143
rect 20260 42100 20312 42109
rect 21088 42168 21140 42220
rect 23664 42236 23716 42288
rect 24216 42236 24268 42288
rect 19800 42032 19852 42084
rect 20352 41964 20404 42016
rect 20444 41964 20496 42016
rect 20812 42100 20864 42152
rect 20996 42100 21048 42152
rect 21640 42100 21692 42152
rect 22008 42100 22060 42152
rect 22376 42143 22428 42152
rect 22376 42109 22385 42143
rect 22385 42109 22419 42143
rect 22419 42109 22428 42143
rect 22376 42100 22428 42109
rect 22928 42100 22980 42152
rect 26792 42168 26844 42220
rect 23204 42100 23256 42152
rect 23388 42143 23440 42152
rect 23388 42109 23397 42143
rect 23397 42109 23431 42143
rect 23431 42109 23440 42143
rect 23388 42100 23440 42109
rect 24032 42143 24084 42152
rect 24032 42109 24041 42143
rect 24041 42109 24075 42143
rect 24075 42109 24084 42143
rect 24032 42100 24084 42109
rect 24124 42143 24176 42152
rect 24124 42109 24133 42143
rect 24133 42109 24167 42143
rect 24167 42109 24176 42143
rect 24124 42100 24176 42109
rect 24400 42143 24452 42152
rect 24400 42109 24409 42143
rect 24409 42109 24443 42143
rect 24443 42109 24452 42143
rect 24400 42100 24452 42109
rect 26240 42100 26292 42152
rect 27528 42100 27580 42152
rect 29552 42143 29604 42152
rect 29552 42109 29561 42143
rect 29561 42109 29595 42143
rect 29595 42109 29604 42143
rect 29552 42100 29604 42109
rect 23572 42032 23624 42084
rect 20996 41964 21048 42016
rect 21272 41964 21324 42016
rect 22836 42007 22888 42016
rect 22836 41973 22845 42007
rect 22845 41973 22879 42007
rect 22879 41973 22888 42007
rect 22836 41964 22888 41973
rect 22928 41964 22980 42016
rect 28724 42032 28776 42084
rect 30748 42100 30800 42152
rect 26424 41964 26476 42016
rect 27988 41964 28040 42016
rect 29000 42007 29052 42016
rect 29000 41973 29009 42007
rect 29009 41973 29043 42007
rect 29043 41973 29052 42007
rect 29000 41964 29052 41973
rect 29276 41964 29328 42016
rect 4322 41862 4374 41914
rect 4386 41862 4438 41914
rect 4450 41862 4502 41914
rect 4514 41862 4566 41914
rect 4578 41862 4630 41914
rect 12096 41862 12148 41914
rect 12160 41862 12212 41914
rect 12224 41862 12276 41914
rect 12288 41862 12340 41914
rect 12352 41862 12404 41914
rect 19870 41862 19922 41914
rect 19934 41862 19986 41914
rect 19998 41862 20050 41914
rect 20062 41862 20114 41914
rect 20126 41862 20178 41914
rect 27644 41862 27696 41914
rect 27708 41862 27760 41914
rect 27772 41862 27824 41914
rect 27836 41862 27888 41914
rect 27900 41862 27952 41914
rect 9680 41803 9732 41812
rect 9680 41769 9689 41803
rect 9689 41769 9723 41803
rect 9723 41769 9732 41803
rect 9680 41760 9732 41769
rect 13820 41803 13872 41812
rect 13820 41769 13829 41803
rect 13829 41769 13863 41803
rect 13863 41769 13872 41803
rect 13820 41760 13872 41769
rect 14280 41760 14332 41812
rect 16764 41760 16816 41812
rect 17132 41760 17184 41812
rect 18512 41760 18564 41812
rect 20076 41760 20128 41812
rect 24032 41760 24084 41812
rect 28816 41760 28868 41812
rect 29552 41760 29604 41812
rect 30748 41803 30800 41812
rect 30748 41769 30757 41803
rect 30757 41769 30791 41803
rect 30791 41769 30800 41803
rect 30748 41760 30800 41769
rect 10968 41692 11020 41744
rect 16212 41692 16264 41744
rect 20260 41692 20312 41744
rect 22652 41692 22704 41744
rect 10140 41667 10192 41676
rect 10140 41633 10149 41667
rect 10149 41633 10183 41667
rect 10183 41633 10192 41667
rect 10140 41624 10192 41633
rect 10324 41667 10376 41676
rect 10324 41633 10333 41667
rect 10333 41633 10367 41667
rect 10367 41633 10376 41667
rect 10324 41624 10376 41633
rect 10784 41624 10836 41676
rect 10416 41556 10468 41608
rect 12716 41556 12768 41608
rect 14004 41624 14056 41676
rect 14832 41624 14884 41676
rect 17868 41667 17920 41676
rect 17868 41633 17877 41667
rect 17877 41633 17911 41667
rect 17911 41633 17920 41667
rect 17868 41624 17920 41633
rect 21272 41667 21324 41676
rect 21272 41633 21281 41667
rect 21281 41633 21315 41667
rect 21315 41633 21324 41667
rect 21272 41624 21324 41633
rect 21364 41624 21416 41676
rect 19616 41556 19668 41608
rect 20444 41556 20496 41608
rect 15016 41488 15068 41540
rect 15844 41488 15896 41540
rect 16120 41488 16172 41540
rect 20996 41488 21048 41540
rect 23204 41667 23256 41676
rect 23204 41633 23213 41667
rect 23213 41633 23247 41667
rect 23247 41633 23256 41667
rect 23204 41624 23256 41633
rect 23940 41667 23992 41676
rect 23940 41633 23949 41667
rect 23949 41633 23983 41667
rect 23983 41633 23992 41667
rect 23940 41624 23992 41633
rect 26424 41667 26476 41676
rect 26424 41633 26433 41667
rect 26433 41633 26467 41667
rect 26467 41633 26476 41667
rect 26424 41624 26476 41633
rect 26700 41667 26752 41676
rect 26700 41633 26734 41667
rect 26734 41633 26752 41667
rect 26700 41624 26752 41633
rect 27988 41624 28040 41676
rect 28172 41667 28224 41676
rect 28172 41633 28206 41667
rect 28206 41633 28224 41667
rect 28172 41624 28224 41633
rect 29368 41667 29420 41676
rect 29368 41633 29377 41667
rect 29377 41633 29411 41667
rect 29411 41633 29420 41667
rect 29368 41624 29420 41633
rect 29460 41624 29512 41676
rect 23940 41488 23992 41540
rect 12440 41463 12492 41472
rect 12440 41429 12449 41463
rect 12449 41429 12483 41463
rect 12483 41429 12492 41463
rect 12440 41420 12492 41429
rect 15384 41420 15436 41472
rect 15660 41420 15712 41472
rect 17592 41420 17644 41472
rect 20536 41420 20588 41472
rect 23480 41463 23532 41472
rect 23480 41429 23489 41463
rect 23489 41429 23523 41463
rect 23523 41429 23532 41463
rect 23480 41420 23532 41429
rect 23756 41463 23808 41472
rect 23756 41429 23765 41463
rect 23765 41429 23799 41463
rect 23799 41429 23808 41463
rect 23756 41420 23808 41429
rect 24584 41420 24636 41472
rect 27804 41463 27856 41472
rect 27804 41429 27813 41463
rect 27813 41429 27847 41463
rect 27847 41429 27856 41463
rect 27804 41420 27856 41429
rect 3662 41318 3714 41370
rect 3726 41318 3778 41370
rect 3790 41318 3842 41370
rect 3854 41318 3906 41370
rect 3918 41318 3970 41370
rect 11436 41318 11488 41370
rect 11500 41318 11552 41370
rect 11564 41318 11616 41370
rect 11628 41318 11680 41370
rect 11692 41318 11744 41370
rect 19210 41318 19262 41370
rect 19274 41318 19326 41370
rect 19338 41318 19390 41370
rect 19402 41318 19454 41370
rect 19466 41318 19518 41370
rect 26984 41318 27036 41370
rect 27048 41318 27100 41370
rect 27112 41318 27164 41370
rect 27176 41318 27228 41370
rect 27240 41318 27292 41370
rect 8300 41012 8352 41064
rect 9680 41216 9732 41268
rect 10140 41216 10192 41268
rect 9220 41148 9272 41200
rect 12624 41216 12676 41268
rect 8944 41055 8996 41064
rect 8944 41021 8953 41055
rect 8953 41021 8987 41055
rect 8987 41021 8996 41055
rect 8944 41012 8996 41021
rect 9220 41055 9272 41064
rect 9220 41021 9229 41055
rect 9229 41021 9263 41055
rect 9263 41021 9272 41055
rect 9220 41012 9272 41021
rect 9496 41080 9548 41132
rect 9772 41012 9824 41064
rect 10600 41080 10652 41132
rect 10784 41080 10836 41132
rect 10140 41055 10192 41064
rect 10140 41021 10149 41055
rect 10149 41021 10183 41055
rect 10183 41021 10192 41055
rect 10140 41012 10192 41021
rect 10324 41055 10376 41064
rect 10324 41021 10333 41055
rect 10333 41021 10367 41055
rect 10367 41021 10376 41055
rect 10324 41012 10376 41021
rect 10968 41012 11020 41064
rect 11060 41055 11112 41064
rect 11060 41021 11069 41055
rect 11069 41021 11103 41055
rect 11103 41021 11112 41055
rect 11060 41012 11112 41021
rect 11796 40944 11848 40996
rect 8116 40876 8168 40928
rect 8668 40919 8720 40928
rect 8668 40885 8677 40919
rect 8677 40885 8711 40919
rect 8711 40885 8720 40919
rect 8668 40876 8720 40885
rect 9128 40876 9180 40928
rect 12808 40987 12860 40996
rect 12808 40953 12817 40987
rect 12817 40953 12851 40987
rect 12851 40953 12860 40987
rect 12808 40944 12860 40953
rect 12532 40876 12584 40928
rect 12716 40919 12768 40928
rect 12716 40885 12725 40919
rect 12725 40885 12759 40919
rect 12759 40885 12768 40919
rect 13084 40944 13136 40996
rect 15200 41148 15252 41200
rect 15568 41259 15620 41268
rect 15568 41225 15577 41259
rect 15577 41225 15611 41259
rect 15611 41225 15620 41259
rect 15568 41216 15620 41225
rect 16488 41216 16540 41268
rect 17316 41216 17368 41268
rect 18144 41259 18196 41268
rect 18144 41225 18153 41259
rect 18153 41225 18187 41259
rect 18187 41225 18196 41259
rect 18144 41216 18196 41225
rect 19064 41216 19116 41268
rect 20352 41216 20404 41268
rect 21364 41216 21416 41268
rect 22652 41216 22704 41268
rect 26608 41216 26660 41268
rect 28172 41259 28224 41268
rect 28172 41225 28181 41259
rect 28181 41225 28215 41259
rect 28215 41225 28224 41259
rect 28172 41216 28224 41225
rect 29460 41216 29512 41268
rect 15108 41055 15160 41064
rect 15108 41021 15117 41055
rect 15117 41021 15151 41055
rect 15151 41021 15160 41055
rect 15108 41012 15160 41021
rect 15200 41055 15252 41064
rect 15200 41021 15209 41055
rect 15209 41021 15243 41055
rect 15243 41021 15252 41055
rect 15200 41012 15252 41021
rect 15384 41012 15436 41064
rect 15568 41012 15620 41064
rect 15936 41012 15988 41064
rect 16120 41055 16172 41064
rect 16120 41021 16129 41055
rect 16129 41021 16163 41055
rect 16163 41021 16172 41055
rect 16120 41012 16172 41021
rect 16304 41012 16356 41064
rect 17132 41080 17184 41132
rect 17592 41080 17644 41132
rect 17040 41012 17092 41064
rect 12716 40876 12768 40885
rect 13268 40876 13320 40928
rect 14096 40876 14148 40928
rect 14372 40876 14424 40928
rect 15200 40876 15252 40928
rect 15292 40876 15344 40928
rect 17408 40944 17460 40996
rect 17592 40987 17644 40996
rect 17592 40953 17601 40987
rect 17601 40953 17635 40987
rect 17635 40953 17644 40987
rect 17592 40944 17644 40953
rect 16672 40919 16724 40928
rect 16672 40885 16681 40919
rect 16681 40885 16715 40919
rect 16715 40885 16724 40919
rect 16672 40876 16724 40885
rect 17316 40876 17368 40928
rect 17868 41012 17920 41064
rect 17960 41012 18012 41064
rect 19340 41012 19392 41064
rect 19524 41012 19576 41064
rect 19708 41012 19760 41064
rect 23480 41080 23532 41132
rect 26332 41148 26384 41200
rect 19248 40944 19300 40996
rect 20260 41012 20312 41064
rect 20352 41055 20404 41064
rect 20352 41021 20361 41055
rect 20361 41021 20395 41055
rect 20395 41021 20404 41055
rect 20352 41012 20404 41021
rect 20444 41055 20496 41064
rect 20444 41021 20453 41055
rect 20453 41021 20487 41055
rect 20487 41021 20496 41055
rect 20444 41012 20496 41021
rect 20076 40944 20128 40996
rect 22100 41012 22152 41064
rect 22376 41012 22428 41064
rect 23756 41012 23808 41064
rect 23940 41055 23992 41064
rect 23940 41021 23949 41055
rect 23949 41021 23983 41055
rect 23983 41021 23992 41055
rect 23940 41012 23992 41021
rect 25320 41012 25372 41064
rect 26148 41012 26200 41064
rect 18052 40876 18104 40928
rect 23480 40944 23532 40996
rect 24676 40944 24728 40996
rect 24860 40944 24912 40996
rect 26792 41080 26844 41132
rect 27804 41080 27856 41132
rect 28908 41080 28960 41132
rect 29552 41080 29604 41132
rect 27436 40944 27488 40996
rect 20352 40876 20404 40928
rect 21916 40876 21968 40928
rect 23296 40919 23348 40928
rect 23296 40885 23305 40919
rect 23305 40885 23339 40919
rect 23339 40885 23348 40919
rect 23296 40876 23348 40885
rect 25228 40876 25280 40928
rect 25504 40919 25556 40928
rect 25504 40885 25513 40919
rect 25513 40885 25547 40919
rect 25547 40885 25556 40919
rect 25504 40876 25556 40885
rect 26516 40876 26568 40928
rect 28632 41055 28684 41064
rect 28632 41021 28641 41055
rect 28641 41021 28675 41055
rect 28675 41021 28684 41055
rect 28632 41012 28684 41021
rect 29276 41055 29328 41064
rect 29276 41021 29285 41055
rect 29285 41021 29319 41055
rect 29319 41021 29328 41055
rect 29276 41012 29328 41021
rect 31116 41012 31168 41064
rect 28540 40876 28592 40928
rect 29460 40919 29512 40928
rect 29460 40885 29469 40919
rect 29469 40885 29503 40919
rect 29503 40885 29512 40919
rect 29460 40876 29512 40885
rect 30748 40944 30800 40996
rect 30932 40876 30984 40928
rect 4322 40774 4374 40826
rect 4386 40774 4438 40826
rect 4450 40774 4502 40826
rect 4514 40774 4566 40826
rect 4578 40774 4630 40826
rect 12096 40774 12148 40826
rect 12160 40774 12212 40826
rect 12224 40774 12276 40826
rect 12288 40774 12340 40826
rect 12352 40774 12404 40826
rect 19870 40774 19922 40826
rect 19934 40774 19986 40826
rect 19998 40774 20050 40826
rect 20062 40774 20114 40826
rect 20126 40774 20178 40826
rect 27644 40774 27696 40826
rect 27708 40774 27760 40826
rect 27772 40774 27824 40826
rect 27836 40774 27888 40826
rect 27900 40774 27952 40826
rect 10140 40672 10192 40724
rect 10968 40715 11020 40724
rect 10968 40681 10977 40715
rect 10977 40681 11011 40715
rect 11011 40681 11020 40715
rect 10968 40672 11020 40681
rect 11796 40715 11848 40724
rect 11796 40681 11805 40715
rect 11805 40681 11839 40715
rect 11839 40681 11848 40715
rect 11796 40672 11848 40681
rect 8944 40604 8996 40656
rect 10232 40604 10284 40656
rect 8116 40579 8168 40588
rect 8116 40545 8125 40579
rect 8125 40545 8159 40579
rect 8159 40545 8168 40579
rect 8116 40536 8168 40545
rect 8852 40536 8904 40588
rect 9588 40536 9640 40588
rect 11980 40604 12032 40656
rect 12440 40672 12492 40724
rect 15108 40672 15160 40724
rect 9864 40400 9916 40452
rect 10692 40468 10744 40520
rect 12164 40579 12216 40588
rect 12164 40545 12173 40579
rect 12173 40545 12207 40579
rect 12207 40545 12216 40579
rect 12164 40536 12216 40545
rect 12256 40579 12308 40588
rect 12256 40545 12265 40579
rect 12265 40545 12299 40579
rect 12299 40545 12308 40579
rect 12256 40536 12308 40545
rect 12716 40604 12768 40656
rect 16764 40672 16816 40724
rect 17224 40672 17276 40724
rect 17408 40672 17460 40724
rect 19248 40672 19300 40724
rect 20352 40672 20404 40724
rect 23204 40672 23256 40724
rect 23940 40672 23992 40724
rect 24860 40715 24912 40724
rect 24860 40681 24869 40715
rect 24869 40681 24903 40715
rect 24903 40681 24912 40715
rect 24860 40672 24912 40681
rect 26700 40672 26752 40724
rect 30748 40672 30800 40724
rect 31116 40715 31168 40724
rect 31116 40681 31125 40715
rect 31125 40681 31159 40715
rect 31159 40681 31168 40715
rect 31116 40672 31168 40681
rect 12532 40536 12584 40588
rect 12900 40579 12952 40588
rect 12900 40545 12909 40579
rect 12909 40545 12943 40579
rect 12943 40545 12952 40579
rect 12900 40536 12952 40545
rect 12992 40579 13044 40588
rect 12992 40545 13001 40579
rect 13001 40545 13035 40579
rect 13035 40545 13044 40579
rect 12992 40536 13044 40545
rect 10968 40400 11020 40452
rect 11796 40400 11848 40452
rect 13268 40579 13320 40588
rect 13268 40545 13277 40579
rect 13277 40545 13311 40579
rect 13311 40545 13320 40579
rect 13268 40536 13320 40545
rect 14096 40579 14148 40588
rect 14096 40545 14105 40579
rect 14105 40545 14139 40579
rect 14139 40545 14148 40579
rect 14096 40536 14148 40545
rect 14372 40579 14424 40588
rect 14372 40545 14381 40579
rect 14381 40545 14415 40579
rect 14415 40545 14424 40579
rect 14372 40536 14424 40545
rect 16212 40536 16264 40588
rect 16764 40579 16816 40588
rect 16764 40545 16773 40579
rect 16773 40545 16807 40579
rect 16807 40545 16816 40579
rect 16764 40536 16816 40545
rect 16856 40468 16908 40520
rect 17132 40536 17184 40588
rect 17592 40604 17644 40656
rect 17776 40604 17828 40656
rect 18420 40604 18472 40656
rect 18604 40604 18656 40656
rect 21456 40647 21508 40656
rect 21456 40613 21465 40647
rect 21465 40613 21499 40647
rect 21499 40613 21508 40647
rect 21456 40604 21508 40613
rect 26240 40604 26292 40656
rect 27344 40604 27396 40656
rect 14096 40400 14148 40452
rect 16764 40400 16816 40452
rect 17316 40511 17368 40520
rect 17316 40477 17325 40511
rect 17325 40477 17359 40511
rect 17359 40477 17368 40511
rect 17316 40468 17368 40477
rect 17960 40536 18012 40588
rect 18880 40579 18932 40588
rect 18880 40545 18889 40579
rect 18889 40545 18923 40579
rect 18923 40545 18932 40579
rect 18880 40536 18932 40545
rect 19340 40536 19392 40588
rect 19616 40536 19668 40588
rect 19800 40536 19852 40588
rect 20720 40536 20772 40588
rect 21916 40579 21968 40588
rect 21916 40545 21925 40579
rect 21925 40545 21959 40579
rect 21959 40545 21968 40579
rect 21916 40536 21968 40545
rect 22192 40579 22244 40588
rect 22192 40545 22226 40579
rect 22226 40545 22244 40579
rect 22192 40536 22244 40545
rect 23572 40536 23624 40588
rect 24952 40536 25004 40588
rect 25504 40536 25556 40588
rect 17684 40400 17736 40452
rect 19064 40400 19116 40452
rect 25044 40511 25096 40520
rect 25044 40477 25053 40511
rect 25053 40477 25087 40511
rect 25087 40477 25096 40511
rect 26516 40536 26568 40588
rect 26608 40579 26660 40588
rect 26608 40545 26617 40579
rect 26617 40545 26651 40579
rect 26651 40545 26660 40579
rect 26608 40536 26660 40545
rect 28356 40579 28408 40588
rect 28356 40545 28365 40579
rect 28365 40545 28399 40579
rect 28399 40545 28408 40579
rect 28356 40536 28408 40545
rect 28540 40536 28592 40588
rect 29460 40536 29512 40588
rect 30932 40579 30984 40588
rect 30932 40545 30941 40579
rect 30941 40545 30975 40579
rect 30975 40545 30984 40579
rect 30932 40536 30984 40545
rect 31024 40579 31076 40588
rect 31024 40545 31033 40579
rect 31033 40545 31067 40579
rect 31067 40545 31076 40579
rect 31024 40536 31076 40545
rect 25044 40468 25096 40477
rect 26148 40468 26200 40520
rect 26792 40511 26844 40520
rect 26792 40477 26801 40511
rect 26801 40477 26835 40511
rect 26835 40477 26844 40511
rect 26792 40468 26844 40477
rect 27436 40468 27488 40520
rect 29552 40468 29604 40520
rect 25136 40400 25188 40452
rect 9496 40375 9548 40384
rect 9496 40341 9505 40375
rect 9505 40341 9539 40375
rect 9539 40341 9548 40375
rect 9496 40332 9548 40341
rect 10692 40332 10744 40384
rect 12624 40375 12676 40384
rect 12624 40341 12633 40375
rect 12633 40341 12667 40375
rect 12667 40341 12676 40375
rect 12624 40332 12676 40341
rect 15844 40332 15896 40384
rect 17408 40332 17460 40384
rect 17500 40332 17552 40384
rect 18696 40375 18748 40384
rect 18696 40341 18705 40375
rect 18705 40341 18739 40375
rect 18739 40341 18748 40375
rect 18696 40332 18748 40341
rect 21456 40332 21508 40384
rect 23480 40332 23532 40384
rect 28632 40375 28684 40384
rect 28632 40341 28641 40375
rect 28641 40341 28675 40375
rect 28675 40341 28684 40375
rect 28632 40332 28684 40341
rect 30380 40332 30432 40384
rect 3662 40230 3714 40282
rect 3726 40230 3778 40282
rect 3790 40230 3842 40282
rect 3854 40230 3906 40282
rect 3918 40230 3970 40282
rect 11436 40230 11488 40282
rect 11500 40230 11552 40282
rect 11564 40230 11616 40282
rect 11628 40230 11680 40282
rect 11692 40230 11744 40282
rect 19210 40230 19262 40282
rect 19274 40230 19326 40282
rect 19338 40230 19390 40282
rect 19402 40230 19454 40282
rect 19466 40230 19518 40282
rect 26984 40230 27036 40282
rect 27048 40230 27100 40282
rect 27112 40230 27164 40282
rect 27176 40230 27228 40282
rect 27240 40230 27292 40282
rect 8852 40171 8904 40180
rect 8852 40137 8861 40171
rect 8861 40137 8895 40171
rect 8895 40137 8904 40171
rect 8852 40128 8904 40137
rect 9680 40171 9732 40180
rect 9680 40137 9689 40171
rect 9689 40137 9723 40171
rect 9723 40137 9732 40171
rect 9680 40128 9732 40137
rect 12256 40128 12308 40180
rect 15384 40171 15436 40180
rect 15384 40137 15393 40171
rect 15393 40137 15427 40171
rect 15427 40137 15436 40171
rect 15384 40128 15436 40137
rect 16120 40171 16172 40180
rect 16120 40137 16129 40171
rect 16129 40137 16163 40171
rect 16163 40137 16172 40171
rect 16120 40128 16172 40137
rect 16856 40128 16908 40180
rect 17868 40128 17920 40180
rect 10140 40060 10192 40112
rect 8668 39992 8720 40044
rect 9128 39967 9180 39976
rect 9128 39933 9137 39967
rect 9137 39933 9171 39967
rect 9171 39933 9180 39967
rect 9128 39924 9180 39933
rect 9220 39967 9272 39976
rect 9220 39933 9229 39967
rect 9229 39933 9263 39967
rect 9263 39933 9272 39967
rect 9220 39924 9272 39933
rect 9588 39992 9640 40044
rect 10968 40060 11020 40112
rect 9956 39924 10008 39976
rect 11336 39992 11388 40044
rect 10600 39967 10652 39976
rect 10600 39933 10609 39967
rect 10609 39933 10643 39967
rect 10643 39933 10652 39967
rect 10600 39924 10652 39933
rect 10692 39967 10744 39976
rect 10692 39933 10701 39967
rect 10701 39933 10735 39967
rect 10735 39933 10744 39967
rect 10692 39924 10744 39933
rect 10876 39967 10928 39976
rect 10876 39933 10885 39967
rect 10885 39933 10919 39967
rect 10919 39933 10928 39967
rect 10876 39924 10928 39933
rect 13084 40035 13136 40044
rect 13084 40001 13093 40035
rect 13093 40001 13127 40035
rect 13127 40001 13136 40035
rect 13084 39992 13136 40001
rect 13268 40060 13320 40112
rect 15016 39992 15068 40044
rect 15384 39992 15436 40044
rect 8392 39831 8444 39840
rect 8392 39797 8401 39831
rect 8401 39797 8435 39831
rect 8435 39797 8444 39831
rect 8392 39788 8444 39797
rect 10232 39856 10284 39908
rect 10324 39856 10376 39908
rect 9588 39788 9640 39840
rect 13544 39967 13596 39976
rect 13544 39933 13553 39967
rect 13553 39933 13587 39967
rect 13587 39933 13596 39967
rect 13544 39924 13596 39933
rect 14096 39924 14148 39976
rect 15568 39967 15620 39976
rect 15568 39933 15577 39967
rect 15577 39933 15611 39967
rect 15611 39933 15620 39967
rect 15568 39924 15620 39933
rect 11336 39856 11388 39908
rect 12164 39856 12216 39908
rect 12716 39856 12768 39908
rect 13452 39856 13504 39908
rect 11612 39831 11664 39840
rect 11612 39797 11621 39831
rect 11621 39797 11655 39831
rect 11655 39797 11664 39831
rect 11612 39788 11664 39797
rect 11888 39788 11940 39840
rect 12532 39788 12584 39840
rect 12900 39788 12952 39840
rect 13636 39788 13688 39840
rect 14924 39831 14976 39840
rect 14924 39797 14933 39831
rect 14933 39797 14967 39831
rect 14967 39797 14976 39831
rect 14924 39788 14976 39797
rect 15844 39967 15896 39976
rect 15844 39933 15853 39967
rect 15853 39933 15887 39967
rect 15887 39933 15896 39967
rect 15844 39924 15896 39933
rect 15936 39967 15988 39976
rect 15936 39933 15945 39967
rect 15945 39933 15979 39967
rect 15979 39933 15988 39967
rect 15936 39924 15988 39933
rect 16764 40060 16816 40112
rect 17776 40060 17828 40112
rect 18144 40060 18196 40112
rect 16672 39992 16724 40044
rect 18880 39992 18932 40044
rect 16580 39967 16632 39976
rect 16580 39933 16589 39967
rect 16589 39933 16623 39967
rect 16623 39933 16632 39967
rect 16580 39924 16632 39933
rect 16948 39924 17000 39976
rect 17132 39967 17184 39976
rect 17132 39933 17141 39967
rect 17141 39933 17175 39967
rect 17175 39933 17184 39967
rect 17132 39924 17184 39933
rect 17408 39924 17460 39976
rect 18972 39967 19024 39976
rect 18972 39933 18981 39967
rect 18981 39933 19015 39967
rect 19015 39933 19024 39967
rect 18972 39924 19024 39933
rect 19800 39924 19852 39976
rect 20352 39856 20404 39908
rect 21088 39924 21140 39976
rect 21456 39967 21508 39976
rect 21456 39933 21465 39967
rect 21465 39933 21499 39967
rect 21499 39933 21508 39967
rect 21456 39924 21508 39933
rect 22192 40060 22244 40112
rect 26884 40128 26936 40180
rect 27436 40171 27488 40180
rect 27436 40137 27445 40171
rect 27445 40137 27479 40171
rect 27479 40137 27488 40171
rect 27436 40128 27488 40137
rect 28540 40128 28592 40180
rect 23020 40060 23072 40112
rect 23388 40060 23440 40112
rect 26056 40060 26108 40112
rect 28448 40060 28500 40112
rect 28908 40060 28960 40112
rect 22376 39967 22428 39976
rect 16396 39788 16448 39840
rect 16488 39788 16540 39840
rect 16672 39788 16724 39840
rect 17316 39788 17368 39840
rect 20536 39831 20588 39840
rect 20536 39797 20545 39831
rect 20545 39797 20579 39831
rect 20579 39797 20588 39831
rect 20536 39788 20588 39797
rect 20628 39788 20680 39840
rect 22376 39933 22385 39967
rect 22385 39933 22419 39967
rect 22419 39933 22428 39967
rect 22376 39924 22428 39933
rect 23204 39924 23256 39976
rect 23388 39924 23440 39976
rect 23664 39967 23716 39976
rect 23664 39933 23673 39967
rect 23673 39933 23707 39967
rect 23707 39933 23716 39967
rect 23664 39924 23716 39933
rect 28356 39992 28408 40044
rect 28724 39992 28776 40044
rect 25596 39924 25648 39976
rect 26332 39967 26384 39976
rect 26332 39933 26341 39967
rect 26341 39933 26375 39967
rect 26375 39933 26384 39967
rect 26332 39924 26384 39933
rect 26516 39924 26568 39976
rect 23572 39856 23624 39908
rect 25044 39856 25096 39908
rect 25228 39856 25280 39908
rect 22100 39831 22152 39840
rect 22100 39797 22109 39831
rect 22109 39797 22143 39831
rect 22143 39797 22152 39831
rect 22100 39788 22152 39797
rect 22744 39788 22796 39840
rect 22928 39788 22980 39840
rect 24216 39788 24268 39840
rect 24860 39788 24912 39840
rect 25412 39831 25464 39840
rect 25412 39797 25421 39831
rect 25421 39797 25455 39831
rect 25455 39797 25464 39831
rect 25412 39788 25464 39797
rect 27712 39788 27764 39840
rect 28540 39924 28592 39976
rect 29920 39924 29972 39976
rect 30564 39924 30616 39976
rect 31024 39967 31076 39976
rect 31024 39933 31033 39967
rect 31033 39933 31067 39967
rect 31067 39933 31076 39967
rect 31024 39924 31076 39933
rect 28356 39856 28408 39908
rect 28816 39899 28868 39908
rect 28816 39865 28825 39899
rect 28825 39865 28859 39899
rect 28859 39865 28868 39899
rect 28816 39856 28868 39865
rect 29276 39856 29328 39908
rect 28632 39831 28684 39840
rect 28632 39797 28659 39831
rect 28659 39797 28684 39831
rect 28632 39788 28684 39797
rect 29828 39831 29880 39840
rect 29828 39797 29837 39831
rect 29837 39797 29871 39831
rect 29871 39797 29880 39831
rect 29828 39788 29880 39797
rect 30380 39788 30432 39840
rect 4322 39686 4374 39738
rect 4386 39686 4438 39738
rect 4450 39686 4502 39738
rect 4514 39686 4566 39738
rect 4578 39686 4630 39738
rect 12096 39686 12148 39738
rect 12160 39686 12212 39738
rect 12224 39686 12276 39738
rect 12288 39686 12340 39738
rect 12352 39686 12404 39738
rect 19870 39686 19922 39738
rect 19934 39686 19986 39738
rect 19998 39686 20050 39738
rect 20062 39686 20114 39738
rect 20126 39686 20178 39738
rect 27644 39686 27696 39738
rect 27708 39686 27760 39738
rect 27772 39686 27824 39738
rect 27836 39686 27888 39738
rect 27900 39686 27952 39738
rect 9772 39584 9824 39636
rect 10692 39584 10744 39636
rect 8392 39448 8444 39500
rect 9772 39491 9824 39500
rect 9772 39457 9781 39491
rect 9781 39457 9815 39491
rect 9815 39457 9824 39491
rect 9772 39448 9824 39457
rect 10048 39516 10100 39568
rect 10968 39516 11020 39568
rect 9956 39491 10008 39500
rect 9956 39457 9965 39491
rect 9965 39457 9999 39491
rect 9999 39457 10008 39491
rect 9956 39448 10008 39457
rect 11612 39584 11664 39636
rect 11980 39516 12032 39568
rect 11704 39491 11756 39500
rect 11704 39457 11713 39491
rect 11713 39457 11747 39491
rect 11747 39457 11756 39491
rect 11704 39448 11756 39457
rect 11888 39491 11940 39500
rect 11888 39457 11897 39491
rect 11897 39457 11931 39491
rect 11931 39457 11940 39491
rect 11888 39448 11940 39457
rect 9220 39380 9272 39432
rect 11336 39380 11388 39432
rect 9772 39312 9824 39364
rect 12440 39584 12492 39636
rect 12532 39516 12584 39568
rect 12624 39491 12676 39500
rect 12624 39457 12633 39491
rect 12633 39457 12667 39491
rect 12667 39457 12676 39491
rect 12624 39448 12676 39457
rect 13452 39627 13504 39636
rect 13452 39593 13461 39627
rect 13461 39593 13495 39627
rect 13495 39593 13504 39627
rect 13452 39584 13504 39593
rect 13544 39584 13596 39636
rect 15476 39584 15528 39636
rect 17684 39584 17736 39636
rect 18972 39584 19024 39636
rect 12532 39380 12584 39432
rect 12624 39312 12676 39364
rect 9680 39244 9732 39296
rect 10416 39244 10468 39296
rect 11888 39244 11940 39296
rect 12440 39244 12492 39296
rect 12992 39491 13044 39500
rect 12992 39457 13001 39491
rect 13001 39457 13035 39491
rect 13035 39457 13044 39491
rect 12992 39448 13044 39457
rect 16488 39516 16540 39568
rect 17132 39516 17184 39568
rect 13636 39312 13688 39364
rect 13728 39312 13780 39364
rect 14924 39380 14976 39432
rect 15568 39448 15620 39500
rect 18512 39491 18564 39500
rect 18512 39457 18521 39491
rect 18521 39457 18555 39491
rect 18555 39457 18564 39491
rect 18512 39448 18564 39457
rect 18696 39491 18748 39500
rect 18696 39457 18705 39491
rect 18705 39457 18739 39491
rect 18739 39457 18748 39491
rect 18696 39448 18748 39457
rect 15844 39380 15896 39432
rect 18880 39491 18932 39500
rect 18880 39457 18889 39491
rect 18889 39457 18923 39491
rect 18923 39457 18932 39491
rect 18880 39448 18932 39457
rect 19248 39491 19300 39500
rect 19248 39457 19257 39491
rect 19257 39457 19291 39491
rect 19291 39457 19300 39491
rect 19248 39448 19300 39457
rect 19616 39448 19668 39500
rect 20168 39491 20220 39500
rect 20168 39457 20177 39491
rect 20177 39457 20211 39491
rect 20211 39457 20220 39491
rect 20168 39448 20220 39457
rect 20352 39491 20404 39500
rect 20352 39457 20361 39491
rect 20361 39457 20395 39491
rect 20395 39457 20404 39491
rect 20352 39448 20404 39457
rect 20444 39491 20496 39500
rect 20444 39457 20453 39491
rect 20453 39457 20487 39491
rect 20487 39457 20496 39491
rect 20444 39448 20496 39457
rect 22100 39516 22152 39568
rect 23572 39584 23624 39636
rect 25596 39627 25648 39636
rect 25596 39593 25605 39627
rect 25605 39593 25639 39627
rect 25639 39593 25648 39627
rect 25596 39584 25648 39593
rect 23204 39516 23256 39568
rect 26332 39516 26384 39568
rect 26792 39516 26844 39568
rect 17776 39312 17828 39364
rect 18880 39312 18932 39364
rect 20168 39312 20220 39364
rect 20628 39312 20680 39364
rect 22744 39491 22796 39500
rect 22744 39457 22753 39491
rect 22753 39457 22787 39491
rect 22787 39457 22796 39491
rect 22744 39448 22796 39457
rect 23572 39448 23624 39500
rect 24216 39491 24268 39500
rect 24216 39457 24225 39491
rect 24225 39457 24259 39491
rect 24259 39457 24268 39491
rect 24216 39448 24268 39457
rect 24492 39491 24544 39500
rect 24492 39457 24526 39491
rect 24526 39457 24544 39491
rect 24492 39448 24544 39457
rect 24860 39448 24912 39500
rect 26516 39380 26568 39432
rect 27344 39491 27396 39500
rect 27344 39457 27353 39491
rect 27353 39457 27387 39491
rect 27387 39457 27396 39491
rect 27344 39448 27396 39457
rect 28356 39448 28408 39500
rect 29460 39516 29512 39568
rect 29828 39491 29880 39500
rect 29828 39457 29837 39491
rect 29837 39457 29871 39491
rect 29871 39457 29880 39491
rect 29828 39448 29880 39457
rect 30196 39448 30248 39500
rect 25228 39312 25280 39364
rect 26884 39423 26936 39432
rect 26884 39389 26893 39423
rect 26893 39389 26927 39423
rect 26927 39389 26936 39423
rect 26884 39380 26936 39389
rect 28080 39380 28132 39432
rect 28540 39423 28592 39432
rect 28540 39389 28549 39423
rect 28549 39389 28583 39423
rect 28583 39389 28592 39423
rect 28540 39380 28592 39389
rect 28724 39380 28776 39432
rect 29552 39423 29604 39432
rect 29552 39389 29561 39423
rect 29561 39389 29595 39423
rect 29595 39389 29604 39423
rect 29552 39380 29604 39389
rect 29184 39312 29236 39364
rect 29920 39355 29972 39364
rect 29920 39321 29929 39355
rect 29929 39321 29963 39355
rect 29963 39321 29972 39355
rect 29920 39312 29972 39321
rect 13360 39244 13412 39296
rect 15384 39244 15436 39296
rect 18420 39244 18472 39296
rect 19248 39244 19300 39296
rect 19892 39287 19944 39296
rect 19892 39253 19901 39287
rect 19901 39253 19935 39287
rect 19935 39253 19944 39287
rect 19892 39244 19944 39253
rect 20444 39244 20496 39296
rect 21088 39244 21140 39296
rect 23848 39244 23900 39296
rect 25136 39244 25188 39296
rect 26056 39287 26108 39296
rect 26056 39253 26065 39287
rect 26065 39253 26099 39287
rect 26099 39253 26108 39287
rect 26056 39244 26108 39253
rect 26792 39244 26844 39296
rect 26884 39244 26936 39296
rect 27436 39244 27488 39296
rect 27712 39244 27764 39296
rect 28724 39244 28776 39296
rect 29644 39287 29696 39296
rect 29644 39253 29653 39287
rect 29653 39253 29687 39287
rect 29687 39253 29696 39287
rect 29644 39244 29696 39253
rect 30564 39244 30616 39296
rect 3662 39142 3714 39194
rect 3726 39142 3778 39194
rect 3790 39142 3842 39194
rect 3854 39142 3906 39194
rect 3918 39142 3970 39194
rect 11436 39142 11488 39194
rect 11500 39142 11552 39194
rect 11564 39142 11616 39194
rect 11628 39142 11680 39194
rect 11692 39142 11744 39194
rect 19210 39142 19262 39194
rect 19274 39142 19326 39194
rect 19338 39142 19390 39194
rect 19402 39142 19454 39194
rect 19466 39142 19518 39194
rect 26984 39142 27036 39194
rect 27048 39142 27100 39194
rect 27112 39142 27164 39194
rect 27176 39142 27228 39194
rect 27240 39142 27292 39194
rect 10600 39040 10652 39092
rect 10876 39040 10928 39092
rect 12532 39040 12584 39092
rect 12808 39040 12860 39092
rect 16948 39040 17000 39092
rect 18512 39040 18564 39092
rect 19432 39040 19484 39092
rect 20260 39040 20312 39092
rect 24492 39040 24544 39092
rect 24860 39040 24912 39092
rect 8300 38836 8352 38888
rect 9128 38879 9180 38888
rect 9128 38845 9137 38879
rect 9137 38845 9171 38879
rect 9171 38845 9180 38879
rect 9128 38836 9180 38845
rect 15568 38972 15620 39024
rect 9588 38904 9640 38956
rect 10968 38904 11020 38956
rect 13636 38904 13688 38956
rect 16948 38947 17000 38956
rect 16948 38913 16957 38947
rect 16957 38913 16991 38947
rect 16991 38913 17000 38947
rect 19524 38972 19576 39024
rect 19892 38972 19944 39024
rect 23480 38972 23532 39024
rect 25412 38972 25464 39024
rect 16948 38904 17000 38913
rect 9680 38836 9732 38888
rect 12440 38836 12492 38888
rect 15660 38836 15712 38888
rect 16212 38836 16264 38888
rect 16488 38836 16540 38888
rect 17224 38879 17276 38888
rect 17224 38845 17233 38879
rect 17233 38845 17267 38879
rect 17267 38845 17276 38879
rect 17224 38836 17276 38845
rect 17316 38836 17368 38888
rect 19800 38836 19852 38888
rect 10048 38768 10100 38820
rect 12716 38768 12768 38820
rect 12900 38768 12952 38820
rect 16948 38768 17000 38820
rect 18420 38768 18472 38820
rect 22928 38904 22980 38956
rect 25044 38836 25096 38888
rect 25228 38879 25280 38888
rect 25228 38845 25237 38879
rect 25237 38845 25271 38879
rect 25271 38845 25280 38879
rect 25228 38836 25280 38845
rect 26332 39040 26384 39092
rect 26608 39040 26660 39092
rect 27344 39040 27396 39092
rect 25596 38972 25648 39024
rect 25872 38947 25924 38956
rect 25872 38913 25881 38947
rect 25881 38913 25915 38947
rect 25915 38913 25924 38947
rect 25872 38904 25924 38913
rect 26608 38904 26660 38956
rect 26792 38904 26844 38956
rect 26424 38879 26476 38888
rect 26424 38845 26433 38879
rect 26433 38845 26467 38879
rect 26467 38845 26476 38879
rect 26424 38836 26476 38845
rect 29460 39040 29512 39092
rect 30196 39083 30248 39092
rect 30196 39049 30205 39083
rect 30205 39049 30239 39083
rect 30239 39049 30248 39083
rect 30196 39040 30248 39049
rect 28908 38972 28960 39024
rect 29276 38836 29328 38888
rect 29644 38836 29696 38888
rect 30380 38879 30432 38888
rect 30380 38845 30389 38879
rect 30389 38845 30423 38879
rect 30423 38845 30432 38879
rect 30380 38836 30432 38845
rect 20352 38768 20404 38820
rect 8484 38743 8536 38752
rect 8484 38709 8493 38743
rect 8493 38709 8527 38743
rect 8527 38709 8536 38743
rect 8484 38700 8536 38709
rect 9864 38700 9916 38752
rect 14096 38700 14148 38752
rect 15476 38700 15528 38752
rect 16212 38743 16264 38752
rect 16212 38709 16221 38743
rect 16221 38709 16255 38743
rect 16255 38709 16264 38743
rect 16212 38700 16264 38709
rect 16672 38700 16724 38752
rect 16856 38743 16908 38752
rect 16856 38709 16865 38743
rect 16865 38709 16899 38743
rect 16899 38709 16908 38743
rect 16856 38700 16908 38709
rect 19708 38700 19760 38752
rect 20168 38743 20220 38752
rect 20168 38709 20177 38743
rect 20177 38709 20211 38743
rect 20211 38709 20220 38743
rect 20168 38700 20220 38709
rect 23848 38700 23900 38752
rect 26424 38700 26476 38752
rect 28080 38768 28132 38820
rect 29184 38768 29236 38820
rect 26976 38700 27028 38752
rect 28816 38700 28868 38752
rect 30564 38768 30616 38820
rect 4322 38598 4374 38650
rect 4386 38598 4438 38650
rect 4450 38598 4502 38650
rect 4514 38598 4566 38650
rect 4578 38598 4630 38650
rect 12096 38598 12148 38650
rect 12160 38598 12212 38650
rect 12224 38598 12276 38650
rect 12288 38598 12340 38650
rect 12352 38598 12404 38650
rect 19870 38598 19922 38650
rect 19934 38598 19986 38650
rect 19998 38598 20050 38650
rect 20062 38598 20114 38650
rect 20126 38598 20178 38650
rect 27644 38598 27696 38650
rect 27708 38598 27760 38650
rect 27772 38598 27824 38650
rect 27836 38598 27888 38650
rect 27900 38598 27952 38650
rect 9588 38496 9640 38548
rect 15108 38496 15160 38548
rect 15660 38496 15712 38548
rect 16396 38496 16448 38548
rect 8484 38428 8536 38480
rect 11336 38428 11388 38480
rect 9864 38403 9916 38412
rect 9864 38369 9873 38403
rect 9873 38369 9907 38403
rect 9907 38369 9916 38403
rect 9864 38360 9916 38369
rect 10048 38403 10100 38412
rect 10048 38369 10057 38403
rect 10057 38369 10091 38403
rect 10091 38369 10100 38403
rect 10048 38360 10100 38369
rect 10232 38403 10284 38412
rect 10232 38369 10241 38403
rect 10241 38369 10275 38403
rect 10275 38369 10284 38403
rect 10232 38360 10284 38369
rect 11888 38428 11940 38480
rect 13452 38428 13504 38480
rect 10508 38292 10560 38344
rect 10968 38292 11020 38344
rect 9864 38224 9916 38276
rect 10232 38224 10284 38276
rect 12440 38403 12492 38412
rect 12440 38369 12449 38403
rect 12449 38369 12483 38403
rect 12483 38369 12492 38403
rect 12440 38360 12492 38369
rect 13268 38335 13320 38344
rect 13268 38301 13277 38335
rect 13277 38301 13311 38335
rect 13311 38301 13320 38335
rect 13268 38292 13320 38301
rect 13820 38403 13872 38412
rect 13820 38369 13829 38403
rect 13829 38369 13863 38403
rect 13863 38369 13872 38403
rect 13820 38360 13872 38369
rect 15200 38428 15252 38480
rect 14096 38403 14148 38412
rect 14096 38369 14105 38403
rect 14105 38369 14139 38403
rect 14139 38369 14148 38403
rect 14096 38360 14148 38369
rect 14924 38360 14976 38412
rect 16028 38360 16080 38412
rect 16212 38360 16264 38412
rect 17684 38360 17736 38412
rect 12992 38224 13044 38276
rect 15936 38292 15988 38344
rect 17500 38292 17552 38344
rect 18420 38360 18472 38412
rect 22284 38496 22336 38548
rect 23572 38539 23624 38548
rect 23572 38505 23581 38539
rect 23581 38505 23615 38539
rect 23615 38505 23624 38539
rect 23572 38496 23624 38505
rect 28540 38496 28592 38548
rect 19064 38360 19116 38412
rect 16120 38224 16172 38276
rect 10140 38156 10192 38208
rect 10324 38156 10376 38208
rect 11244 38156 11296 38208
rect 12716 38156 12768 38208
rect 14188 38199 14240 38208
rect 14188 38165 14197 38199
rect 14197 38165 14231 38199
rect 14231 38165 14240 38199
rect 14188 38156 14240 38165
rect 14372 38199 14424 38208
rect 14372 38165 14381 38199
rect 14381 38165 14415 38199
rect 14415 38165 14424 38199
rect 14372 38156 14424 38165
rect 15660 38199 15712 38208
rect 15660 38165 15669 38199
rect 15669 38165 15703 38199
rect 15703 38165 15712 38199
rect 15660 38156 15712 38165
rect 15752 38156 15804 38208
rect 17868 38156 17920 38208
rect 18972 38335 19024 38344
rect 18972 38301 18981 38335
rect 18981 38301 19015 38335
rect 19015 38301 19024 38335
rect 18972 38292 19024 38301
rect 19708 38403 19760 38412
rect 19708 38369 19717 38403
rect 19717 38369 19751 38403
rect 19751 38369 19760 38403
rect 19708 38360 19760 38369
rect 20812 38428 20864 38480
rect 25136 38428 25188 38480
rect 27988 38428 28040 38480
rect 19984 38403 20036 38412
rect 19984 38369 20018 38403
rect 20018 38369 20036 38403
rect 19984 38360 20036 38369
rect 20536 38360 20588 38412
rect 22376 38360 22428 38412
rect 23756 38403 23808 38412
rect 23756 38369 23765 38403
rect 23765 38369 23799 38403
rect 23799 38369 23808 38403
rect 23756 38360 23808 38369
rect 26884 38360 26936 38412
rect 29276 38360 29328 38412
rect 23940 38335 23992 38344
rect 23940 38301 23949 38335
rect 23949 38301 23983 38335
rect 23983 38301 23992 38335
rect 23940 38292 23992 38301
rect 22836 38224 22888 38276
rect 20904 38156 20956 38208
rect 22192 38156 22244 38208
rect 29092 38156 29144 38208
rect 3662 38054 3714 38106
rect 3726 38054 3778 38106
rect 3790 38054 3842 38106
rect 3854 38054 3906 38106
rect 3918 38054 3970 38106
rect 11436 38054 11488 38106
rect 11500 38054 11552 38106
rect 11564 38054 11616 38106
rect 11628 38054 11680 38106
rect 11692 38054 11744 38106
rect 19210 38054 19262 38106
rect 19274 38054 19326 38106
rect 19338 38054 19390 38106
rect 19402 38054 19454 38106
rect 19466 38054 19518 38106
rect 26984 38054 27036 38106
rect 27048 38054 27100 38106
rect 27112 38054 27164 38106
rect 27176 38054 27228 38106
rect 27240 38054 27292 38106
rect 9680 37995 9732 38004
rect 9680 37961 9689 37995
rect 9689 37961 9723 37995
rect 9723 37961 9732 37995
rect 9680 37952 9732 37961
rect 8300 37884 8352 37936
rect 10140 37859 10192 37868
rect 10140 37825 10149 37859
rect 10149 37825 10183 37859
rect 10183 37825 10192 37859
rect 10140 37816 10192 37825
rect 10324 37859 10376 37868
rect 10324 37825 10333 37859
rect 10333 37825 10367 37859
rect 10367 37825 10376 37859
rect 10324 37816 10376 37825
rect 12440 37952 12492 38004
rect 13084 37952 13136 38004
rect 14924 37952 14976 38004
rect 15936 37995 15988 38004
rect 15936 37961 15945 37995
rect 15945 37961 15979 37995
rect 15979 37961 15988 37995
rect 15936 37952 15988 37961
rect 16856 37952 16908 38004
rect 9496 37748 9548 37800
rect 10876 37791 10928 37800
rect 10876 37757 10885 37791
rect 10885 37757 10919 37791
rect 10919 37757 10928 37791
rect 10876 37748 10928 37757
rect 11244 37748 11296 37800
rect 12900 37884 12952 37936
rect 16488 37884 16540 37936
rect 18052 37952 18104 38004
rect 18880 37952 18932 38004
rect 19984 37952 20036 38004
rect 20444 37952 20496 38004
rect 20720 37952 20772 38004
rect 17684 37884 17736 37936
rect 23296 37952 23348 38004
rect 24032 37952 24084 38004
rect 25872 37952 25924 38004
rect 12716 37791 12768 37800
rect 12716 37757 12725 37791
rect 12725 37757 12759 37791
rect 12759 37757 12768 37791
rect 12716 37748 12768 37757
rect 12808 37748 12860 37800
rect 12992 37791 13044 37800
rect 12992 37757 13001 37791
rect 13001 37757 13035 37791
rect 13035 37757 13044 37791
rect 12992 37748 13044 37757
rect 17868 37859 17920 37868
rect 17868 37825 17877 37859
rect 17877 37825 17911 37859
rect 17911 37825 17920 37859
rect 17868 37816 17920 37825
rect 19340 37859 19392 37868
rect 19340 37825 19349 37859
rect 19349 37825 19383 37859
rect 19383 37825 19392 37859
rect 19340 37816 19392 37825
rect 15384 37748 15436 37800
rect 15476 37791 15528 37800
rect 15476 37757 15485 37791
rect 15485 37757 15519 37791
rect 15519 37757 15528 37791
rect 15476 37748 15528 37757
rect 15568 37791 15620 37800
rect 15568 37757 15577 37791
rect 15577 37757 15611 37791
rect 15611 37757 15620 37791
rect 15568 37748 15620 37757
rect 15844 37748 15896 37800
rect 16212 37748 16264 37800
rect 16948 37791 17000 37800
rect 16948 37757 16957 37791
rect 16957 37757 16991 37791
rect 16991 37757 17000 37791
rect 16948 37748 17000 37757
rect 9496 37612 9548 37664
rect 10600 37612 10652 37664
rect 13912 37680 13964 37732
rect 14188 37680 14240 37732
rect 16396 37680 16448 37732
rect 16856 37612 16908 37664
rect 17868 37612 17920 37664
rect 18328 37748 18380 37800
rect 18972 37791 19024 37800
rect 18972 37757 18981 37791
rect 18981 37757 19015 37791
rect 19015 37757 19024 37791
rect 18972 37748 19024 37757
rect 19800 37816 19852 37868
rect 20076 37791 20128 37800
rect 20076 37757 20085 37791
rect 20085 37757 20119 37791
rect 20119 37757 20128 37791
rect 20076 37748 20128 37757
rect 20168 37791 20220 37800
rect 20168 37757 20177 37791
rect 20177 37757 20211 37791
rect 20211 37757 20220 37791
rect 20168 37748 20220 37757
rect 20352 37748 20404 37800
rect 18788 37723 18840 37732
rect 18788 37689 18797 37723
rect 18797 37689 18831 37723
rect 18831 37689 18840 37723
rect 18788 37680 18840 37689
rect 18880 37723 18932 37732
rect 18880 37689 18889 37723
rect 18889 37689 18923 37723
rect 18923 37689 18932 37723
rect 18880 37680 18932 37689
rect 19616 37680 19668 37732
rect 20536 37748 20588 37800
rect 20904 37791 20956 37800
rect 20904 37757 20913 37791
rect 20913 37757 20947 37791
rect 20947 37757 20956 37791
rect 20904 37748 20956 37757
rect 21272 37816 21324 37868
rect 22192 37859 22244 37868
rect 22192 37825 22201 37859
rect 22201 37825 22235 37859
rect 22235 37825 22244 37859
rect 22192 37816 22244 37825
rect 29092 37859 29144 37868
rect 29092 37825 29101 37859
rect 29101 37825 29135 37859
rect 29135 37825 29144 37859
rect 29092 37816 29144 37825
rect 22284 37748 22336 37800
rect 24952 37791 25004 37800
rect 24952 37757 24961 37791
rect 24961 37757 24995 37791
rect 24995 37757 25004 37791
rect 24952 37748 25004 37757
rect 31116 37816 31168 37868
rect 21640 37723 21692 37732
rect 21640 37689 21649 37723
rect 21649 37689 21683 37723
rect 21683 37689 21692 37723
rect 21640 37680 21692 37689
rect 23388 37680 23440 37732
rect 19524 37612 19576 37664
rect 20628 37655 20680 37664
rect 20628 37621 20637 37655
rect 20637 37621 20671 37655
rect 20671 37621 20680 37655
rect 20628 37612 20680 37621
rect 21824 37612 21876 37664
rect 30472 37655 30524 37664
rect 30472 37621 30481 37655
rect 30481 37621 30515 37655
rect 30515 37621 30524 37655
rect 30472 37612 30524 37621
rect 4322 37510 4374 37562
rect 4386 37510 4438 37562
rect 4450 37510 4502 37562
rect 4514 37510 4566 37562
rect 4578 37510 4630 37562
rect 12096 37510 12148 37562
rect 12160 37510 12212 37562
rect 12224 37510 12276 37562
rect 12288 37510 12340 37562
rect 12352 37510 12404 37562
rect 19870 37510 19922 37562
rect 19934 37510 19986 37562
rect 19998 37510 20050 37562
rect 20062 37510 20114 37562
rect 20126 37510 20178 37562
rect 27644 37510 27696 37562
rect 27708 37510 27760 37562
rect 27772 37510 27824 37562
rect 27836 37510 27888 37562
rect 27900 37510 27952 37562
rect 9128 37408 9180 37460
rect 9128 37315 9180 37324
rect 9128 37281 9137 37315
rect 9137 37281 9171 37315
rect 9171 37281 9180 37315
rect 9128 37272 9180 37281
rect 9956 37408 10008 37460
rect 10416 37408 10468 37460
rect 14372 37408 14424 37460
rect 15660 37408 15712 37460
rect 16488 37408 16540 37460
rect 20352 37451 20404 37460
rect 20352 37417 20361 37451
rect 20361 37417 20395 37451
rect 20395 37417 20404 37451
rect 20352 37408 20404 37417
rect 9772 37340 9824 37392
rect 10876 37340 10928 37392
rect 9496 37315 9548 37324
rect 9496 37281 9505 37315
rect 9505 37281 9539 37315
rect 9539 37281 9548 37315
rect 9496 37272 9548 37281
rect 10140 37315 10192 37324
rect 10140 37281 10149 37315
rect 10149 37281 10183 37315
rect 10183 37281 10192 37315
rect 10140 37272 10192 37281
rect 10324 37315 10376 37324
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 10416 37272 10468 37324
rect 14556 37272 14608 37324
rect 15200 37272 15252 37324
rect 16396 37272 16448 37324
rect 15292 37204 15344 37256
rect 15660 37204 15712 37256
rect 15108 37136 15160 37188
rect 16948 37315 17000 37324
rect 16948 37281 16957 37315
rect 16957 37281 16991 37315
rect 16991 37281 17000 37315
rect 16948 37272 17000 37281
rect 18880 37340 18932 37392
rect 19340 37204 19392 37256
rect 20168 37315 20220 37324
rect 20168 37281 20177 37315
rect 20177 37281 20211 37315
rect 20211 37281 20220 37315
rect 20168 37272 20220 37281
rect 20720 37315 20772 37324
rect 20720 37281 20729 37315
rect 20729 37281 20763 37315
rect 20763 37281 20772 37315
rect 20720 37272 20772 37281
rect 20444 37204 20496 37256
rect 20536 37204 20588 37256
rect 20904 37315 20956 37324
rect 20904 37281 20913 37315
rect 20913 37281 20947 37315
rect 20947 37281 20956 37315
rect 20904 37272 20956 37281
rect 21088 37315 21140 37324
rect 21088 37281 21097 37315
rect 21097 37281 21131 37315
rect 21131 37281 21140 37315
rect 21088 37272 21140 37281
rect 21272 37315 21324 37324
rect 21272 37281 21281 37315
rect 21281 37281 21315 37315
rect 21315 37281 21324 37315
rect 21272 37272 21324 37281
rect 21640 37408 21692 37460
rect 23388 37451 23440 37460
rect 23388 37417 23397 37451
rect 23397 37417 23431 37451
rect 23431 37417 23440 37451
rect 23388 37408 23440 37417
rect 23480 37340 23532 37392
rect 24952 37340 25004 37392
rect 29000 37408 29052 37460
rect 30472 37408 30524 37460
rect 30564 37408 30616 37460
rect 31300 37408 31352 37460
rect 22376 37272 22428 37324
rect 23572 37315 23624 37324
rect 23572 37281 23581 37315
rect 23581 37281 23615 37315
rect 23615 37281 23624 37315
rect 23572 37272 23624 37281
rect 23664 37272 23716 37324
rect 24584 37315 24636 37324
rect 24584 37281 24593 37315
rect 24593 37281 24627 37315
rect 24627 37281 24636 37315
rect 24584 37272 24636 37281
rect 25136 37272 25188 37324
rect 27344 37340 27396 37392
rect 26884 37315 26936 37324
rect 26884 37281 26893 37315
rect 26893 37281 26927 37315
rect 26927 37281 26936 37315
rect 26884 37272 26936 37281
rect 29000 37315 29052 37324
rect 29000 37281 29018 37315
rect 29018 37281 29052 37315
rect 29000 37272 29052 37281
rect 29092 37315 29144 37324
rect 29092 37281 29101 37315
rect 29101 37281 29135 37315
rect 29135 37281 29144 37315
rect 29092 37272 29144 37281
rect 30196 37272 30248 37324
rect 22928 37204 22980 37256
rect 9312 37068 9364 37120
rect 10692 37111 10744 37120
rect 10692 37077 10701 37111
rect 10701 37077 10735 37111
rect 10735 37077 10744 37111
rect 10692 37068 10744 37077
rect 13728 37111 13780 37120
rect 13728 37077 13737 37111
rect 13737 37077 13771 37111
rect 13771 37077 13780 37111
rect 13728 37068 13780 37077
rect 15568 37111 15620 37120
rect 15568 37077 15577 37111
rect 15577 37077 15611 37111
rect 15611 37077 15620 37111
rect 15568 37068 15620 37077
rect 18328 37068 18380 37120
rect 18972 37136 19024 37188
rect 20628 37136 20680 37188
rect 23296 37136 23348 37188
rect 26700 37204 26752 37256
rect 28264 37204 28316 37256
rect 28816 37247 28868 37256
rect 28816 37213 28825 37247
rect 28825 37213 28859 37247
rect 28859 37213 28868 37247
rect 28816 37204 28868 37213
rect 26884 37136 26936 37188
rect 27436 37136 27488 37188
rect 18604 37111 18656 37120
rect 18604 37077 18613 37111
rect 18613 37077 18647 37111
rect 18647 37077 18656 37111
rect 18604 37068 18656 37077
rect 23480 37068 23532 37120
rect 24952 37068 25004 37120
rect 25872 37068 25924 37120
rect 26792 37068 26844 37120
rect 27804 37068 27856 37120
rect 28724 37068 28776 37120
rect 29460 37068 29512 37120
rect 30748 37247 30800 37256
rect 30748 37213 30757 37247
rect 30757 37213 30791 37247
rect 30791 37213 30800 37247
rect 30748 37204 30800 37213
rect 31300 37315 31352 37324
rect 31300 37281 31309 37315
rect 31309 37281 31343 37315
rect 31343 37281 31352 37315
rect 31300 37272 31352 37281
rect 30288 37136 30340 37188
rect 31024 37136 31076 37188
rect 31116 37179 31168 37188
rect 31116 37145 31125 37179
rect 31125 37145 31159 37179
rect 31159 37145 31168 37179
rect 31116 37136 31168 37145
rect 30564 37068 30616 37120
rect 3662 36966 3714 37018
rect 3726 36966 3778 37018
rect 3790 36966 3842 37018
rect 3854 36966 3906 37018
rect 3918 36966 3970 37018
rect 11436 36966 11488 37018
rect 11500 36966 11552 37018
rect 11564 36966 11616 37018
rect 11628 36966 11680 37018
rect 11692 36966 11744 37018
rect 19210 36966 19262 37018
rect 19274 36966 19326 37018
rect 19338 36966 19390 37018
rect 19402 36966 19454 37018
rect 19466 36966 19518 37018
rect 26984 36966 27036 37018
rect 27048 36966 27100 37018
rect 27112 36966 27164 37018
rect 27176 36966 27228 37018
rect 27240 36966 27292 37018
rect 10140 36864 10192 36916
rect 8300 36728 8352 36780
rect 12900 36864 12952 36916
rect 13268 36864 13320 36916
rect 14556 36864 14608 36916
rect 15108 36907 15160 36916
rect 15108 36873 15117 36907
rect 15117 36873 15151 36907
rect 15151 36873 15160 36907
rect 15108 36864 15160 36873
rect 16212 36907 16264 36916
rect 16212 36873 16221 36907
rect 16221 36873 16255 36907
rect 16255 36873 16264 36907
rect 16212 36864 16264 36873
rect 17868 36907 17920 36916
rect 17868 36873 17877 36907
rect 17877 36873 17911 36907
rect 17911 36873 17920 36907
rect 17868 36864 17920 36873
rect 18972 36907 19024 36916
rect 18972 36873 18981 36907
rect 18981 36873 19015 36907
rect 19015 36873 19024 36907
rect 18972 36864 19024 36873
rect 20720 36864 20772 36916
rect 13820 36839 13872 36848
rect 13820 36805 13829 36839
rect 13829 36805 13863 36839
rect 13863 36805 13872 36839
rect 13820 36796 13872 36805
rect 15660 36796 15712 36848
rect 16120 36796 16172 36848
rect 20904 36864 20956 36916
rect 21088 36864 21140 36916
rect 22928 36864 22980 36916
rect 23572 36864 23624 36916
rect 27344 36864 27396 36916
rect 30288 36864 30340 36916
rect 14556 36771 14608 36780
rect 14556 36737 14565 36771
rect 14565 36737 14599 36771
rect 14599 36737 14608 36771
rect 14556 36728 14608 36737
rect 9588 36660 9640 36712
rect 9036 36592 9088 36644
rect 10416 36635 10468 36644
rect 10416 36601 10425 36635
rect 10425 36601 10459 36635
rect 10459 36601 10468 36635
rect 10416 36592 10468 36601
rect 11244 36703 11296 36712
rect 11244 36669 11253 36703
rect 11253 36669 11287 36703
rect 11287 36669 11296 36703
rect 11244 36660 11296 36669
rect 11428 36703 11480 36712
rect 11428 36669 11437 36703
rect 11437 36669 11471 36703
rect 11471 36669 11480 36703
rect 11428 36660 11480 36669
rect 11060 36592 11112 36644
rect 12624 36660 12676 36712
rect 15568 36728 15620 36780
rect 14188 36592 14240 36644
rect 10968 36567 11020 36576
rect 10968 36533 10977 36567
rect 10977 36533 11011 36567
rect 11011 36533 11020 36567
rect 10968 36524 11020 36533
rect 12992 36524 13044 36576
rect 14556 36524 14608 36576
rect 15660 36660 15712 36712
rect 16028 36660 16080 36712
rect 16396 36771 16448 36780
rect 16396 36737 16405 36771
rect 16405 36737 16439 36771
rect 16439 36737 16448 36771
rect 16396 36728 16448 36737
rect 18696 36728 18748 36780
rect 16212 36592 16264 36644
rect 16488 36703 16540 36712
rect 16488 36669 16497 36703
rect 16497 36669 16531 36703
rect 16531 36669 16540 36703
rect 16488 36660 16540 36669
rect 19064 36728 19116 36780
rect 22836 36728 22888 36780
rect 17960 36592 18012 36644
rect 15568 36524 15620 36576
rect 16120 36524 16172 36576
rect 18144 36524 18196 36576
rect 18788 36592 18840 36644
rect 19248 36703 19300 36712
rect 19248 36669 19257 36703
rect 19257 36669 19291 36703
rect 19291 36669 19300 36703
rect 19248 36660 19300 36669
rect 18972 36592 19024 36644
rect 21456 36660 21508 36712
rect 21916 36660 21968 36712
rect 23020 36703 23072 36712
rect 23020 36669 23029 36703
rect 23029 36669 23063 36703
rect 23063 36669 23072 36703
rect 23020 36660 23072 36669
rect 23940 36771 23992 36780
rect 23940 36737 23949 36771
rect 23949 36737 23983 36771
rect 23983 36737 23992 36771
rect 23940 36728 23992 36737
rect 23664 36660 23716 36712
rect 24124 36703 24176 36712
rect 24124 36669 24133 36703
rect 24133 36669 24167 36703
rect 24167 36669 24176 36703
rect 24124 36660 24176 36669
rect 24400 36703 24452 36712
rect 24400 36669 24409 36703
rect 24409 36669 24443 36703
rect 24443 36669 24452 36703
rect 24400 36660 24452 36669
rect 25872 36771 25924 36780
rect 25872 36737 25881 36771
rect 25881 36737 25915 36771
rect 25915 36737 25924 36771
rect 25872 36728 25924 36737
rect 27804 36771 27856 36780
rect 27804 36737 27813 36771
rect 27813 36737 27847 36771
rect 27847 36737 27856 36771
rect 27804 36728 27856 36737
rect 29184 36703 29236 36712
rect 29184 36669 29193 36703
rect 29193 36669 29227 36703
rect 29227 36669 29236 36703
rect 29184 36660 29236 36669
rect 20352 36635 20404 36644
rect 20352 36601 20361 36635
rect 20361 36601 20395 36635
rect 20395 36601 20404 36635
rect 20352 36592 20404 36601
rect 20536 36635 20588 36644
rect 20536 36601 20545 36635
rect 20545 36601 20579 36635
rect 20579 36601 20588 36635
rect 20536 36592 20588 36601
rect 20628 36635 20680 36644
rect 20628 36601 20637 36635
rect 20637 36601 20671 36635
rect 20671 36601 20680 36635
rect 20628 36592 20680 36601
rect 20812 36635 20864 36644
rect 20812 36601 20821 36635
rect 20821 36601 20855 36635
rect 20855 36601 20864 36635
rect 20812 36592 20864 36601
rect 20260 36524 20312 36576
rect 24032 36592 24084 36644
rect 24768 36592 24820 36644
rect 25228 36592 25280 36644
rect 26608 36592 26660 36644
rect 23480 36524 23532 36576
rect 25780 36567 25832 36576
rect 25780 36533 25789 36567
rect 25789 36533 25823 36567
rect 25823 36533 25832 36567
rect 25780 36524 25832 36533
rect 29460 36635 29512 36644
rect 29460 36601 29469 36635
rect 29469 36601 29503 36635
rect 29503 36601 29512 36635
rect 29460 36592 29512 36601
rect 30012 36592 30064 36644
rect 28080 36524 28132 36576
rect 29644 36567 29696 36576
rect 29644 36533 29669 36567
rect 29669 36533 29696 36567
rect 29644 36524 29696 36533
rect 30564 36524 30616 36576
rect 4322 36422 4374 36474
rect 4386 36422 4438 36474
rect 4450 36422 4502 36474
rect 4514 36422 4566 36474
rect 4578 36422 4630 36474
rect 12096 36422 12148 36474
rect 12160 36422 12212 36474
rect 12224 36422 12276 36474
rect 12288 36422 12340 36474
rect 12352 36422 12404 36474
rect 19870 36422 19922 36474
rect 19934 36422 19986 36474
rect 19998 36422 20050 36474
rect 20062 36422 20114 36474
rect 20126 36422 20178 36474
rect 27644 36422 27696 36474
rect 27708 36422 27760 36474
rect 27772 36422 27824 36474
rect 27836 36422 27888 36474
rect 27900 36422 27952 36474
rect 9036 36363 9088 36372
rect 9036 36329 9045 36363
rect 9045 36329 9079 36363
rect 9079 36329 9088 36363
rect 9036 36320 9088 36329
rect 9312 36227 9364 36236
rect 9312 36193 9321 36227
rect 9321 36193 9355 36227
rect 9355 36193 9364 36227
rect 9312 36184 9364 36193
rect 9864 36320 9916 36372
rect 11428 36320 11480 36372
rect 13176 36363 13228 36372
rect 13176 36329 13185 36363
rect 13185 36329 13219 36363
rect 13219 36329 13228 36363
rect 13176 36320 13228 36329
rect 14556 36363 14608 36372
rect 14556 36329 14565 36363
rect 14565 36329 14599 36363
rect 14599 36329 14608 36363
rect 14556 36320 14608 36329
rect 16028 36320 16080 36372
rect 17960 36320 18012 36372
rect 18972 36320 19024 36372
rect 10968 36252 11020 36304
rect 11244 36252 11296 36304
rect 10232 36184 10284 36236
rect 9588 36116 9640 36168
rect 10508 36227 10560 36236
rect 10508 36193 10517 36227
rect 10517 36193 10551 36227
rect 10551 36193 10560 36227
rect 10508 36184 10560 36193
rect 10692 36227 10744 36236
rect 10692 36193 10701 36227
rect 10701 36193 10735 36227
rect 10735 36193 10744 36227
rect 10692 36184 10744 36193
rect 11980 36227 12032 36236
rect 11980 36193 11989 36227
rect 11989 36193 12023 36227
rect 12023 36193 12032 36227
rect 11980 36184 12032 36193
rect 12164 36184 12216 36236
rect 11244 36116 11296 36168
rect 11520 36116 11572 36168
rect 11888 36116 11940 36168
rect 12624 36184 12676 36236
rect 12808 36184 12860 36236
rect 12900 36227 12952 36236
rect 12900 36193 12909 36227
rect 12909 36193 12943 36227
rect 12943 36193 12952 36227
rect 12900 36184 12952 36193
rect 12716 36116 12768 36168
rect 13820 36184 13872 36236
rect 14280 36116 14332 36168
rect 15476 36184 15528 36236
rect 16212 36184 16264 36236
rect 18880 36252 18932 36304
rect 20444 36320 20496 36372
rect 20628 36320 20680 36372
rect 23480 36320 23532 36372
rect 23756 36320 23808 36372
rect 24124 36320 24176 36372
rect 24400 36320 24452 36372
rect 19616 36252 19668 36304
rect 16396 36184 16448 36236
rect 15292 36116 15344 36168
rect 11888 35980 11940 36032
rect 13636 36091 13688 36100
rect 13636 36057 13645 36091
rect 13645 36057 13679 36091
rect 13679 36057 13688 36091
rect 13636 36048 13688 36057
rect 14004 36048 14056 36100
rect 16488 36116 16540 36168
rect 16856 36227 16908 36236
rect 16856 36193 16865 36227
rect 16865 36193 16899 36227
rect 16899 36193 16908 36227
rect 16856 36184 16908 36193
rect 17960 36227 18012 36236
rect 17960 36193 17969 36227
rect 17969 36193 18003 36227
rect 18003 36193 18012 36227
rect 17960 36184 18012 36193
rect 18420 36227 18472 36236
rect 18420 36193 18429 36227
rect 18429 36193 18463 36227
rect 18463 36193 18472 36227
rect 18420 36184 18472 36193
rect 18788 36184 18840 36236
rect 18144 36116 18196 36168
rect 18328 36116 18380 36168
rect 18512 36116 18564 36168
rect 19248 36116 19300 36168
rect 20260 36227 20312 36236
rect 20260 36193 20269 36227
rect 20269 36193 20303 36227
rect 20303 36193 20312 36227
rect 20260 36184 20312 36193
rect 12624 36023 12676 36032
rect 12624 35989 12633 36023
rect 12633 35989 12667 36023
rect 12667 35989 12676 36023
rect 12624 35980 12676 35989
rect 13912 35980 13964 36032
rect 14740 35980 14792 36032
rect 16396 36023 16448 36032
rect 16396 35989 16405 36023
rect 16405 35989 16439 36023
rect 16439 35989 16448 36023
rect 16396 35980 16448 35989
rect 16488 35980 16540 36032
rect 19524 36048 19576 36100
rect 18696 35980 18748 36032
rect 18972 35980 19024 36032
rect 20812 36184 20864 36236
rect 21548 36227 21600 36236
rect 21548 36193 21557 36227
rect 21557 36193 21591 36227
rect 21591 36193 21600 36227
rect 21548 36184 21600 36193
rect 22376 36184 22428 36236
rect 22560 36227 22612 36236
rect 22560 36193 22569 36227
rect 22569 36193 22603 36227
rect 22603 36193 22612 36227
rect 22560 36184 22612 36193
rect 23480 36227 23532 36236
rect 23480 36193 23489 36227
rect 23489 36193 23523 36227
rect 23523 36193 23532 36227
rect 23480 36184 23532 36193
rect 23204 36159 23256 36168
rect 23204 36125 23213 36159
rect 23213 36125 23247 36159
rect 23247 36125 23256 36159
rect 23204 36116 23256 36125
rect 23664 36227 23716 36236
rect 23664 36193 23673 36227
rect 23673 36193 23707 36227
rect 23707 36193 23716 36227
rect 23664 36184 23716 36193
rect 25228 36252 25280 36304
rect 25780 36252 25832 36304
rect 26700 36320 26752 36372
rect 30012 36363 30064 36372
rect 30012 36329 30021 36363
rect 30021 36329 30055 36363
rect 30055 36329 30064 36363
rect 30012 36320 30064 36329
rect 30288 36320 30340 36372
rect 24124 36184 24176 36236
rect 23848 36116 23900 36168
rect 24032 36159 24084 36168
rect 24032 36125 24041 36159
rect 24041 36125 24075 36159
rect 24075 36125 24084 36159
rect 24032 36116 24084 36125
rect 22284 36091 22336 36100
rect 22284 36057 22293 36091
rect 22293 36057 22327 36091
rect 22327 36057 22336 36091
rect 22284 36048 22336 36057
rect 22836 36048 22888 36100
rect 24584 36184 24636 36236
rect 24768 36227 24820 36236
rect 24768 36193 24777 36227
rect 24777 36193 24811 36227
rect 24811 36193 24820 36227
rect 24768 36184 24820 36193
rect 24952 36227 25004 36236
rect 24952 36193 24961 36227
rect 24961 36193 24995 36227
rect 24995 36193 25004 36227
rect 24952 36184 25004 36193
rect 25412 36227 25464 36236
rect 25412 36193 25421 36227
rect 25421 36193 25455 36227
rect 25455 36193 25464 36227
rect 25412 36184 25464 36193
rect 31024 36363 31076 36372
rect 31024 36329 31033 36363
rect 31033 36329 31067 36363
rect 31067 36329 31076 36363
rect 31024 36320 31076 36329
rect 31300 36320 31352 36372
rect 26424 36227 26476 36236
rect 26424 36193 26433 36227
rect 26433 36193 26467 36227
rect 26467 36193 26476 36227
rect 26424 36184 26476 36193
rect 26608 36227 26660 36236
rect 26608 36193 26616 36227
rect 26616 36193 26650 36227
rect 26650 36193 26660 36227
rect 26608 36184 26660 36193
rect 26700 36227 26752 36236
rect 26700 36193 26709 36227
rect 26709 36193 26743 36227
rect 26743 36193 26752 36227
rect 26700 36184 26752 36193
rect 26792 36227 26844 36236
rect 26792 36193 26801 36227
rect 26801 36193 26835 36227
rect 26835 36193 26844 36227
rect 26792 36184 26844 36193
rect 26884 36184 26936 36236
rect 30564 36227 30616 36236
rect 30564 36193 30573 36227
rect 30573 36193 30607 36227
rect 30607 36193 30616 36227
rect 30564 36184 30616 36193
rect 29644 36116 29696 36168
rect 30288 36116 30340 36168
rect 20628 36023 20680 36032
rect 20628 35989 20637 36023
rect 20637 35989 20671 36023
rect 20671 35989 20680 36023
rect 20628 35980 20680 35989
rect 21456 35980 21508 36032
rect 21824 35980 21876 36032
rect 25688 36023 25740 36032
rect 25688 35989 25697 36023
rect 25697 35989 25731 36023
rect 25731 35989 25740 36023
rect 25688 35980 25740 35989
rect 26792 35980 26844 36032
rect 29552 35980 29604 36032
rect 30748 35980 30800 36032
rect 3662 35878 3714 35930
rect 3726 35878 3778 35930
rect 3790 35878 3842 35930
rect 3854 35878 3906 35930
rect 3918 35878 3970 35930
rect 11436 35878 11488 35930
rect 11500 35878 11552 35930
rect 11564 35878 11616 35930
rect 11628 35878 11680 35930
rect 11692 35878 11744 35930
rect 19210 35878 19262 35930
rect 19274 35878 19326 35930
rect 19338 35878 19390 35930
rect 19402 35878 19454 35930
rect 19466 35878 19518 35930
rect 26984 35878 27036 35930
rect 27048 35878 27100 35930
rect 27112 35878 27164 35930
rect 27176 35878 27228 35930
rect 27240 35878 27292 35930
rect 10048 35776 10100 35828
rect 12624 35776 12676 35828
rect 12716 35819 12768 35828
rect 12716 35785 12725 35819
rect 12725 35785 12759 35819
rect 12759 35785 12768 35819
rect 12716 35776 12768 35785
rect 12808 35776 12860 35828
rect 14648 35776 14700 35828
rect 12256 35708 12308 35760
rect 8300 35640 8352 35692
rect 9496 35615 9548 35624
rect 9496 35581 9505 35615
rect 9505 35581 9539 35615
rect 9539 35581 9548 35615
rect 9496 35572 9548 35581
rect 9772 35615 9824 35624
rect 9772 35581 9781 35615
rect 9781 35581 9815 35615
rect 9815 35581 9824 35615
rect 9772 35572 9824 35581
rect 10140 35572 10192 35624
rect 12808 35640 12860 35692
rect 10508 35504 10560 35556
rect 11520 35547 11572 35556
rect 11520 35513 11554 35547
rect 11554 35513 11572 35547
rect 11520 35504 11572 35513
rect 11704 35504 11756 35556
rect 13084 35615 13136 35624
rect 13084 35581 13093 35615
rect 13093 35581 13127 35615
rect 13127 35581 13136 35615
rect 13084 35572 13136 35581
rect 13452 35640 13504 35692
rect 15016 35640 15068 35692
rect 15752 35708 15804 35760
rect 17132 35776 17184 35828
rect 21548 35776 21600 35828
rect 22560 35776 22612 35828
rect 23664 35776 23716 35828
rect 24584 35776 24636 35828
rect 26516 35776 26568 35828
rect 27160 35776 27212 35828
rect 28448 35776 28500 35828
rect 15292 35572 15344 35624
rect 15476 35615 15528 35624
rect 15476 35581 15485 35615
rect 15485 35581 15519 35615
rect 15519 35581 15528 35615
rect 15476 35572 15528 35581
rect 10324 35436 10376 35488
rect 11612 35436 11664 35488
rect 13268 35504 13320 35556
rect 13544 35547 13596 35556
rect 13544 35513 13553 35547
rect 13553 35513 13587 35547
rect 13587 35513 13596 35547
rect 13544 35504 13596 35513
rect 13728 35547 13780 35556
rect 13728 35513 13737 35547
rect 13737 35513 13771 35547
rect 13771 35513 13780 35547
rect 15660 35572 15712 35624
rect 16488 35708 16540 35760
rect 16028 35640 16080 35692
rect 13728 35504 13780 35513
rect 16212 35615 16264 35624
rect 16212 35581 16221 35615
rect 16221 35581 16255 35615
rect 16255 35581 16264 35615
rect 16212 35572 16264 35581
rect 12900 35436 12952 35488
rect 15476 35436 15528 35488
rect 16488 35615 16540 35624
rect 16488 35581 16497 35615
rect 16497 35581 16531 35615
rect 16531 35581 16540 35615
rect 16488 35572 16540 35581
rect 16764 35615 16816 35624
rect 16764 35581 16773 35615
rect 16773 35581 16807 35615
rect 16807 35581 16816 35615
rect 16764 35572 16816 35581
rect 21824 35683 21876 35692
rect 21824 35649 21833 35683
rect 21833 35649 21867 35683
rect 21867 35649 21876 35683
rect 21824 35640 21876 35649
rect 26884 35640 26936 35692
rect 18604 35572 18656 35624
rect 19800 35572 19852 35624
rect 20628 35615 20680 35624
rect 20628 35581 20662 35615
rect 20662 35581 20680 35615
rect 20628 35572 20680 35581
rect 23940 35572 23992 35624
rect 24124 35572 24176 35624
rect 26700 35572 26752 35624
rect 27988 35640 28040 35692
rect 28908 35640 28960 35692
rect 29644 35572 29696 35624
rect 20812 35504 20864 35556
rect 22192 35504 22244 35556
rect 25320 35504 25372 35556
rect 16488 35436 16540 35488
rect 18144 35479 18196 35488
rect 18144 35445 18153 35479
rect 18153 35445 18187 35479
rect 18187 35445 18196 35479
rect 18144 35436 18196 35445
rect 18788 35436 18840 35488
rect 19708 35436 19760 35488
rect 20260 35436 20312 35488
rect 27252 35436 27304 35488
rect 27988 35479 28040 35488
rect 27988 35445 27997 35479
rect 27997 35445 28031 35479
rect 28031 35445 28040 35479
rect 27988 35436 28040 35445
rect 28448 35436 28500 35488
rect 30840 35436 30892 35488
rect 4322 35334 4374 35386
rect 4386 35334 4438 35386
rect 4450 35334 4502 35386
rect 4514 35334 4566 35386
rect 4578 35334 4630 35386
rect 12096 35334 12148 35386
rect 12160 35334 12212 35386
rect 12224 35334 12276 35386
rect 12288 35334 12340 35386
rect 12352 35334 12404 35386
rect 19870 35334 19922 35386
rect 19934 35334 19986 35386
rect 19998 35334 20050 35386
rect 20062 35334 20114 35386
rect 20126 35334 20178 35386
rect 27644 35334 27696 35386
rect 27708 35334 27760 35386
rect 27772 35334 27824 35386
rect 27836 35334 27888 35386
rect 27900 35334 27952 35386
rect 10140 35232 10192 35284
rect 11520 35232 11572 35284
rect 11980 35232 12032 35284
rect 12624 35164 12676 35216
rect 10048 35096 10100 35148
rect 11612 35096 11664 35148
rect 9772 35028 9824 35080
rect 11244 35028 11296 35080
rect 11888 35139 11940 35148
rect 11888 35105 11897 35139
rect 11897 35105 11931 35139
rect 11931 35105 11940 35139
rect 11888 35096 11940 35105
rect 12072 35139 12124 35148
rect 12072 35105 12081 35139
rect 12081 35105 12115 35139
rect 12115 35105 12124 35139
rect 12072 35096 12124 35105
rect 12164 35096 12216 35148
rect 12716 35028 12768 35080
rect 15476 35232 15528 35284
rect 16212 35232 16264 35284
rect 16764 35232 16816 35284
rect 19800 35232 19852 35284
rect 22192 35275 22244 35284
rect 22192 35241 22201 35275
rect 22201 35241 22235 35275
rect 22235 35241 22244 35275
rect 22192 35232 22244 35241
rect 13360 35139 13412 35148
rect 13360 35105 13369 35139
rect 13369 35105 13403 35139
rect 13403 35105 13412 35139
rect 13360 35096 13412 35105
rect 15016 35164 15068 35216
rect 13636 35139 13688 35148
rect 13636 35105 13645 35139
rect 13645 35105 13679 35139
rect 13679 35105 13688 35139
rect 13636 35096 13688 35105
rect 13728 35139 13780 35148
rect 13728 35105 13737 35139
rect 13737 35105 13771 35139
rect 13771 35105 13780 35139
rect 13728 35096 13780 35105
rect 14280 35139 14332 35148
rect 14280 35105 14289 35139
rect 14289 35105 14323 35139
rect 14323 35105 14332 35139
rect 14280 35096 14332 35105
rect 13636 34960 13688 35012
rect 10048 34892 10100 34944
rect 11704 34892 11756 34944
rect 11888 34892 11940 34944
rect 12164 34892 12216 34944
rect 13452 34892 13504 34944
rect 13912 34892 13964 34944
rect 14556 35139 14608 35148
rect 14556 35105 14565 35139
rect 14565 35105 14599 35139
rect 14599 35105 14608 35139
rect 14556 35096 14608 35105
rect 14648 35139 14700 35148
rect 14648 35105 14657 35139
rect 14657 35105 14691 35139
rect 14691 35105 14700 35139
rect 14648 35096 14700 35105
rect 14740 35139 14792 35148
rect 14740 35105 14749 35139
rect 14749 35105 14783 35139
rect 14783 35105 14792 35139
rect 14740 35096 14792 35105
rect 15108 35096 15160 35148
rect 18696 35164 18748 35216
rect 16396 35139 16448 35148
rect 16396 35105 16405 35139
rect 16405 35105 16439 35139
rect 16439 35105 16448 35139
rect 16396 35096 16448 35105
rect 16948 35096 17000 35148
rect 18788 35139 18840 35148
rect 18788 35105 18797 35139
rect 18797 35105 18831 35139
rect 18831 35105 18840 35139
rect 18788 35096 18840 35105
rect 21916 35164 21968 35216
rect 22560 35232 22612 35284
rect 25320 35275 25372 35284
rect 25320 35241 25329 35275
rect 25329 35241 25363 35275
rect 25363 35241 25372 35275
rect 25320 35232 25372 35241
rect 26700 35207 26752 35216
rect 26700 35173 26709 35207
rect 26709 35173 26743 35207
rect 26743 35173 26752 35207
rect 26700 35164 26752 35173
rect 26884 35207 26936 35216
rect 26884 35173 26893 35207
rect 26893 35173 26927 35207
rect 26927 35173 26936 35207
rect 26884 35164 26936 35173
rect 27252 35275 27304 35284
rect 27252 35241 27277 35275
rect 27277 35241 27304 35275
rect 27252 35232 27304 35241
rect 28080 35232 28132 35284
rect 29184 35232 29236 35284
rect 30288 35232 30340 35284
rect 18052 35028 18104 35080
rect 20720 35096 20772 35148
rect 16028 34960 16080 35012
rect 17408 34960 17460 35012
rect 15292 34892 15344 34944
rect 15476 34892 15528 34944
rect 17224 34892 17276 34944
rect 18880 34960 18932 35012
rect 19708 34960 19760 35012
rect 20812 35028 20864 35080
rect 22928 35071 22980 35080
rect 22928 35037 22937 35071
rect 22937 35037 22971 35071
rect 22971 35037 22980 35071
rect 22928 35028 22980 35037
rect 23848 35028 23900 35080
rect 24860 35096 24912 35148
rect 25044 35028 25096 35080
rect 25688 35096 25740 35148
rect 28172 35139 28224 35148
rect 28172 35105 28181 35139
rect 28181 35105 28215 35139
rect 28215 35105 28224 35139
rect 28172 35096 28224 35105
rect 28356 35096 28408 35148
rect 30196 35164 30248 35216
rect 29644 35139 29696 35148
rect 27988 35028 28040 35080
rect 29644 35105 29653 35139
rect 29653 35105 29687 35139
rect 29687 35105 29696 35139
rect 29644 35096 29696 35105
rect 29736 35139 29788 35148
rect 29736 35105 29745 35139
rect 29745 35105 29779 35139
rect 29779 35105 29788 35139
rect 29736 35096 29788 35105
rect 22744 34960 22796 35012
rect 24032 34960 24084 35012
rect 19892 34892 19944 34944
rect 22100 34892 22152 34944
rect 27160 34892 27212 34944
rect 27344 34892 27396 34944
rect 28724 35003 28776 35012
rect 28724 34969 28733 35003
rect 28733 34969 28767 35003
rect 28767 34969 28776 35003
rect 28724 34960 28776 34969
rect 28908 34960 28960 35012
rect 27988 34892 28040 34944
rect 28632 34892 28684 34944
rect 29920 34960 29972 35012
rect 30564 35139 30616 35148
rect 30564 35105 30573 35139
rect 30573 35105 30607 35139
rect 30607 35105 30616 35139
rect 30564 35096 30616 35105
rect 30840 35071 30892 35080
rect 30840 35037 30849 35071
rect 30849 35037 30883 35071
rect 30883 35037 30892 35071
rect 30840 35028 30892 35037
rect 30288 34892 30340 34944
rect 3662 34790 3714 34842
rect 3726 34790 3778 34842
rect 3790 34790 3842 34842
rect 3854 34790 3906 34842
rect 3918 34790 3970 34842
rect 11436 34790 11488 34842
rect 11500 34790 11552 34842
rect 11564 34790 11616 34842
rect 11628 34790 11680 34842
rect 11692 34790 11744 34842
rect 19210 34790 19262 34842
rect 19274 34790 19326 34842
rect 19338 34790 19390 34842
rect 19402 34790 19454 34842
rect 19466 34790 19518 34842
rect 26984 34790 27036 34842
rect 27048 34790 27100 34842
rect 27112 34790 27164 34842
rect 27176 34790 27228 34842
rect 27240 34790 27292 34842
rect 9680 34688 9732 34740
rect 10416 34688 10468 34740
rect 11796 34688 11848 34740
rect 12072 34688 12124 34740
rect 14556 34688 14608 34740
rect 14740 34688 14792 34740
rect 9128 34484 9180 34536
rect 8852 34416 8904 34468
rect 10048 34527 10100 34536
rect 10048 34493 10057 34527
rect 10057 34493 10091 34527
rect 10091 34493 10100 34527
rect 10048 34484 10100 34493
rect 12440 34620 12492 34672
rect 13452 34620 13504 34672
rect 16488 34688 16540 34740
rect 11060 34484 11112 34536
rect 12808 34484 12860 34536
rect 12900 34527 12952 34536
rect 12900 34493 12909 34527
rect 12909 34493 12943 34527
rect 12943 34493 12952 34527
rect 12900 34484 12952 34493
rect 13268 34484 13320 34536
rect 13912 34527 13964 34536
rect 13912 34493 13946 34527
rect 13946 34493 13964 34527
rect 13912 34484 13964 34493
rect 13176 34416 13228 34468
rect 13728 34416 13780 34468
rect 16672 34552 16724 34604
rect 19064 34688 19116 34740
rect 20720 34731 20772 34740
rect 20720 34697 20729 34731
rect 20729 34697 20763 34731
rect 20763 34697 20772 34731
rect 20720 34688 20772 34697
rect 15108 34527 15160 34536
rect 15108 34493 15117 34527
rect 15117 34493 15151 34527
rect 15151 34493 15160 34527
rect 15108 34484 15160 34493
rect 16028 34527 16080 34536
rect 16028 34493 16037 34527
rect 16037 34493 16071 34527
rect 16071 34493 16080 34527
rect 16028 34484 16080 34493
rect 18052 34552 18104 34604
rect 18144 34552 18196 34604
rect 18972 34595 19024 34604
rect 18972 34561 18981 34595
rect 18981 34561 19015 34595
rect 19015 34561 19024 34595
rect 18972 34552 19024 34561
rect 22100 34688 22152 34740
rect 22928 34688 22980 34740
rect 23940 34731 23992 34740
rect 23940 34697 23949 34731
rect 23949 34697 23983 34731
rect 23983 34697 23992 34731
rect 23940 34688 23992 34697
rect 25688 34688 25740 34740
rect 26700 34688 26752 34740
rect 28356 34731 28408 34740
rect 28356 34697 28365 34731
rect 28365 34697 28399 34731
rect 28399 34697 28408 34731
rect 28356 34688 28408 34697
rect 29644 34688 29696 34740
rect 29736 34688 29788 34740
rect 30196 34688 30248 34740
rect 30564 34688 30616 34740
rect 22836 34620 22888 34672
rect 24952 34620 25004 34672
rect 17960 34484 18012 34536
rect 9312 34348 9364 34400
rect 10324 34348 10376 34400
rect 13912 34348 13964 34400
rect 14188 34348 14240 34400
rect 18236 34348 18288 34400
rect 19616 34484 19668 34536
rect 19892 34484 19944 34536
rect 19524 34416 19576 34468
rect 21088 34484 21140 34536
rect 22008 34484 22060 34536
rect 22376 34484 22428 34536
rect 23480 34484 23532 34536
rect 25412 34552 25464 34604
rect 26240 34552 26292 34604
rect 24768 34527 24820 34536
rect 24768 34493 24777 34527
rect 24777 34493 24811 34527
rect 24811 34493 24820 34527
rect 24768 34484 24820 34493
rect 25044 34527 25096 34536
rect 25044 34493 25053 34527
rect 25053 34493 25087 34527
rect 25087 34493 25096 34527
rect 25044 34484 25096 34493
rect 28632 34527 28684 34536
rect 28632 34493 28641 34527
rect 28641 34493 28675 34527
rect 28675 34493 28684 34527
rect 28632 34484 28684 34493
rect 31300 34527 31352 34536
rect 31300 34493 31309 34527
rect 31309 34493 31343 34527
rect 31343 34493 31352 34527
rect 31300 34484 31352 34493
rect 19800 34348 19852 34400
rect 21088 34348 21140 34400
rect 22560 34459 22612 34468
rect 22560 34425 22569 34459
rect 22569 34425 22603 34459
rect 22603 34425 22612 34459
rect 22560 34416 22612 34425
rect 24124 34459 24176 34468
rect 24124 34425 24133 34459
rect 24133 34425 24167 34459
rect 24167 34425 24176 34459
rect 24124 34416 24176 34425
rect 24492 34416 24544 34468
rect 25136 34459 25188 34468
rect 25136 34425 25145 34459
rect 25145 34425 25179 34459
rect 25179 34425 25188 34459
rect 25136 34416 25188 34425
rect 27344 34416 27396 34468
rect 29276 34459 29328 34468
rect 29276 34425 29310 34459
rect 29310 34425 29328 34459
rect 29276 34416 29328 34425
rect 22376 34391 22428 34400
rect 22376 34357 22385 34391
rect 22385 34357 22419 34391
rect 22419 34357 22428 34391
rect 22376 34348 22428 34357
rect 23572 34391 23624 34400
rect 23572 34357 23581 34391
rect 23581 34357 23615 34391
rect 23615 34357 23624 34391
rect 23572 34348 23624 34357
rect 24584 34391 24636 34400
rect 24584 34357 24593 34391
rect 24593 34357 24627 34391
rect 24627 34357 24636 34391
rect 24584 34348 24636 34357
rect 25596 34348 25648 34400
rect 4322 34246 4374 34298
rect 4386 34246 4438 34298
rect 4450 34246 4502 34298
rect 4514 34246 4566 34298
rect 4578 34246 4630 34298
rect 12096 34246 12148 34298
rect 12160 34246 12212 34298
rect 12224 34246 12276 34298
rect 12288 34246 12340 34298
rect 12352 34246 12404 34298
rect 19870 34246 19922 34298
rect 19934 34246 19986 34298
rect 19998 34246 20050 34298
rect 20062 34246 20114 34298
rect 20126 34246 20178 34298
rect 27644 34246 27696 34298
rect 27708 34246 27760 34298
rect 27772 34246 27824 34298
rect 27836 34246 27888 34298
rect 27900 34246 27952 34298
rect 8852 34187 8904 34196
rect 8852 34153 8861 34187
rect 8861 34153 8895 34187
rect 8895 34153 8904 34187
rect 8852 34144 8904 34153
rect 9496 34144 9548 34196
rect 11336 34144 11388 34196
rect 11796 34144 11848 34196
rect 12900 34144 12952 34196
rect 9220 34051 9272 34060
rect 9220 34017 9229 34051
rect 9229 34017 9263 34051
rect 9263 34017 9272 34051
rect 9220 34008 9272 34017
rect 9312 34051 9364 34060
rect 9312 34017 9321 34051
rect 9321 34017 9355 34051
rect 9355 34017 9364 34051
rect 9312 34008 9364 34017
rect 10232 34076 10284 34128
rect 12440 34076 12492 34128
rect 13544 34076 13596 34128
rect 14280 34144 14332 34196
rect 9772 34051 9824 34060
rect 9772 34017 9781 34051
rect 9781 34017 9815 34051
rect 9815 34017 9824 34051
rect 9772 34008 9824 34017
rect 11888 34008 11940 34060
rect 12992 34051 13044 34060
rect 12992 34017 13001 34051
rect 13001 34017 13035 34051
rect 13035 34017 13044 34051
rect 12992 34008 13044 34017
rect 14740 34008 14792 34060
rect 9680 33940 9732 33992
rect 13544 33940 13596 33992
rect 13912 33983 13964 33992
rect 13912 33949 13921 33983
rect 13921 33949 13955 33983
rect 13955 33949 13964 33983
rect 13912 33940 13964 33949
rect 9312 33872 9364 33924
rect 11244 33872 11296 33924
rect 12072 33872 12124 33924
rect 12716 33872 12768 33924
rect 13268 33872 13320 33924
rect 11796 33804 11848 33856
rect 12808 33804 12860 33856
rect 15476 34051 15528 34060
rect 15476 34017 15485 34051
rect 15485 34017 15519 34051
rect 15519 34017 15528 34051
rect 15476 34008 15528 34017
rect 15568 34008 15620 34060
rect 16304 34008 16356 34060
rect 16580 34051 16632 34060
rect 16580 34017 16589 34051
rect 16589 34017 16623 34051
rect 16623 34017 16632 34051
rect 16580 34008 16632 34017
rect 18144 34187 18196 34196
rect 18144 34153 18153 34187
rect 18153 34153 18187 34187
rect 18187 34153 18196 34187
rect 18144 34144 18196 34153
rect 18236 34187 18288 34196
rect 18236 34153 18245 34187
rect 18245 34153 18279 34187
rect 18279 34153 18288 34187
rect 18236 34144 18288 34153
rect 18972 34144 19024 34196
rect 22284 34144 22336 34196
rect 16764 34076 16816 34128
rect 22100 34076 22152 34128
rect 25136 34144 25188 34196
rect 29276 34144 29328 34196
rect 31300 34187 31352 34196
rect 31300 34153 31309 34187
rect 31309 34153 31343 34187
rect 31343 34153 31352 34187
rect 31300 34144 31352 34153
rect 17960 33940 18012 33992
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18512 34051 18564 34060
rect 18512 34017 18521 34051
rect 18521 34017 18555 34051
rect 18555 34017 18564 34051
rect 18512 34008 18564 34017
rect 18880 34051 18932 34060
rect 18880 34017 18889 34051
rect 18889 34017 18923 34051
rect 18923 34017 18932 34051
rect 18880 34008 18932 34017
rect 19156 34008 19208 34060
rect 19616 34008 19668 34060
rect 19708 34008 19760 34060
rect 19800 34051 19852 34060
rect 19800 34017 19809 34051
rect 19809 34017 19843 34051
rect 19843 34017 19852 34051
rect 19800 34008 19852 34017
rect 23572 34076 23624 34128
rect 26424 34076 26476 34128
rect 26792 34076 26844 34128
rect 27344 34119 27396 34128
rect 27344 34085 27353 34119
rect 27353 34085 27387 34119
rect 27387 34085 27396 34119
rect 27344 34076 27396 34085
rect 27988 34076 28040 34128
rect 22560 34008 22612 34060
rect 24584 34051 24636 34060
rect 24584 34017 24593 34051
rect 24593 34017 24627 34051
rect 24627 34017 24636 34051
rect 24584 34008 24636 34017
rect 24860 34051 24912 34060
rect 24860 34017 24894 34051
rect 24894 34017 24912 34051
rect 24860 34008 24912 34017
rect 26240 34051 26292 34060
rect 26240 34017 26249 34051
rect 26249 34017 26283 34051
rect 26283 34017 26292 34051
rect 26240 34008 26292 34017
rect 18052 33940 18104 33949
rect 16948 33872 17000 33924
rect 18880 33872 18932 33924
rect 21732 33983 21784 33992
rect 21732 33949 21741 33983
rect 21741 33949 21775 33983
rect 21775 33949 21784 33983
rect 21732 33940 21784 33949
rect 21824 33983 21876 33992
rect 21824 33949 21833 33983
rect 21833 33949 21867 33983
rect 21867 33949 21876 33983
rect 21824 33940 21876 33949
rect 25688 33940 25740 33992
rect 29184 34008 29236 34060
rect 29644 34076 29696 34128
rect 30288 34076 30340 34128
rect 29736 34051 29788 34060
rect 29736 34017 29745 34051
rect 29745 34017 29779 34051
rect 29779 34017 29788 34051
rect 29736 34008 29788 34017
rect 29920 34051 29972 34060
rect 29920 34017 29929 34051
rect 29929 34017 29963 34051
rect 29963 34017 29972 34051
rect 29920 34008 29972 34017
rect 25596 33872 25648 33924
rect 26516 33872 26568 33924
rect 29552 33983 29604 33992
rect 29552 33949 29561 33983
rect 29561 33949 29595 33983
rect 29595 33949 29604 33983
rect 29552 33940 29604 33949
rect 27988 33872 28040 33924
rect 28908 33872 28960 33924
rect 15384 33804 15436 33856
rect 16120 33804 16172 33856
rect 16856 33804 16908 33856
rect 18604 33804 18656 33856
rect 18788 33804 18840 33856
rect 19524 33804 19576 33856
rect 19616 33804 19668 33856
rect 20720 33804 20772 33856
rect 21272 33847 21324 33856
rect 21272 33813 21281 33847
rect 21281 33813 21315 33847
rect 21315 33813 21324 33847
rect 21272 33804 21324 33813
rect 22284 33804 22336 33856
rect 23112 33804 23164 33856
rect 24400 33804 24452 33856
rect 26148 33847 26200 33856
rect 26148 33813 26157 33847
rect 26157 33813 26191 33847
rect 26191 33813 26200 33847
rect 26148 33804 26200 33813
rect 26332 33804 26384 33856
rect 27528 33847 27580 33856
rect 27528 33813 27537 33847
rect 27537 33813 27571 33847
rect 27571 33813 27580 33847
rect 27528 33804 27580 33813
rect 28448 33804 28500 33856
rect 3662 33702 3714 33754
rect 3726 33702 3778 33754
rect 3790 33702 3842 33754
rect 3854 33702 3906 33754
rect 3918 33702 3970 33754
rect 11436 33702 11488 33754
rect 11500 33702 11552 33754
rect 11564 33702 11616 33754
rect 11628 33702 11680 33754
rect 11692 33702 11744 33754
rect 19210 33702 19262 33754
rect 19274 33702 19326 33754
rect 19338 33702 19390 33754
rect 19402 33702 19454 33754
rect 19466 33702 19518 33754
rect 26984 33702 27036 33754
rect 27048 33702 27100 33754
rect 27112 33702 27164 33754
rect 27176 33702 27228 33754
rect 27240 33702 27292 33754
rect 13636 33600 13688 33652
rect 17132 33600 17184 33652
rect 18880 33643 18932 33652
rect 18880 33609 18889 33643
rect 18889 33609 18923 33643
rect 18923 33609 18932 33643
rect 18880 33600 18932 33609
rect 21732 33643 21784 33652
rect 21732 33609 21741 33643
rect 21741 33609 21775 33643
rect 21775 33609 21784 33643
rect 21732 33600 21784 33609
rect 23848 33643 23900 33652
rect 23848 33609 23857 33643
rect 23857 33609 23891 33643
rect 23891 33609 23900 33643
rect 23848 33600 23900 33609
rect 10508 33532 10560 33584
rect 9864 33464 9916 33516
rect 10416 33464 10468 33516
rect 12348 33532 12400 33584
rect 12808 33532 12860 33584
rect 15568 33532 15620 33584
rect 16764 33532 16816 33584
rect 19064 33532 19116 33584
rect 22376 33532 22428 33584
rect 10232 33396 10284 33448
rect 9864 33328 9916 33380
rect 10048 33328 10100 33380
rect 10968 33439 11020 33448
rect 10968 33405 10977 33439
rect 10977 33405 11011 33439
rect 11011 33405 11020 33439
rect 10968 33396 11020 33405
rect 11336 33439 11388 33448
rect 11336 33405 11345 33439
rect 11345 33405 11379 33439
rect 11379 33405 11388 33439
rect 11336 33396 11388 33405
rect 11796 33464 11848 33516
rect 15292 33464 15344 33516
rect 12072 33396 12124 33448
rect 12348 33396 12400 33448
rect 12532 33439 12584 33448
rect 12532 33405 12541 33439
rect 12541 33405 12575 33439
rect 12575 33405 12584 33439
rect 12532 33396 12584 33405
rect 12624 33439 12676 33448
rect 12624 33405 12633 33439
rect 12633 33405 12667 33439
rect 12667 33405 12676 33439
rect 12624 33396 12676 33405
rect 14004 33439 14056 33448
rect 14004 33405 14013 33439
rect 14013 33405 14047 33439
rect 14047 33405 14056 33439
rect 14004 33396 14056 33405
rect 14188 33439 14240 33448
rect 14188 33405 14197 33439
rect 14197 33405 14231 33439
rect 14231 33405 14240 33439
rect 14188 33396 14240 33405
rect 16856 33507 16908 33516
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 18512 33464 18564 33516
rect 19616 33464 19668 33516
rect 11612 33328 11664 33380
rect 9956 33260 10008 33312
rect 10692 33260 10744 33312
rect 11060 33303 11112 33312
rect 11060 33269 11069 33303
rect 11069 33269 11103 33303
rect 11103 33269 11112 33303
rect 11060 33260 11112 33269
rect 12440 33260 12492 33312
rect 13636 33260 13688 33312
rect 16672 33396 16724 33448
rect 18052 33396 18104 33448
rect 18144 33396 18196 33448
rect 18972 33396 19024 33448
rect 17132 33371 17184 33380
rect 17132 33337 17166 33371
rect 17166 33337 17184 33371
rect 17132 33328 17184 33337
rect 19064 33371 19116 33380
rect 19064 33337 19073 33371
rect 19073 33337 19107 33371
rect 19107 33337 19116 33371
rect 19064 33328 19116 33337
rect 18144 33260 18196 33312
rect 18512 33260 18564 33312
rect 18972 33303 19024 33312
rect 18972 33269 18981 33303
rect 18981 33269 19015 33303
rect 19015 33269 19024 33303
rect 18972 33260 19024 33269
rect 21732 33396 21784 33448
rect 22376 33439 22428 33448
rect 22376 33405 22385 33439
rect 22385 33405 22419 33439
rect 22419 33405 22428 33439
rect 22376 33396 22428 33405
rect 21272 33328 21324 33380
rect 22100 33328 22152 33380
rect 23480 33439 23532 33448
rect 23480 33405 23489 33439
rect 23489 33405 23523 33439
rect 23523 33405 23532 33439
rect 23480 33396 23532 33405
rect 24768 33464 24820 33516
rect 25136 33464 25188 33516
rect 26148 33600 26200 33652
rect 27344 33643 27396 33652
rect 27344 33609 27353 33643
rect 27353 33609 27387 33643
rect 27387 33609 27396 33643
rect 27344 33600 27396 33609
rect 28356 33575 28408 33584
rect 28356 33541 28365 33575
rect 28365 33541 28399 33575
rect 28399 33541 28408 33575
rect 28356 33532 28408 33541
rect 28448 33507 28500 33516
rect 28448 33473 28457 33507
rect 28457 33473 28491 33507
rect 28491 33473 28500 33507
rect 28448 33464 28500 33473
rect 24216 33439 24268 33448
rect 24216 33405 24225 33439
rect 24225 33405 24259 33439
rect 24259 33405 24268 33439
rect 24216 33396 24268 33405
rect 24308 33439 24360 33448
rect 24308 33405 24317 33439
rect 24317 33405 24351 33439
rect 24351 33405 24360 33439
rect 24308 33396 24360 33405
rect 24400 33439 24452 33448
rect 24400 33405 24409 33439
rect 24409 33405 24443 33439
rect 24443 33405 24452 33439
rect 24400 33396 24452 33405
rect 24492 33396 24544 33448
rect 26056 33396 26108 33448
rect 28080 33439 28132 33448
rect 28080 33405 28089 33439
rect 28089 33405 28123 33439
rect 28123 33405 28132 33439
rect 29552 33464 29604 33516
rect 28080 33396 28132 33405
rect 28908 33396 28960 33448
rect 26424 33328 26476 33380
rect 20812 33260 20864 33312
rect 29092 33260 29144 33312
rect 4322 33158 4374 33210
rect 4386 33158 4438 33210
rect 4450 33158 4502 33210
rect 4514 33158 4566 33210
rect 4578 33158 4630 33210
rect 12096 33158 12148 33210
rect 12160 33158 12212 33210
rect 12224 33158 12276 33210
rect 12288 33158 12340 33210
rect 12352 33158 12404 33210
rect 19870 33158 19922 33210
rect 19934 33158 19986 33210
rect 19998 33158 20050 33210
rect 20062 33158 20114 33210
rect 20126 33158 20178 33210
rect 27644 33158 27696 33210
rect 27708 33158 27760 33210
rect 27772 33158 27824 33210
rect 27836 33158 27888 33210
rect 27900 33158 27952 33210
rect 10416 33099 10468 33108
rect 10416 33065 10425 33099
rect 10425 33065 10459 33099
rect 10459 33065 10468 33099
rect 10416 33056 10468 33065
rect 8852 32963 8904 32972
rect 8852 32929 8861 32963
rect 8861 32929 8895 32963
rect 8895 32929 8904 32963
rect 8852 32920 8904 32929
rect 9220 32963 9272 32972
rect 9220 32929 9229 32963
rect 9229 32929 9263 32963
rect 9263 32929 9272 32963
rect 9220 32920 9272 32929
rect 9588 32963 9640 32972
rect 9588 32929 9597 32963
rect 9597 32929 9631 32963
rect 9631 32929 9640 32963
rect 9588 32920 9640 32929
rect 10048 32988 10100 33040
rect 10140 32988 10192 33040
rect 9956 32963 10008 32972
rect 9956 32929 9965 32963
rect 9965 32929 9999 32963
rect 9999 32929 10008 32963
rect 9956 32920 10008 32929
rect 10876 32988 10928 33040
rect 12624 32988 12676 33040
rect 10508 32852 10560 32904
rect 10784 32920 10836 32972
rect 11336 32920 11388 32972
rect 11796 32920 11848 32972
rect 16672 33056 16724 33108
rect 16856 33056 16908 33108
rect 14188 33031 14240 33040
rect 14188 32997 14197 33031
rect 14197 32997 14231 33031
rect 14231 32997 14240 33031
rect 14188 32988 14240 32997
rect 15200 32988 15252 33040
rect 16488 32988 16540 33040
rect 16580 32988 16632 33040
rect 19064 33056 19116 33108
rect 21824 33056 21876 33108
rect 22560 33099 22612 33108
rect 22560 33065 22569 33099
rect 22569 33065 22603 33099
rect 22603 33065 22612 33099
rect 22560 33056 22612 33065
rect 24216 33099 24268 33108
rect 24216 33065 24225 33099
rect 24225 33065 24259 33099
rect 24259 33065 24268 33099
rect 24216 33056 24268 33065
rect 24860 33056 24912 33108
rect 26424 33099 26476 33108
rect 26424 33065 26433 33099
rect 26433 33065 26467 33099
rect 26467 33065 26476 33099
rect 26424 33056 26476 33065
rect 27528 33056 27580 33108
rect 29092 33099 29144 33108
rect 29092 33065 29101 33099
rect 29101 33065 29135 33099
rect 29135 33065 29144 33099
rect 29092 33056 29144 33065
rect 13452 32963 13504 32972
rect 13452 32929 13461 32963
rect 13461 32929 13495 32963
rect 13495 32929 13504 32963
rect 13452 32920 13504 32929
rect 13636 32963 13688 32972
rect 13636 32929 13645 32963
rect 13645 32929 13679 32963
rect 13679 32929 13688 32963
rect 13636 32920 13688 32929
rect 13820 32920 13872 32972
rect 14648 32920 14700 32972
rect 15384 32963 15436 32972
rect 15384 32929 15393 32963
rect 15393 32929 15427 32963
rect 15427 32929 15436 32963
rect 15384 32920 15436 32929
rect 16028 32920 16080 32972
rect 18420 32920 18472 32972
rect 21456 32920 21508 32972
rect 22008 32920 22060 32972
rect 22468 32920 22520 32972
rect 24124 32920 24176 32972
rect 12716 32852 12768 32904
rect 16304 32895 16356 32904
rect 16304 32861 16313 32895
rect 16313 32861 16347 32895
rect 16347 32861 16356 32895
rect 16304 32852 16356 32861
rect 15200 32827 15252 32836
rect 15200 32793 15209 32827
rect 15209 32793 15243 32827
rect 15243 32793 15252 32827
rect 15200 32784 15252 32793
rect 9404 32716 9456 32768
rect 10416 32716 10468 32768
rect 10508 32716 10560 32768
rect 11336 32716 11388 32768
rect 11428 32716 11480 32768
rect 12348 32716 12400 32768
rect 12532 32716 12584 32768
rect 16948 32852 17000 32904
rect 17684 32852 17736 32904
rect 19708 32895 19760 32904
rect 19708 32861 19717 32895
rect 19717 32861 19751 32895
rect 19751 32861 19760 32895
rect 19708 32852 19760 32861
rect 21180 32852 21232 32904
rect 16764 32784 16816 32836
rect 24952 32963 25004 32972
rect 24952 32929 24961 32963
rect 24961 32929 24995 32963
rect 24995 32929 25004 32963
rect 24952 32920 25004 32929
rect 26332 32988 26384 33040
rect 28908 32988 28960 33040
rect 25688 32920 25740 32972
rect 26608 32920 26660 32972
rect 26884 32920 26936 32972
rect 27436 32920 27488 32972
rect 28356 32963 28408 32972
rect 28356 32929 28365 32963
rect 28365 32929 28399 32963
rect 28399 32929 28408 32963
rect 28356 32920 28408 32929
rect 25044 32852 25096 32904
rect 25136 32895 25188 32904
rect 25136 32861 25145 32895
rect 25145 32861 25179 32895
rect 25179 32861 25188 32895
rect 25136 32852 25188 32861
rect 17040 32716 17092 32768
rect 19800 32759 19852 32768
rect 19800 32725 19809 32759
rect 19809 32725 19843 32759
rect 19843 32725 19852 32759
rect 19800 32716 19852 32725
rect 25504 32716 25556 32768
rect 27896 32852 27948 32904
rect 28448 32784 28500 32836
rect 27712 32716 27764 32768
rect 29000 32759 29052 32768
rect 29000 32725 29009 32759
rect 29009 32725 29043 32759
rect 29043 32725 29052 32759
rect 29000 32716 29052 32725
rect 3662 32614 3714 32666
rect 3726 32614 3778 32666
rect 3790 32614 3842 32666
rect 3854 32614 3906 32666
rect 3918 32614 3970 32666
rect 11436 32614 11488 32666
rect 11500 32614 11552 32666
rect 11564 32614 11616 32666
rect 11628 32614 11680 32666
rect 11692 32614 11744 32666
rect 19210 32614 19262 32666
rect 19274 32614 19326 32666
rect 19338 32614 19390 32666
rect 19402 32614 19454 32666
rect 19466 32614 19518 32666
rect 26984 32614 27036 32666
rect 27048 32614 27100 32666
rect 27112 32614 27164 32666
rect 27176 32614 27228 32666
rect 27240 32614 27292 32666
rect 8852 32512 8904 32564
rect 9864 32512 9916 32564
rect 10784 32512 10836 32564
rect 11244 32512 11296 32564
rect 13452 32512 13504 32564
rect 15384 32512 15436 32564
rect 15844 32555 15896 32564
rect 15844 32521 15853 32555
rect 15853 32521 15887 32555
rect 15887 32521 15896 32555
rect 15844 32512 15896 32521
rect 16120 32512 16172 32564
rect 9220 32444 9272 32496
rect 10140 32376 10192 32428
rect 9680 32308 9732 32360
rect 10416 32351 10468 32360
rect 10416 32317 10425 32351
rect 10425 32317 10459 32351
rect 10459 32317 10468 32351
rect 10416 32308 10468 32317
rect 10508 32351 10560 32360
rect 10508 32317 10517 32351
rect 10517 32317 10551 32351
rect 10551 32317 10560 32351
rect 10508 32308 10560 32317
rect 10692 32351 10744 32360
rect 10692 32317 10701 32351
rect 10701 32317 10735 32351
rect 10735 32317 10744 32351
rect 10692 32308 10744 32317
rect 13820 32444 13872 32496
rect 16672 32512 16724 32564
rect 17684 32555 17736 32564
rect 17684 32521 17693 32555
rect 17693 32521 17727 32555
rect 17727 32521 17736 32555
rect 17684 32512 17736 32521
rect 18880 32512 18932 32564
rect 11796 32376 11848 32428
rect 11060 32351 11112 32360
rect 11060 32317 11069 32351
rect 11069 32317 11103 32351
rect 11103 32317 11112 32351
rect 11060 32308 11112 32317
rect 11244 32351 11296 32360
rect 11244 32317 11253 32351
rect 11253 32317 11287 32351
rect 11287 32317 11296 32351
rect 11244 32308 11296 32317
rect 11336 32351 11388 32360
rect 11336 32317 11345 32351
rect 11345 32317 11379 32351
rect 11379 32317 11388 32351
rect 11336 32308 11388 32317
rect 12348 32351 12400 32360
rect 12348 32317 12357 32351
rect 12357 32317 12391 32351
rect 12391 32317 12400 32351
rect 12348 32308 12400 32317
rect 12532 32351 12584 32360
rect 12532 32317 12541 32351
rect 12541 32317 12575 32351
rect 12575 32317 12584 32351
rect 12532 32308 12584 32317
rect 16120 32419 16172 32428
rect 16120 32385 16129 32419
rect 16129 32385 16163 32419
rect 16163 32385 16172 32419
rect 16120 32376 16172 32385
rect 10048 32240 10100 32292
rect 9680 32172 9732 32224
rect 9864 32215 9916 32224
rect 9864 32181 9873 32215
rect 9873 32181 9907 32215
rect 9907 32181 9916 32215
rect 9864 32172 9916 32181
rect 9956 32172 10008 32224
rect 11244 32172 11296 32224
rect 11888 32172 11940 32224
rect 12440 32240 12492 32292
rect 12808 32308 12860 32360
rect 16028 32308 16080 32360
rect 13820 32172 13872 32224
rect 14924 32240 14976 32292
rect 16396 32419 16448 32428
rect 16396 32385 16405 32419
rect 16405 32385 16439 32419
rect 16439 32385 16448 32419
rect 16396 32376 16448 32385
rect 17316 32308 17368 32360
rect 19432 32444 19484 32496
rect 20168 32444 20220 32496
rect 17500 32308 17552 32360
rect 18972 32376 19024 32428
rect 20904 32487 20956 32496
rect 20904 32453 20913 32487
rect 20913 32453 20947 32487
rect 20947 32453 20956 32487
rect 20904 32444 20956 32453
rect 21824 32444 21876 32496
rect 22468 32555 22520 32564
rect 22468 32521 22477 32555
rect 22477 32521 22511 32555
rect 22511 32521 22520 32555
rect 22468 32512 22520 32521
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 23480 32512 23532 32564
rect 28908 32512 28960 32564
rect 16764 32240 16816 32292
rect 16948 32283 17000 32292
rect 16948 32249 16957 32283
rect 16957 32249 16991 32283
rect 16991 32249 17000 32283
rect 16948 32240 17000 32249
rect 17960 32308 18012 32360
rect 19064 32308 19116 32360
rect 20168 32351 20220 32360
rect 20168 32317 20177 32351
rect 20177 32317 20211 32351
rect 20211 32317 20220 32351
rect 20168 32308 20220 32317
rect 20260 32351 20312 32360
rect 20260 32317 20270 32351
rect 20270 32317 20304 32351
rect 20304 32317 20312 32351
rect 20260 32308 20312 32317
rect 21088 32308 21140 32360
rect 21180 32351 21232 32360
rect 21180 32317 21189 32351
rect 21189 32317 21223 32351
rect 21223 32317 21232 32351
rect 21180 32308 21232 32317
rect 21272 32351 21324 32360
rect 21272 32317 21281 32351
rect 21281 32317 21315 32351
rect 21315 32317 21324 32351
rect 21272 32308 21324 32317
rect 21732 32351 21784 32360
rect 21732 32317 21741 32351
rect 21741 32317 21775 32351
rect 21775 32317 21784 32351
rect 21732 32308 21784 32317
rect 22192 32351 22244 32360
rect 22192 32317 22201 32351
rect 22201 32317 22235 32351
rect 22235 32317 22244 32351
rect 22192 32308 22244 32317
rect 22560 32308 22612 32360
rect 24400 32444 24452 32496
rect 22836 32351 22888 32360
rect 22836 32317 22845 32351
rect 22845 32317 22879 32351
rect 22879 32317 22888 32351
rect 22836 32308 22888 32317
rect 23020 32308 23072 32360
rect 23112 32351 23164 32360
rect 23112 32317 23121 32351
rect 23121 32317 23155 32351
rect 23155 32317 23164 32351
rect 23112 32308 23164 32317
rect 23480 32308 23532 32360
rect 26240 32308 26292 32360
rect 19156 32240 19208 32292
rect 20076 32240 20128 32292
rect 20996 32240 21048 32292
rect 27344 32240 27396 32292
rect 27712 32283 27764 32292
rect 27712 32249 27746 32283
rect 27746 32249 27764 32283
rect 27712 32240 27764 32249
rect 15660 32172 15712 32224
rect 15936 32215 15988 32224
rect 15936 32181 15945 32215
rect 15945 32181 15979 32215
rect 15979 32181 15988 32215
rect 15936 32172 15988 32181
rect 17316 32215 17368 32224
rect 17316 32181 17325 32215
rect 17325 32181 17359 32215
rect 17359 32181 17368 32215
rect 17316 32172 17368 32181
rect 17408 32172 17460 32224
rect 19524 32172 19576 32224
rect 21548 32172 21600 32224
rect 21640 32215 21692 32224
rect 21640 32181 21649 32215
rect 21649 32181 21683 32215
rect 21683 32181 21692 32215
rect 21640 32172 21692 32181
rect 22376 32215 22428 32224
rect 22376 32181 22385 32215
rect 22385 32181 22419 32215
rect 22419 32181 22428 32215
rect 22376 32172 22428 32181
rect 23296 32215 23348 32224
rect 23296 32181 23305 32215
rect 23305 32181 23339 32215
rect 23339 32181 23348 32215
rect 23296 32172 23348 32181
rect 25320 32215 25372 32224
rect 25320 32181 25329 32215
rect 25329 32181 25363 32215
rect 25363 32181 25372 32215
rect 25320 32172 25372 32181
rect 29368 32172 29420 32224
rect 4322 32070 4374 32122
rect 4386 32070 4438 32122
rect 4450 32070 4502 32122
rect 4514 32070 4566 32122
rect 4578 32070 4630 32122
rect 12096 32070 12148 32122
rect 12160 32070 12212 32122
rect 12224 32070 12276 32122
rect 12288 32070 12340 32122
rect 12352 32070 12404 32122
rect 19870 32070 19922 32122
rect 19934 32070 19986 32122
rect 19998 32070 20050 32122
rect 20062 32070 20114 32122
rect 20126 32070 20178 32122
rect 27644 32070 27696 32122
rect 27708 32070 27760 32122
rect 27772 32070 27824 32122
rect 27836 32070 27888 32122
rect 27900 32070 27952 32122
rect 10968 31968 11020 32020
rect 14924 32011 14976 32020
rect 14924 31977 14933 32011
rect 14933 31977 14967 32011
rect 14967 31977 14976 32011
rect 14924 31968 14976 31977
rect 10232 31900 10284 31952
rect 10876 31900 10928 31952
rect 11336 31900 11388 31952
rect 14464 31900 14516 31952
rect 16764 31968 16816 32020
rect 17316 31968 17368 32020
rect 9128 31875 9180 31884
rect 9128 31841 9137 31875
rect 9137 31841 9171 31875
rect 9171 31841 9180 31875
rect 9128 31832 9180 31841
rect 12716 31832 12768 31884
rect 13544 31875 13596 31884
rect 13544 31841 13553 31875
rect 13553 31841 13587 31875
rect 13587 31841 13596 31875
rect 13544 31832 13596 31841
rect 13728 31832 13780 31884
rect 15200 31875 15252 31884
rect 15200 31841 15209 31875
rect 15209 31841 15243 31875
rect 15243 31841 15252 31875
rect 15200 31832 15252 31841
rect 15292 31875 15344 31884
rect 15292 31841 15301 31875
rect 15301 31841 15335 31875
rect 15335 31841 15344 31875
rect 15292 31832 15344 31841
rect 15936 31900 15988 31952
rect 16672 31943 16724 31952
rect 16672 31909 16699 31943
rect 16699 31909 16724 31943
rect 16672 31900 16724 31909
rect 15660 31832 15712 31884
rect 15752 31832 15804 31884
rect 21364 31968 21416 32020
rect 12808 31807 12860 31816
rect 12808 31773 12817 31807
rect 12817 31773 12851 31807
rect 12851 31773 12860 31807
rect 12808 31764 12860 31773
rect 12716 31696 12768 31748
rect 14556 31764 14608 31816
rect 16856 31764 16908 31816
rect 18052 31832 18104 31884
rect 18880 31832 18932 31884
rect 19156 31875 19208 31884
rect 19156 31841 19165 31875
rect 19165 31841 19199 31875
rect 19199 31841 19208 31875
rect 19156 31832 19208 31841
rect 19524 31875 19576 31884
rect 19524 31841 19533 31875
rect 19533 31841 19567 31875
rect 19567 31841 19576 31875
rect 19524 31832 19576 31841
rect 21640 31900 21692 31952
rect 21548 31875 21600 31884
rect 21548 31841 21582 31875
rect 21582 31841 21600 31875
rect 21548 31832 21600 31841
rect 23296 31900 23348 31952
rect 19432 31764 19484 31816
rect 22376 31764 22428 31816
rect 24308 31968 24360 32020
rect 28080 31968 28132 32020
rect 24492 31900 24544 31952
rect 29000 31900 29052 31952
rect 17132 31696 17184 31748
rect 24032 31696 24084 31748
rect 26332 31832 26384 31884
rect 26700 31832 26752 31884
rect 29368 31875 29420 31884
rect 29368 31841 29377 31875
rect 29377 31841 29411 31875
rect 29411 31841 29420 31875
rect 29368 31832 29420 31841
rect 26884 31696 26936 31748
rect 8852 31628 8904 31680
rect 9312 31628 9364 31680
rect 11060 31628 11112 31680
rect 12348 31628 12400 31680
rect 14464 31671 14516 31680
rect 14464 31637 14473 31671
rect 14473 31637 14507 31671
rect 14507 31637 14516 31671
rect 14464 31628 14516 31637
rect 16948 31628 17000 31680
rect 17776 31628 17828 31680
rect 22376 31628 22428 31680
rect 25136 31628 25188 31680
rect 26516 31671 26568 31680
rect 26516 31637 26525 31671
rect 26525 31637 26559 31671
rect 26559 31637 26568 31671
rect 26516 31628 26568 31637
rect 3662 31526 3714 31578
rect 3726 31526 3778 31578
rect 3790 31526 3842 31578
rect 3854 31526 3906 31578
rect 3918 31526 3970 31578
rect 11436 31526 11488 31578
rect 11500 31526 11552 31578
rect 11564 31526 11616 31578
rect 11628 31526 11680 31578
rect 11692 31526 11744 31578
rect 19210 31526 19262 31578
rect 19274 31526 19326 31578
rect 19338 31526 19390 31578
rect 19402 31526 19454 31578
rect 19466 31526 19518 31578
rect 26984 31526 27036 31578
rect 27048 31526 27100 31578
rect 27112 31526 27164 31578
rect 27176 31526 27228 31578
rect 27240 31526 27292 31578
rect 11152 31424 11204 31476
rect 12808 31424 12860 31476
rect 20260 31424 20312 31476
rect 22192 31424 22244 31476
rect 22652 31424 22704 31476
rect 24032 31424 24084 31476
rect 8944 31263 8996 31272
rect 8944 31229 8953 31263
rect 8953 31229 8987 31263
rect 8987 31229 8996 31263
rect 8944 31220 8996 31229
rect 9312 31356 9364 31408
rect 9404 31288 9456 31340
rect 9680 31263 9732 31272
rect 9680 31229 9689 31263
rect 9689 31229 9723 31263
rect 9723 31229 9732 31263
rect 9680 31220 9732 31229
rect 8668 31127 8720 31136
rect 8668 31093 8677 31127
rect 8677 31093 8711 31127
rect 8711 31093 8720 31127
rect 8668 31084 8720 31093
rect 9588 31084 9640 31136
rect 9956 31220 10008 31272
rect 11888 31356 11940 31408
rect 12348 31356 12400 31408
rect 11244 31288 11296 31340
rect 11060 31263 11112 31272
rect 11060 31229 11069 31263
rect 11069 31229 11103 31263
rect 11103 31229 11112 31263
rect 11060 31220 11112 31229
rect 11336 31220 11388 31272
rect 11888 31220 11940 31272
rect 13452 31288 13504 31340
rect 16856 31356 16908 31408
rect 18512 31356 18564 31408
rect 20996 31356 21048 31408
rect 11336 31084 11388 31136
rect 12348 31263 12400 31272
rect 12348 31229 12357 31263
rect 12357 31229 12391 31263
rect 12391 31229 12400 31263
rect 12348 31220 12400 31229
rect 12440 31220 12492 31272
rect 13820 31263 13872 31272
rect 13820 31229 13854 31263
rect 13854 31229 13872 31263
rect 12808 31152 12860 31204
rect 13820 31220 13872 31229
rect 15200 31220 15252 31272
rect 15384 31263 15436 31272
rect 15384 31229 15393 31263
rect 15393 31229 15427 31263
rect 15427 31229 15436 31263
rect 15384 31220 15436 31229
rect 14188 31152 14240 31204
rect 15844 31263 15896 31272
rect 15844 31229 15853 31263
rect 15853 31229 15887 31263
rect 15887 31229 15896 31263
rect 15844 31220 15896 31229
rect 15936 31220 15988 31272
rect 16120 31263 16172 31272
rect 16120 31229 16129 31263
rect 16129 31229 16163 31263
rect 16163 31229 16172 31263
rect 16120 31220 16172 31229
rect 21272 31288 21324 31340
rect 21824 31356 21876 31408
rect 21916 31288 21968 31340
rect 22284 31288 22336 31340
rect 23664 31356 23716 31408
rect 24124 31356 24176 31408
rect 16580 31220 16632 31272
rect 16856 31220 16908 31272
rect 17500 31220 17552 31272
rect 17040 31152 17092 31204
rect 17776 31263 17828 31272
rect 17776 31229 17785 31263
rect 17785 31229 17819 31263
rect 17819 31229 17828 31263
rect 17776 31220 17828 31229
rect 17960 31263 18012 31272
rect 17960 31229 17969 31263
rect 17969 31229 18003 31263
rect 18003 31229 18012 31263
rect 17960 31220 18012 31229
rect 13084 31084 13136 31136
rect 15752 31084 15804 31136
rect 16488 31084 16540 31136
rect 16856 31127 16908 31136
rect 16856 31093 16865 31127
rect 16865 31093 16899 31127
rect 16899 31093 16908 31127
rect 16856 31084 16908 31093
rect 18052 31152 18104 31204
rect 18696 31263 18748 31272
rect 18696 31229 18705 31263
rect 18705 31229 18739 31263
rect 18739 31229 18748 31263
rect 18696 31220 18748 31229
rect 20812 31263 20864 31272
rect 20812 31229 20821 31263
rect 20821 31229 20855 31263
rect 20855 31229 20864 31263
rect 20812 31220 20864 31229
rect 20996 31263 21048 31272
rect 20996 31229 21005 31263
rect 21005 31229 21039 31263
rect 21039 31229 21048 31263
rect 20996 31220 21048 31229
rect 21364 31263 21416 31272
rect 21364 31229 21373 31263
rect 21373 31229 21407 31263
rect 21407 31229 21416 31263
rect 21364 31220 21416 31229
rect 22376 31220 22428 31272
rect 22560 31263 22612 31272
rect 22560 31229 22569 31263
rect 22569 31229 22603 31263
rect 22603 31229 22612 31263
rect 22560 31220 22612 31229
rect 26424 31331 26476 31340
rect 26424 31297 26433 31331
rect 26433 31297 26467 31331
rect 26467 31297 26476 31331
rect 26424 31288 26476 31297
rect 23020 31263 23072 31272
rect 23020 31229 23029 31263
rect 23029 31229 23063 31263
rect 23063 31229 23072 31263
rect 23020 31220 23072 31229
rect 23480 31263 23532 31272
rect 23480 31229 23489 31263
rect 23489 31229 23523 31263
rect 23523 31229 23532 31263
rect 23480 31220 23532 31229
rect 26056 31263 26108 31272
rect 26056 31229 26065 31263
rect 26065 31229 26099 31263
rect 26099 31229 26108 31263
rect 26056 31220 26108 31229
rect 26884 31220 26936 31272
rect 18420 31084 18472 31136
rect 21824 31195 21876 31204
rect 21824 31161 21833 31195
rect 21833 31161 21867 31195
rect 21867 31161 21876 31195
rect 21824 31152 21876 31161
rect 21916 31195 21968 31204
rect 21916 31161 21951 31195
rect 21951 31161 21968 31195
rect 21916 31152 21968 31161
rect 22468 31084 22520 31136
rect 22652 31195 22704 31204
rect 22652 31161 22661 31195
rect 22661 31161 22695 31195
rect 22695 31161 22704 31195
rect 22652 31152 22704 31161
rect 23664 31152 23716 31204
rect 23112 31084 23164 31136
rect 24216 31084 24268 31136
rect 24952 31084 25004 31136
rect 26332 31084 26384 31136
rect 26700 31195 26752 31204
rect 26700 31161 26709 31195
rect 26709 31161 26743 31195
rect 26743 31161 26752 31195
rect 26700 31152 26752 31161
rect 27988 31220 28040 31272
rect 26884 31127 26936 31136
rect 26884 31093 26893 31127
rect 26893 31093 26927 31127
rect 26927 31093 26936 31127
rect 26884 31084 26936 31093
rect 26976 31127 27028 31136
rect 26976 31093 26985 31127
rect 26985 31093 27019 31127
rect 27019 31093 27028 31127
rect 26976 31084 27028 31093
rect 27528 31127 27580 31136
rect 27528 31093 27537 31127
rect 27537 31093 27571 31127
rect 27571 31093 27580 31127
rect 27528 31084 27580 31093
rect 4322 30982 4374 31034
rect 4386 30982 4438 31034
rect 4450 30982 4502 31034
rect 4514 30982 4566 31034
rect 4578 30982 4630 31034
rect 12096 30982 12148 31034
rect 12160 30982 12212 31034
rect 12224 30982 12276 31034
rect 12288 30982 12340 31034
rect 12352 30982 12404 31034
rect 19870 30982 19922 31034
rect 19934 30982 19986 31034
rect 19998 30982 20050 31034
rect 20062 30982 20114 31034
rect 20126 30982 20178 31034
rect 27644 30982 27696 31034
rect 27708 30982 27760 31034
rect 27772 30982 27824 31034
rect 27836 30982 27888 31034
rect 27900 30982 27952 31034
rect 8944 30880 8996 30932
rect 10324 30880 10376 30932
rect 11612 30880 11664 30932
rect 12716 30880 12768 30932
rect 12808 30923 12860 30932
rect 12808 30889 12817 30923
rect 12817 30889 12851 30923
rect 12851 30889 12860 30923
rect 12808 30880 12860 30889
rect 13452 30880 13504 30932
rect 15844 30923 15896 30932
rect 15844 30889 15853 30923
rect 15853 30889 15887 30923
rect 15887 30889 15896 30923
rect 15844 30880 15896 30889
rect 16304 30880 16356 30932
rect 8668 30812 8720 30864
rect 8852 30787 8904 30796
rect 8852 30753 8861 30787
rect 8861 30753 8895 30787
rect 8895 30753 8904 30787
rect 8852 30744 8904 30753
rect 10048 30744 10100 30796
rect 11888 30787 11940 30796
rect 11888 30753 11897 30787
rect 11897 30753 11931 30787
rect 11931 30753 11940 30787
rect 11888 30744 11940 30753
rect 13084 30744 13136 30796
rect 13268 30787 13320 30796
rect 13268 30753 13277 30787
rect 13277 30753 13311 30787
rect 13311 30753 13320 30787
rect 13268 30744 13320 30753
rect 14464 30812 14516 30864
rect 15292 30812 15344 30864
rect 17868 30880 17920 30932
rect 18144 30880 18196 30932
rect 18696 30880 18748 30932
rect 23664 30923 23716 30932
rect 23664 30889 23673 30923
rect 23673 30889 23707 30923
rect 23707 30889 23716 30923
rect 23664 30880 23716 30889
rect 26056 30880 26108 30932
rect 26332 30880 26384 30932
rect 16580 30812 16632 30864
rect 26884 30880 26936 30932
rect 26976 30880 27028 30932
rect 14556 30787 14608 30796
rect 14556 30753 14565 30787
rect 14565 30753 14599 30787
rect 14599 30753 14608 30787
rect 14556 30744 14608 30753
rect 10324 30676 10376 30728
rect 11612 30719 11664 30728
rect 11612 30685 11621 30719
rect 11621 30685 11655 30719
rect 11655 30685 11664 30719
rect 11612 30676 11664 30685
rect 12072 30676 12124 30728
rect 12164 30719 12216 30728
rect 12164 30685 12173 30719
rect 12173 30685 12207 30719
rect 12207 30685 12216 30719
rect 12164 30676 12216 30685
rect 12716 30608 12768 30660
rect 14188 30608 14240 30660
rect 15568 30787 15620 30796
rect 15568 30753 15577 30787
rect 15577 30753 15611 30787
rect 15611 30753 15620 30787
rect 15568 30744 15620 30753
rect 16488 30787 16540 30796
rect 16488 30753 16497 30787
rect 16497 30753 16531 30787
rect 16531 30753 16540 30787
rect 16488 30744 16540 30753
rect 16856 30744 16908 30796
rect 17132 30719 17184 30728
rect 17132 30685 17141 30719
rect 17141 30685 17175 30719
rect 17175 30685 17184 30719
rect 17132 30676 17184 30685
rect 16304 30608 16356 30660
rect 18512 30744 18564 30796
rect 19064 30744 19116 30796
rect 22008 30744 22060 30796
rect 22376 30744 22428 30796
rect 27436 30812 27488 30864
rect 28448 30812 28500 30864
rect 11888 30540 11940 30592
rect 12532 30540 12584 30592
rect 16396 30540 16448 30592
rect 16672 30583 16724 30592
rect 16672 30549 16681 30583
rect 16681 30549 16715 30583
rect 16715 30549 16724 30583
rect 16672 30540 16724 30549
rect 23940 30787 23992 30796
rect 23940 30753 23949 30787
rect 23949 30753 23983 30787
rect 23983 30753 23992 30787
rect 23940 30744 23992 30753
rect 24216 30787 24268 30796
rect 24216 30753 24225 30787
rect 24225 30753 24259 30787
rect 24259 30753 24268 30787
rect 24216 30744 24268 30753
rect 26424 30787 26476 30796
rect 26424 30753 26433 30787
rect 26433 30753 26467 30787
rect 26467 30753 26476 30787
rect 26424 30744 26476 30753
rect 26516 30787 26568 30796
rect 26516 30753 26526 30787
rect 26526 30753 26560 30787
rect 26560 30753 26568 30787
rect 26516 30744 26568 30753
rect 27528 30744 27580 30796
rect 27988 30744 28040 30796
rect 28908 30744 28960 30796
rect 25228 30540 25280 30592
rect 25596 30583 25648 30592
rect 25596 30549 25605 30583
rect 25605 30549 25639 30583
rect 25639 30549 25648 30583
rect 25596 30540 25648 30549
rect 26700 30540 26752 30592
rect 27988 30540 28040 30592
rect 3662 30438 3714 30490
rect 3726 30438 3778 30490
rect 3790 30438 3842 30490
rect 3854 30438 3906 30490
rect 3918 30438 3970 30490
rect 11436 30438 11488 30490
rect 11500 30438 11552 30490
rect 11564 30438 11616 30490
rect 11628 30438 11680 30490
rect 11692 30438 11744 30490
rect 19210 30438 19262 30490
rect 19274 30438 19326 30490
rect 19338 30438 19390 30490
rect 19402 30438 19454 30490
rect 19466 30438 19518 30490
rect 26984 30438 27036 30490
rect 27048 30438 27100 30490
rect 27112 30438 27164 30490
rect 27176 30438 27228 30490
rect 27240 30438 27292 30490
rect 9680 30336 9732 30388
rect 12072 30336 12124 30388
rect 15568 30379 15620 30388
rect 15568 30345 15577 30379
rect 15577 30345 15611 30379
rect 15611 30345 15620 30379
rect 15568 30336 15620 30345
rect 12532 30268 12584 30320
rect 16212 30311 16264 30320
rect 16212 30277 16221 30311
rect 16221 30277 16255 30311
rect 16255 30277 16264 30311
rect 16212 30268 16264 30277
rect 15384 30200 15436 30252
rect 16672 30379 16724 30388
rect 16672 30345 16681 30379
rect 16681 30345 16715 30379
rect 16715 30345 16724 30379
rect 16672 30336 16724 30345
rect 23020 30336 23072 30388
rect 16488 30268 16540 30320
rect 17040 30311 17092 30320
rect 17040 30277 17049 30311
rect 17049 30277 17083 30311
rect 17083 30277 17092 30311
rect 17040 30268 17092 30277
rect 23940 30336 23992 30388
rect 24124 30336 24176 30388
rect 24860 30336 24912 30388
rect 9036 30175 9088 30184
rect 9036 30141 9045 30175
rect 9045 30141 9079 30175
rect 9079 30141 9088 30175
rect 9036 30132 9088 30141
rect 9404 30064 9456 30116
rect 11336 30175 11388 30184
rect 11336 30141 11370 30175
rect 11370 30141 11388 30175
rect 11336 30132 11388 30141
rect 14280 30132 14332 30184
rect 9588 30107 9640 30116
rect 9588 30073 9622 30107
rect 9622 30073 9640 30107
rect 16212 30132 16264 30184
rect 16396 30132 16448 30184
rect 16580 30132 16632 30184
rect 16672 30132 16724 30184
rect 9588 30064 9640 30073
rect 16856 30064 16908 30116
rect 14096 29996 14148 30048
rect 16120 29996 16172 30048
rect 16304 29996 16356 30048
rect 17224 30175 17276 30184
rect 17224 30141 17233 30175
rect 17233 30141 17267 30175
rect 17267 30141 17276 30175
rect 17224 30132 17276 30141
rect 23204 30200 23256 30252
rect 23848 30200 23900 30252
rect 25228 30311 25280 30320
rect 25228 30277 25237 30311
rect 25237 30277 25271 30311
rect 25271 30277 25280 30311
rect 25228 30268 25280 30277
rect 17592 30175 17644 30184
rect 17592 30141 17601 30175
rect 17601 30141 17635 30175
rect 17635 30141 17644 30175
rect 17592 30132 17644 30141
rect 17868 30175 17920 30184
rect 17868 30141 17877 30175
rect 17877 30141 17911 30175
rect 17911 30141 17920 30175
rect 17868 30132 17920 30141
rect 19064 30132 19116 30184
rect 22008 30132 22060 30184
rect 23940 30132 23992 30184
rect 24860 30175 24912 30184
rect 24860 30141 24869 30175
rect 24869 30141 24903 30175
rect 24903 30141 24912 30175
rect 24860 30132 24912 30141
rect 18512 30064 18564 30116
rect 18972 29996 19024 30048
rect 24216 30107 24268 30116
rect 24216 30073 24225 30107
rect 24225 30073 24259 30107
rect 24259 30073 24268 30107
rect 24216 30064 24268 30073
rect 24308 30107 24360 30116
rect 24308 30073 24343 30107
rect 24343 30073 24360 30107
rect 24308 30064 24360 30073
rect 24952 30107 25004 30116
rect 24952 30073 24961 30107
rect 24961 30073 24995 30107
rect 24995 30073 25004 30107
rect 24952 30064 25004 30073
rect 27344 30064 27396 30116
rect 27528 30064 27580 30116
rect 25596 29996 25648 30048
rect 28908 29996 28960 30048
rect 4322 29894 4374 29946
rect 4386 29894 4438 29946
rect 4450 29894 4502 29946
rect 4514 29894 4566 29946
rect 4578 29894 4630 29946
rect 12096 29894 12148 29946
rect 12160 29894 12212 29946
rect 12224 29894 12276 29946
rect 12288 29894 12340 29946
rect 12352 29894 12404 29946
rect 19870 29894 19922 29946
rect 19934 29894 19986 29946
rect 19998 29894 20050 29946
rect 20062 29894 20114 29946
rect 20126 29894 20178 29946
rect 27644 29894 27696 29946
rect 27708 29894 27760 29946
rect 27772 29894 27824 29946
rect 27836 29894 27888 29946
rect 27900 29894 27952 29946
rect 16764 29835 16816 29844
rect 16764 29801 16773 29835
rect 16773 29801 16807 29835
rect 16807 29801 16816 29835
rect 16764 29792 16816 29801
rect 17592 29835 17644 29844
rect 17592 29801 17601 29835
rect 17601 29801 17635 29835
rect 17635 29801 17644 29835
rect 17592 29792 17644 29801
rect 11888 29724 11940 29776
rect 14648 29724 14700 29776
rect 16672 29724 16724 29776
rect 17408 29767 17460 29776
rect 17408 29733 17433 29767
rect 17433 29733 17460 29767
rect 17408 29724 17460 29733
rect 18144 29724 18196 29776
rect 19616 29792 19668 29844
rect 21732 29792 21784 29844
rect 24308 29792 24360 29844
rect 26516 29792 26568 29844
rect 26792 29792 26844 29844
rect 27620 29835 27672 29844
rect 27620 29801 27629 29835
rect 27629 29801 27663 29835
rect 27663 29801 27672 29835
rect 27620 29792 27672 29801
rect 28080 29792 28132 29844
rect 14096 29699 14148 29708
rect 14096 29665 14105 29699
rect 14105 29665 14139 29699
rect 14139 29665 14148 29699
rect 14096 29656 14148 29665
rect 14740 29656 14792 29708
rect 15936 29656 15988 29708
rect 16488 29656 16540 29708
rect 17316 29656 17368 29708
rect 17040 29588 17092 29640
rect 17224 29588 17276 29640
rect 17960 29699 18012 29708
rect 17960 29665 17969 29699
rect 17969 29665 18003 29699
rect 18003 29665 18012 29699
rect 19892 29724 19944 29776
rect 17960 29656 18012 29665
rect 18972 29699 19024 29708
rect 18972 29665 18981 29699
rect 18981 29665 19015 29699
rect 19015 29665 19024 29699
rect 18972 29656 19024 29665
rect 19616 29656 19668 29708
rect 20260 29724 20312 29776
rect 20444 29656 20496 29708
rect 21732 29699 21784 29708
rect 21732 29665 21741 29699
rect 21741 29665 21775 29699
rect 21775 29665 21784 29699
rect 21732 29656 21784 29665
rect 21824 29699 21876 29708
rect 21824 29665 21833 29699
rect 21833 29665 21867 29699
rect 21867 29665 21876 29699
rect 21824 29656 21876 29665
rect 22008 29699 22060 29708
rect 22008 29665 22017 29699
rect 22017 29665 22051 29699
rect 22051 29665 22060 29699
rect 22008 29656 22060 29665
rect 22284 29699 22336 29708
rect 22284 29665 22293 29699
rect 22293 29665 22327 29699
rect 22327 29665 22336 29699
rect 22284 29656 22336 29665
rect 22376 29699 22428 29708
rect 22376 29665 22385 29699
rect 22385 29665 22419 29699
rect 22419 29665 22428 29699
rect 22376 29656 22428 29665
rect 23480 29724 23532 29776
rect 23572 29699 23624 29708
rect 23572 29665 23581 29699
rect 23581 29665 23615 29699
rect 23615 29665 23624 29699
rect 23572 29656 23624 29665
rect 26608 29724 26660 29776
rect 25228 29699 25280 29708
rect 25228 29665 25237 29699
rect 25237 29665 25271 29699
rect 25271 29665 25280 29699
rect 25228 29656 25280 29665
rect 20812 29588 20864 29640
rect 21180 29520 21232 29572
rect 25136 29588 25188 29640
rect 26700 29699 26752 29708
rect 26700 29665 26709 29699
rect 26709 29665 26743 29699
rect 26743 29665 26752 29699
rect 26700 29656 26752 29665
rect 28448 29699 28500 29708
rect 28448 29665 28457 29699
rect 28457 29665 28491 29699
rect 28491 29665 28500 29699
rect 28448 29656 28500 29665
rect 26608 29631 26660 29640
rect 26608 29597 26617 29631
rect 26617 29597 26651 29631
rect 26651 29597 26660 29631
rect 26608 29588 26660 29597
rect 26792 29631 26844 29640
rect 26792 29597 26801 29631
rect 26801 29597 26835 29631
rect 26835 29597 26844 29631
rect 26792 29588 26844 29597
rect 27436 29588 27488 29640
rect 28908 29588 28960 29640
rect 23112 29520 23164 29572
rect 25780 29520 25832 29572
rect 28172 29563 28224 29572
rect 28172 29529 28181 29563
rect 28181 29529 28215 29563
rect 28215 29529 28224 29563
rect 28172 29520 28224 29529
rect 16120 29495 16172 29504
rect 16120 29461 16129 29495
rect 16129 29461 16163 29495
rect 16163 29461 16172 29495
rect 16120 29452 16172 29461
rect 16488 29495 16540 29504
rect 16488 29461 16497 29495
rect 16497 29461 16531 29495
rect 16531 29461 16540 29495
rect 16488 29452 16540 29461
rect 16580 29452 16632 29504
rect 18052 29452 18104 29504
rect 20352 29452 20404 29504
rect 20444 29452 20496 29504
rect 22192 29452 22244 29504
rect 22652 29495 22704 29504
rect 22652 29461 22661 29495
rect 22661 29461 22695 29495
rect 22695 29461 22704 29495
rect 22652 29452 22704 29461
rect 23204 29452 23256 29504
rect 27988 29452 28040 29504
rect 3662 29350 3714 29402
rect 3726 29350 3778 29402
rect 3790 29350 3842 29402
rect 3854 29350 3906 29402
rect 3918 29350 3970 29402
rect 11436 29350 11488 29402
rect 11500 29350 11552 29402
rect 11564 29350 11616 29402
rect 11628 29350 11680 29402
rect 11692 29350 11744 29402
rect 19210 29350 19262 29402
rect 19274 29350 19326 29402
rect 19338 29350 19390 29402
rect 19402 29350 19454 29402
rect 19466 29350 19518 29402
rect 26984 29350 27036 29402
rect 27048 29350 27100 29402
rect 27112 29350 27164 29402
rect 27176 29350 27228 29402
rect 27240 29350 27292 29402
rect 11520 29248 11572 29300
rect 11888 29248 11940 29300
rect 13084 29248 13136 29300
rect 14372 29248 14424 29300
rect 14740 29291 14792 29300
rect 14740 29257 14749 29291
rect 14749 29257 14783 29291
rect 14783 29257 14792 29291
rect 14740 29248 14792 29257
rect 16672 29248 16724 29300
rect 17960 29248 18012 29300
rect 18144 29291 18196 29300
rect 18144 29257 18153 29291
rect 18153 29257 18187 29291
rect 18187 29257 18196 29291
rect 18144 29248 18196 29257
rect 19616 29291 19668 29300
rect 19616 29257 19625 29291
rect 19625 29257 19659 29291
rect 19659 29257 19668 29291
rect 19616 29248 19668 29257
rect 25596 29248 25648 29300
rect 11336 29180 11388 29232
rect 11704 29180 11756 29232
rect 9404 29044 9456 29096
rect 11520 29044 11572 29096
rect 11704 29087 11756 29096
rect 11704 29053 11713 29087
rect 11713 29053 11747 29087
rect 11747 29053 11756 29087
rect 11704 29044 11756 29053
rect 12440 29044 12492 29096
rect 11980 28976 12032 29028
rect 11060 28908 11112 28960
rect 12440 28951 12492 28960
rect 12440 28917 12449 28951
rect 12449 28917 12483 28951
rect 12483 28917 12492 28951
rect 12440 28908 12492 28917
rect 12624 28951 12676 28960
rect 12624 28917 12633 28951
rect 12633 28917 12667 28951
rect 12667 28917 12676 28951
rect 12624 28908 12676 28917
rect 13084 29087 13136 29096
rect 13084 29053 13093 29087
rect 13093 29053 13127 29087
rect 13127 29053 13136 29087
rect 13084 29044 13136 29053
rect 13176 29087 13228 29096
rect 13176 29053 13185 29087
rect 13185 29053 13219 29087
rect 13219 29053 13228 29087
rect 13176 29044 13228 29053
rect 14188 29087 14240 29096
rect 14188 29053 14197 29087
rect 14197 29053 14231 29087
rect 14231 29053 14240 29087
rect 14188 29044 14240 29053
rect 14372 29044 14424 29096
rect 15292 29180 15344 29232
rect 16212 29180 16264 29232
rect 16120 29112 16172 29164
rect 15660 29044 15712 29096
rect 18512 29112 18564 29164
rect 19432 29044 19484 29096
rect 19892 29180 19944 29232
rect 26884 29180 26936 29232
rect 20352 29112 20404 29164
rect 20444 29155 20496 29164
rect 20444 29121 20453 29155
rect 20453 29121 20487 29155
rect 20487 29121 20496 29155
rect 20444 29112 20496 29121
rect 23664 29155 23716 29164
rect 23664 29121 23673 29155
rect 23673 29121 23707 29155
rect 23707 29121 23716 29155
rect 23664 29112 23716 29121
rect 25780 29155 25832 29164
rect 25780 29121 25789 29155
rect 25789 29121 25823 29155
rect 25823 29121 25832 29155
rect 25780 29112 25832 29121
rect 28356 29112 28408 29164
rect 16672 28976 16724 29028
rect 18420 28976 18472 29028
rect 19800 29019 19852 29028
rect 19800 28985 19809 29019
rect 19809 28985 19843 29019
rect 19843 28985 19852 29019
rect 19800 28976 19852 28985
rect 22652 29044 22704 29096
rect 23388 29044 23440 29096
rect 24032 29087 24084 29096
rect 24032 29053 24041 29087
rect 24041 29053 24075 29087
rect 24075 29053 24084 29087
rect 24032 29044 24084 29053
rect 25136 29087 25188 29096
rect 25136 29053 25145 29087
rect 25145 29053 25179 29087
rect 25179 29053 25188 29087
rect 25136 29044 25188 29053
rect 25228 29087 25280 29096
rect 25228 29053 25238 29087
rect 25238 29053 25272 29087
rect 25272 29053 25280 29087
rect 25228 29044 25280 29053
rect 20444 28976 20496 29028
rect 20536 28976 20588 29028
rect 22192 29019 22244 29028
rect 19340 28908 19392 28960
rect 22192 28985 22226 29019
rect 22226 28985 22244 29019
rect 22192 28976 22244 28985
rect 23204 28976 23256 29028
rect 25872 29087 25924 29096
rect 25872 29053 25881 29087
rect 25881 29053 25915 29087
rect 25915 29053 25924 29087
rect 25872 29044 25924 29053
rect 25964 29044 26016 29096
rect 27344 29044 27396 29096
rect 28172 29019 28224 29028
rect 28172 28985 28181 29019
rect 28181 28985 28215 29019
rect 28215 28985 28224 29019
rect 28172 28976 28224 28985
rect 29092 28976 29144 29028
rect 21732 28908 21784 28960
rect 21916 28908 21968 28960
rect 22468 28908 22520 28960
rect 23296 28951 23348 28960
rect 23296 28917 23305 28951
rect 23305 28917 23339 28951
rect 23339 28917 23348 28951
rect 23296 28908 23348 28917
rect 28080 28908 28132 28960
rect 4322 28806 4374 28858
rect 4386 28806 4438 28858
rect 4450 28806 4502 28858
rect 4514 28806 4566 28858
rect 4578 28806 4630 28858
rect 12096 28806 12148 28858
rect 12160 28806 12212 28858
rect 12224 28806 12276 28858
rect 12288 28806 12340 28858
rect 12352 28806 12404 28858
rect 19870 28806 19922 28858
rect 19934 28806 19986 28858
rect 19998 28806 20050 28858
rect 20062 28806 20114 28858
rect 20126 28806 20178 28858
rect 27644 28806 27696 28858
rect 27708 28806 27760 28858
rect 27772 28806 27824 28858
rect 27836 28806 27888 28858
rect 27900 28806 27952 28858
rect 11980 28704 12032 28756
rect 14280 28747 14332 28756
rect 14280 28713 14289 28747
rect 14289 28713 14323 28747
rect 14323 28713 14332 28747
rect 14280 28704 14332 28713
rect 14832 28704 14884 28756
rect 14188 28679 14240 28688
rect 14188 28645 14197 28679
rect 14197 28645 14231 28679
rect 14231 28645 14240 28679
rect 14188 28636 14240 28645
rect 11060 28568 11112 28620
rect 11244 28611 11296 28620
rect 11244 28577 11278 28611
rect 11278 28577 11296 28611
rect 11244 28568 11296 28577
rect 12440 28568 12492 28620
rect 12624 28568 12676 28620
rect 16304 28704 16356 28756
rect 17408 28747 17460 28756
rect 17408 28713 17417 28747
rect 17417 28713 17451 28747
rect 17451 28713 17460 28747
rect 17408 28704 17460 28713
rect 20536 28747 20588 28756
rect 20536 28713 20545 28747
rect 20545 28713 20579 28747
rect 20579 28713 20588 28747
rect 20536 28704 20588 28713
rect 20904 28704 20956 28756
rect 15108 28679 15160 28688
rect 15108 28645 15117 28679
rect 15117 28645 15151 28679
rect 15151 28645 15160 28679
rect 15108 28636 15160 28645
rect 13176 28500 13228 28552
rect 14464 28543 14516 28552
rect 14464 28509 14473 28543
rect 14473 28509 14507 28543
rect 14507 28509 14516 28543
rect 14464 28500 14516 28509
rect 14556 28543 14608 28552
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 14740 28543 14792 28552
rect 14740 28509 14749 28543
rect 14749 28509 14783 28543
rect 14783 28509 14792 28543
rect 14740 28500 14792 28509
rect 16304 28568 16356 28620
rect 16856 28568 16908 28620
rect 18512 28636 18564 28688
rect 21640 28679 21692 28688
rect 21640 28645 21649 28679
rect 21649 28645 21683 28679
rect 21683 28645 21692 28679
rect 21640 28636 21692 28645
rect 21916 28704 21968 28756
rect 22284 28704 22336 28756
rect 26792 28704 26844 28756
rect 15936 28500 15988 28552
rect 17868 28611 17920 28620
rect 17868 28577 17877 28611
rect 17877 28577 17911 28611
rect 17911 28577 17920 28611
rect 17868 28568 17920 28577
rect 18420 28500 18472 28552
rect 16212 28432 16264 28484
rect 19340 28568 19392 28620
rect 20260 28568 20312 28620
rect 21456 28611 21508 28620
rect 21456 28577 21465 28611
rect 21465 28577 21499 28611
rect 21499 28577 21508 28611
rect 21456 28568 21508 28577
rect 20536 28500 20588 28552
rect 21180 28500 21232 28552
rect 16672 28364 16724 28416
rect 17960 28407 18012 28416
rect 17960 28373 17969 28407
rect 17969 28373 18003 28407
rect 18003 28373 18012 28407
rect 17960 28364 18012 28373
rect 19984 28407 20036 28416
rect 19984 28373 19993 28407
rect 19993 28373 20027 28407
rect 20027 28373 20036 28407
rect 19984 28364 20036 28373
rect 21916 28611 21968 28620
rect 21916 28577 21925 28611
rect 21925 28577 21959 28611
rect 21959 28577 21968 28611
rect 21916 28568 21968 28577
rect 23204 28636 23256 28688
rect 23388 28679 23440 28688
rect 23388 28645 23422 28679
rect 23422 28645 23440 28679
rect 23388 28636 23440 28645
rect 25596 28679 25648 28688
rect 25596 28645 25605 28679
rect 25605 28645 25639 28679
rect 25639 28645 25648 28679
rect 25596 28636 25648 28645
rect 22008 28500 22060 28552
rect 21640 28432 21692 28484
rect 22468 28611 22520 28620
rect 22468 28577 22477 28611
rect 22477 28577 22511 28611
rect 22511 28577 22520 28611
rect 22468 28568 22520 28577
rect 22560 28611 22612 28620
rect 22560 28577 22569 28611
rect 22569 28577 22603 28611
rect 22603 28577 22612 28611
rect 22560 28568 22612 28577
rect 23112 28611 23164 28620
rect 23112 28577 23121 28611
rect 23121 28577 23155 28611
rect 23155 28577 23164 28611
rect 23112 28568 23164 28577
rect 21732 28364 21784 28416
rect 24584 28568 24636 28620
rect 26884 28611 26936 28620
rect 26884 28577 26893 28611
rect 26893 28577 26927 28611
rect 26927 28577 26936 28611
rect 26884 28568 26936 28577
rect 28264 28568 28316 28620
rect 29092 28611 29144 28620
rect 29092 28577 29101 28611
rect 29101 28577 29135 28611
rect 29135 28577 29144 28611
rect 29092 28568 29144 28577
rect 27344 28500 27396 28552
rect 25964 28432 26016 28484
rect 24952 28364 25004 28416
rect 26792 28407 26844 28416
rect 26792 28373 26801 28407
rect 26801 28373 26835 28407
rect 26835 28373 26844 28407
rect 26792 28364 26844 28373
rect 28080 28364 28132 28416
rect 28448 28364 28500 28416
rect 3662 28262 3714 28314
rect 3726 28262 3778 28314
rect 3790 28262 3842 28314
rect 3854 28262 3906 28314
rect 3918 28262 3970 28314
rect 11436 28262 11488 28314
rect 11500 28262 11552 28314
rect 11564 28262 11616 28314
rect 11628 28262 11680 28314
rect 11692 28262 11744 28314
rect 19210 28262 19262 28314
rect 19274 28262 19326 28314
rect 19338 28262 19390 28314
rect 19402 28262 19454 28314
rect 19466 28262 19518 28314
rect 26984 28262 27036 28314
rect 27048 28262 27100 28314
rect 27112 28262 27164 28314
rect 27176 28262 27228 28314
rect 27240 28262 27292 28314
rect 11244 28160 11296 28212
rect 14556 28160 14608 28212
rect 16396 28160 16448 28212
rect 17500 28203 17552 28212
rect 15936 28135 15988 28144
rect 15936 28101 15945 28135
rect 15945 28101 15979 28135
rect 15979 28101 15988 28135
rect 15936 28092 15988 28101
rect 16120 28092 16172 28144
rect 17500 28169 17509 28203
rect 17509 28169 17543 28203
rect 17543 28169 17552 28203
rect 17500 28160 17552 28169
rect 18144 28160 18196 28212
rect 22100 28160 22152 28212
rect 24032 28160 24084 28212
rect 11336 27999 11388 28008
rect 11336 27965 11345 27999
rect 11345 27965 11379 27999
rect 11379 27965 11388 27999
rect 11336 27956 11388 27965
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 11796 27956 11848 28008
rect 13268 27956 13320 28008
rect 15108 27956 15160 28008
rect 16764 28024 16816 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 16120 27999 16172 28008
rect 16120 27965 16129 27999
rect 16129 27965 16163 27999
rect 16163 27965 16172 27999
rect 16120 27956 16172 27965
rect 11980 27888 12032 27940
rect 13820 27931 13872 27940
rect 13820 27897 13829 27931
rect 13829 27897 13863 27931
rect 13863 27897 13872 27931
rect 13820 27888 13872 27897
rect 15384 27888 15436 27940
rect 16304 27999 16356 28008
rect 16304 27965 16313 27999
rect 16313 27965 16347 27999
rect 16347 27965 16356 27999
rect 16304 27956 16356 27965
rect 16672 27888 16724 27940
rect 17316 27931 17368 27940
rect 17316 27897 17325 27931
rect 17325 27897 17359 27931
rect 17359 27897 17368 27931
rect 17316 27888 17368 27897
rect 16304 27820 16356 27872
rect 18420 28092 18472 28144
rect 21456 28092 21508 28144
rect 22376 28092 22428 28144
rect 22560 28092 22612 28144
rect 24952 28160 25004 28212
rect 25872 28160 25924 28212
rect 19984 28024 20036 28076
rect 20444 28024 20496 28076
rect 21732 28024 21784 28076
rect 19064 27956 19116 28008
rect 20904 27999 20956 28008
rect 20904 27965 20913 27999
rect 20913 27965 20947 27999
rect 20947 27965 20956 27999
rect 20904 27956 20956 27965
rect 22284 27999 22336 28008
rect 22284 27965 22293 27999
rect 22293 27965 22327 27999
rect 22327 27965 22336 27999
rect 22284 27956 22336 27965
rect 23756 27956 23808 28008
rect 23940 27956 23992 28008
rect 24860 28092 24912 28144
rect 28264 28203 28316 28212
rect 28264 28169 28273 28203
rect 28273 28169 28307 28203
rect 28307 28169 28316 28203
rect 28264 28160 28316 28169
rect 28356 28092 28408 28144
rect 24216 27999 24268 28008
rect 24216 27965 24225 27999
rect 24225 27965 24259 27999
rect 24259 27965 24268 27999
rect 24216 27956 24268 27965
rect 24492 27999 24544 28008
rect 24492 27965 24501 27999
rect 24501 27965 24535 27999
rect 24535 27965 24544 27999
rect 24492 27956 24544 27965
rect 25504 27956 25556 28008
rect 25780 27999 25832 28008
rect 25780 27965 25793 27999
rect 25793 27965 25832 27999
rect 22836 27888 22888 27940
rect 24308 27931 24360 27940
rect 24308 27897 24343 27931
rect 24343 27897 24360 27931
rect 24308 27888 24360 27897
rect 18696 27820 18748 27872
rect 22192 27863 22244 27872
rect 22192 27829 22201 27863
rect 22201 27829 22235 27863
rect 22235 27829 22244 27863
rect 22192 27820 22244 27829
rect 23940 27820 23992 27872
rect 24676 27888 24728 27940
rect 25780 27956 25832 27965
rect 27620 27956 27672 28008
rect 26056 27888 26108 27940
rect 27988 27888 28040 27940
rect 28264 27888 28316 27940
rect 25136 27820 25188 27872
rect 4322 27718 4374 27770
rect 4386 27718 4438 27770
rect 4450 27718 4502 27770
rect 4514 27718 4566 27770
rect 4578 27718 4630 27770
rect 12096 27718 12148 27770
rect 12160 27718 12212 27770
rect 12224 27718 12276 27770
rect 12288 27718 12340 27770
rect 12352 27718 12404 27770
rect 19870 27718 19922 27770
rect 19934 27718 19986 27770
rect 19998 27718 20050 27770
rect 20062 27718 20114 27770
rect 20126 27718 20178 27770
rect 27644 27718 27696 27770
rect 27708 27718 27760 27770
rect 27772 27718 27824 27770
rect 27836 27718 27888 27770
rect 27900 27718 27952 27770
rect 14464 27616 14516 27668
rect 16304 27616 16356 27668
rect 18144 27616 18196 27668
rect 23296 27616 23348 27668
rect 11796 27480 11848 27532
rect 12532 27480 12584 27532
rect 13268 27480 13320 27532
rect 13728 27523 13780 27532
rect 13728 27489 13737 27523
rect 13737 27489 13771 27523
rect 13771 27489 13780 27523
rect 13728 27480 13780 27489
rect 14004 27523 14056 27532
rect 14004 27489 14013 27523
rect 14013 27489 14047 27523
rect 14047 27489 14056 27523
rect 14004 27480 14056 27489
rect 15108 27548 15160 27600
rect 16764 27591 16816 27600
rect 16764 27557 16773 27591
rect 16773 27557 16807 27591
rect 16807 27557 16816 27591
rect 16764 27548 16816 27557
rect 18236 27591 18288 27600
rect 18236 27557 18245 27591
rect 18245 27557 18279 27591
rect 18279 27557 18288 27591
rect 18236 27548 18288 27557
rect 21640 27591 21692 27600
rect 21640 27557 21649 27591
rect 21649 27557 21683 27591
rect 21683 27557 21692 27591
rect 21640 27548 21692 27557
rect 23664 27548 23716 27600
rect 11796 27344 11848 27396
rect 13176 27412 13228 27464
rect 14740 27480 14792 27532
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15384 27412 15436 27421
rect 16488 27412 16540 27464
rect 17408 27480 17460 27532
rect 18696 27523 18748 27532
rect 18696 27489 18705 27523
rect 18705 27489 18739 27523
rect 18739 27489 18748 27523
rect 18696 27480 18748 27489
rect 17316 27412 17368 27464
rect 17960 27455 18012 27464
rect 17960 27421 17969 27455
rect 17969 27421 18003 27455
rect 18003 27421 18012 27455
rect 17960 27412 18012 27421
rect 20444 27523 20496 27532
rect 20444 27489 20453 27523
rect 20453 27489 20487 27523
rect 20487 27489 20496 27523
rect 20444 27480 20496 27489
rect 20536 27523 20588 27532
rect 20536 27489 20545 27523
rect 20545 27489 20579 27523
rect 20579 27489 20588 27523
rect 20536 27480 20588 27489
rect 21088 27480 21140 27532
rect 23296 27480 23348 27532
rect 24032 27523 24084 27532
rect 24032 27489 24041 27523
rect 24041 27489 24075 27523
rect 24075 27489 24084 27523
rect 24032 27480 24084 27489
rect 11336 27276 11388 27328
rect 11980 27276 12032 27328
rect 14280 27344 14332 27396
rect 15108 27344 15160 27396
rect 21732 27412 21784 27464
rect 22744 27412 22796 27464
rect 22468 27344 22520 27396
rect 22560 27344 22612 27396
rect 23480 27412 23532 27464
rect 24400 27480 24452 27532
rect 24492 27523 24544 27532
rect 24492 27489 24501 27523
rect 24501 27489 24535 27523
rect 24535 27489 24544 27523
rect 24492 27480 24544 27489
rect 25044 27659 25096 27668
rect 25044 27625 25053 27659
rect 25053 27625 25087 27659
rect 25087 27625 25096 27659
rect 25044 27616 25096 27625
rect 24860 27548 24912 27600
rect 24216 27412 24268 27464
rect 24676 27344 24728 27396
rect 19800 27276 19852 27328
rect 20260 27319 20312 27328
rect 20260 27285 20269 27319
rect 20269 27285 20303 27319
rect 20303 27285 20312 27319
rect 20260 27276 20312 27285
rect 20812 27319 20864 27328
rect 20812 27285 20821 27319
rect 20821 27285 20855 27319
rect 20855 27285 20864 27319
rect 20812 27276 20864 27285
rect 21456 27276 21508 27328
rect 22376 27276 22428 27328
rect 22744 27276 22796 27328
rect 23020 27276 23072 27328
rect 24124 27276 24176 27328
rect 24584 27319 24636 27328
rect 24584 27285 24593 27319
rect 24593 27285 24627 27319
rect 24627 27285 24636 27319
rect 24584 27276 24636 27285
rect 25136 27523 25188 27532
rect 25136 27489 25145 27523
rect 25145 27489 25179 27523
rect 25179 27489 25188 27523
rect 25136 27480 25188 27489
rect 25228 27480 25280 27532
rect 25780 27455 25832 27464
rect 25780 27421 25789 27455
rect 25789 27421 25823 27455
rect 25823 27421 25832 27455
rect 25780 27412 25832 27421
rect 25872 27344 25924 27396
rect 26056 27387 26108 27396
rect 26056 27353 26065 27387
rect 26065 27353 26099 27387
rect 26099 27353 26108 27387
rect 26056 27344 26108 27353
rect 27528 27480 27580 27532
rect 28356 27480 28408 27532
rect 26332 27412 26384 27464
rect 26700 27412 26752 27464
rect 28080 27412 28132 27464
rect 27528 27344 27580 27396
rect 26332 27276 26384 27328
rect 26424 27319 26476 27328
rect 26424 27285 26433 27319
rect 26433 27285 26467 27319
rect 26467 27285 26476 27319
rect 26424 27276 26476 27285
rect 26884 27276 26936 27328
rect 29092 27319 29144 27328
rect 29092 27285 29101 27319
rect 29101 27285 29135 27319
rect 29135 27285 29144 27319
rect 29092 27276 29144 27285
rect 3662 27174 3714 27226
rect 3726 27174 3778 27226
rect 3790 27174 3842 27226
rect 3854 27174 3906 27226
rect 3918 27174 3970 27226
rect 11436 27174 11488 27226
rect 11500 27174 11552 27226
rect 11564 27174 11616 27226
rect 11628 27174 11680 27226
rect 11692 27174 11744 27226
rect 19210 27174 19262 27226
rect 19274 27174 19326 27226
rect 19338 27174 19390 27226
rect 19402 27174 19454 27226
rect 19466 27174 19518 27226
rect 26984 27174 27036 27226
rect 27048 27174 27100 27226
rect 27112 27174 27164 27226
rect 27176 27174 27228 27226
rect 27240 27174 27292 27226
rect 12532 27115 12584 27124
rect 12532 27081 12541 27115
rect 12541 27081 12575 27115
rect 12575 27081 12584 27115
rect 12532 27072 12584 27081
rect 14004 27072 14056 27124
rect 20720 27072 20772 27124
rect 24216 27072 24268 27124
rect 26148 27072 26200 27124
rect 26332 27115 26384 27124
rect 26332 27081 26341 27115
rect 26341 27081 26375 27115
rect 26375 27081 26384 27115
rect 26332 27072 26384 27081
rect 26424 27115 26476 27124
rect 26424 27081 26433 27115
rect 26433 27081 26467 27115
rect 26467 27081 26476 27115
rect 26424 27072 26476 27081
rect 26792 27115 26844 27124
rect 26792 27081 26801 27115
rect 26801 27081 26835 27115
rect 26835 27081 26844 27115
rect 26792 27072 26844 27081
rect 17776 27004 17828 27056
rect 24952 27004 25004 27056
rect 11244 26868 11296 26920
rect 11428 26911 11480 26920
rect 11428 26877 11462 26911
rect 11462 26877 11480 26911
rect 11428 26868 11480 26877
rect 13728 26868 13780 26920
rect 14280 26911 14332 26920
rect 14280 26877 14289 26911
rect 14289 26877 14323 26911
rect 14323 26877 14332 26911
rect 14280 26868 14332 26877
rect 14556 26911 14608 26920
rect 14556 26877 14565 26911
rect 14565 26877 14599 26911
rect 14599 26877 14608 26911
rect 14556 26868 14608 26877
rect 22468 26936 22520 26988
rect 17040 26868 17092 26920
rect 17960 26868 18012 26920
rect 18512 26868 18564 26920
rect 19616 26911 19668 26920
rect 19616 26877 19625 26911
rect 19625 26877 19659 26911
rect 19659 26877 19668 26911
rect 19616 26868 19668 26877
rect 20260 26868 20312 26920
rect 21180 26911 21232 26920
rect 21180 26877 21189 26911
rect 21189 26877 21223 26911
rect 21223 26877 21232 26911
rect 21180 26868 21232 26877
rect 21456 26911 21508 26920
rect 21456 26877 21490 26911
rect 21490 26877 21508 26911
rect 21456 26868 21508 26877
rect 22744 26868 22796 26920
rect 23020 26911 23072 26920
rect 23020 26877 23029 26911
rect 23029 26877 23063 26911
rect 23063 26877 23072 26911
rect 23020 26868 23072 26877
rect 23296 26911 23348 26920
rect 23296 26877 23305 26911
rect 23305 26877 23339 26911
rect 23339 26877 23348 26911
rect 23296 26868 23348 26877
rect 23388 26868 23440 26920
rect 24124 26911 24176 26920
rect 24124 26877 24158 26911
rect 24158 26877 24176 26911
rect 24124 26868 24176 26877
rect 24400 26868 24452 26920
rect 25228 26868 25280 26920
rect 25320 26868 25372 26920
rect 26056 26911 26108 26920
rect 26056 26877 26065 26911
rect 26065 26877 26099 26911
rect 26099 26877 26108 26911
rect 26056 26868 26108 26877
rect 26332 26868 26384 26920
rect 27988 26868 28040 26920
rect 20536 26800 20588 26852
rect 22376 26800 22428 26852
rect 13912 26732 13964 26784
rect 14188 26732 14240 26784
rect 16948 26775 17000 26784
rect 16948 26741 16957 26775
rect 16957 26741 16991 26775
rect 16991 26741 17000 26775
rect 16948 26732 17000 26741
rect 17500 26732 17552 26784
rect 18328 26732 18380 26784
rect 20996 26732 21048 26784
rect 22008 26732 22060 26784
rect 22560 26775 22612 26784
rect 22560 26741 22569 26775
rect 22569 26741 22603 26775
rect 22603 26741 22612 26775
rect 22560 26732 22612 26741
rect 22652 26775 22704 26784
rect 22652 26741 22661 26775
rect 22661 26741 22695 26775
rect 22695 26741 22704 26775
rect 22652 26732 22704 26741
rect 22744 26732 22796 26784
rect 26516 26800 26568 26852
rect 23572 26732 23624 26784
rect 24584 26732 24636 26784
rect 24768 26732 24820 26784
rect 25412 26732 25464 26784
rect 25872 26732 25924 26784
rect 28448 26800 28500 26852
rect 29092 26800 29144 26852
rect 26700 26732 26752 26784
rect 27528 26732 27580 26784
rect 4322 26630 4374 26682
rect 4386 26630 4438 26682
rect 4450 26630 4502 26682
rect 4514 26630 4566 26682
rect 4578 26630 4630 26682
rect 12096 26630 12148 26682
rect 12160 26630 12212 26682
rect 12224 26630 12276 26682
rect 12288 26630 12340 26682
rect 12352 26630 12404 26682
rect 19870 26630 19922 26682
rect 19934 26630 19986 26682
rect 19998 26630 20050 26682
rect 20062 26630 20114 26682
rect 20126 26630 20178 26682
rect 27644 26630 27696 26682
rect 27708 26630 27760 26682
rect 27772 26630 27824 26682
rect 27836 26630 27888 26682
rect 27900 26630 27952 26682
rect 13820 26528 13872 26580
rect 14740 26571 14792 26580
rect 14740 26537 14749 26571
rect 14749 26537 14783 26571
rect 14783 26537 14792 26571
rect 14740 26528 14792 26537
rect 17040 26571 17092 26580
rect 17040 26537 17049 26571
rect 17049 26537 17083 26571
rect 17083 26537 17092 26571
rect 17040 26528 17092 26537
rect 17316 26528 17368 26580
rect 17500 26571 17552 26580
rect 17500 26537 17509 26571
rect 17509 26537 17543 26571
rect 17543 26537 17552 26571
rect 17500 26528 17552 26537
rect 18144 26528 18196 26580
rect 18328 26571 18380 26580
rect 18328 26537 18337 26571
rect 18337 26537 18371 26571
rect 18371 26537 18380 26571
rect 18328 26528 18380 26537
rect 18420 26528 18472 26580
rect 19708 26571 19760 26580
rect 19708 26537 19717 26571
rect 19717 26537 19751 26571
rect 19751 26537 19760 26571
rect 19708 26528 19760 26537
rect 20444 26528 20496 26580
rect 15292 26460 15344 26512
rect 16764 26435 16816 26444
rect 16764 26401 16773 26435
rect 16773 26401 16807 26435
rect 16807 26401 16816 26435
rect 16764 26392 16816 26401
rect 12624 26367 12676 26376
rect 12624 26333 12633 26367
rect 12633 26333 12667 26367
rect 12667 26333 12676 26367
rect 12624 26324 12676 26333
rect 12808 26367 12860 26376
rect 12808 26333 12817 26367
rect 12817 26333 12851 26367
rect 12851 26333 12860 26367
rect 12808 26324 12860 26333
rect 13176 26324 13228 26376
rect 13636 26367 13688 26376
rect 13636 26333 13670 26367
rect 13670 26333 13688 26367
rect 13636 26324 13688 26333
rect 14188 26324 14240 26376
rect 15200 26367 15252 26376
rect 15200 26333 15209 26367
rect 15209 26333 15243 26367
rect 15243 26333 15252 26367
rect 15200 26324 15252 26333
rect 18052 26324 18104 26376
rect 19616 26460 19668 26512
rect 20352 26460 20404 26512
rect 20444 26435 20496 26444
rect 20444 26401 20453 26435
rect 20453 26401 20487 26435
rect 20487 26401 20496 26435
rect 20444 26392 20496 26401
rect 13912 26188 13964 26240
rect 15016 26188 15068 26240
rect 18144 26256 18196 26308
rect 16580 26188 16632 26240
rect 17868 26231 17920 26240
rect 17868 26197 17877 26231
rect 17877 26197 17911 26231
rect 17911 26197 17920 26231
rect 17868 26188 17920 26197
rect 18696 26231 18748 26240
rect 18696 26197 18705 26231
rect 18705 26197 18739 26231
rect 18739 26197 18748 26231
rect 18696 26188 18748 26197
rect 19064 26256 19116 26308
rect 20996 26392 21048 26444
rect 21180 26528 21232 26580
rect 22284 26528 22336 26580
rect 23112 26528 23164 26580
rect 23296 26528 23348 26580
rect 24032 26528 24084 26580
rect 26608 26528 26660 26580
rect 22192 26460 22244 26512
rect 22652 26460 22704 26512
rect 22836 26460 22888 26512
rect 24492 26460 24544 26512
rect 25504 26460 25556 26512
rect 26700 26503 26752 26512
rect 26700 26469 26709 26503
rect 26709 26469 26743 26503
rect 26743 26469 26752 26503
rect 26700 26460 26752 26469
rect 26792 26503 26844 26512
rect 26792 26469 26801 26503
rect 26801 26469 26835 26503
rect 26835 26469 26844 26503
rect 26792 26460 26844 26469
rect 27712 26460 27764 26512
rect 28172 26528 28224 26580
rect 28356 26571 28408 26580
rect 28356 26537 28365 26571
rect 28365 26537 28399 26571
rect 28399 26537 28408 26571
rect 28356 26528 28408 26537
rect 23388 26392 23440 26444
rect 20904 26367 20956 26376
rect 20904 26333 20913 26367
rect 20913 26333 20947 26367
rect 20947 26333 20956 26367
rect 20904 26324 20956 26333
rect 23572 26324 23624 26376
rect 18880 26188 18932 26240
rect 20720 26256 20772 26308
rect 20812 26256 20864 26308
rect 21640 26256 21692 26308
rect 19800 26188 19852 26240
rect 23480 26188 23532 26240
rect 23572 26188 23624 26240
rect 23756 26188 23808 26240
rect 26332 26392 26384 26444
rect 26424 26435 26476 26444
rect 26424 26401 26433 26435
rect 26433 26401 26467 26435
rect 26467 26401 26476 26435
rect 26424 26392 26476 26401
rect 26516 26435 26568 26444
rect 26516 26401 26526 26435
rect 26526 26401 26560 26435
rect 26560 26401 26568 26435
rect 26516 26392 26568 26401
rect 26884 26435 26936 26444
rect 26884 26401 26898 26435
rect 26898 26401 26932 26435
rect 26932 26401 26936 26435
rect 26884 26392 26936 26401
rect 27528 26392 27580 26444
rect 26056 26256 26108 26308
rect 26332 26256 26384 26308
rect 27896 26324 27948 26376
rect 28264 26324 28316 26376
rect 26792 26256 26844 26308
rect 28080 26256 28132 26308
rect 28172 26256 28224 26308
rect 28448 26256 28500 26308
rect 28908 26188 28960 26240
rect 3662 26086 3714 26138
rect 3726 26086 3778 26138
rect 3790 26086 3842 26138
rect 3854 26086 3906 26138
rect 3918 26086 3970 26138
rect 11436 26086 11488 26138
rect 11500 26086 11552 26138
rect 11564 26086 11616 26138
rect 11628 26086 11680 26138
rect 11692 26086 11744 26138
rect 19210 26086 19262 26138
rect 19274 26086 19326 26138
rect 19338 26086 19390 26138
rect 19402 26086 19454 26138
rect 19466 26086 19518 26138
rect 26984 26086 27036 26138
rect 27048 26086 27100 26138
rect 27112 26086 27164 26138
rect 27176 26086 27228 26138
rect 27240 26086 27292 26138
rect 12992 26027 13044 26036
rect 12992 25993 13001 26027
rect 13001 25993 13035 26027
rect 13035 25993 13044 26027
rect 12992 25984 13044 25993
rect 14556 25984 14608 26036
rect 15292 26027 15344 26036
rect 15292 25993 15301 26027
rect 15301 25993 15335 26027
rect 15335 25993 15344 26027
rect 15292 25984 15344 25993
rect 15384 25984 15436 26036
rect 12624 25848 12676 25900
rect 13636 25848 13688 25900
rect 15016 25891 15068 25900
rect 15016 25857 15025 25891
rect 15025 25857 15059 25891
rect 15059 25857 15068 25891
rect 15016 25848 15068 25857
rect 11336 25780 11388 25832
rect 12808 25780 12860 25832
rect 13176 25823 13228 25832
rect 13176 25789 13185 25823
rect 13185 25789 13219 25823
rect 13219 25789 13228 25823
rect 13176 25780 13228 25789
rect 11888 25644 11940 25696
rect 14188 25687 14240 25696
rect 14188 25653 14197 25687
rect 14197 25653 14231 25687
rect 14231 25653 14240 25687
rect 14188 25644 14240 25653
rect 14280 25644 14332 25696
rect 15200 25780 15252 25832
rect 15752 25780 15804 25832
rect 16764 25984 16816 26036
rect 17132 25984 17184 26036
rect 17776 25916 17828 25968
rect 17960 25891 18012 25900
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 17960 25848 18012 25857
rect 15476 25712 15528 25764
rect 16580 25780 16632 25832
rect 17868 25780 17920 25832
rect 18512 26027 18564 26036
rect 18512 25993 18521 26027
rect 18521 25993 18555 26027
rect 18555 25993 18564 26027
rect 18512 25984 18564 25993
rect 20996 25984 21048 26036
rect 28816 25848 28868 25900
rect 19064 25823 19116 25832
rect 19064 25789 19073 25823
rect 19073 25789 19107 25823
rect 19107 25789 19116 25823
rect 19064 25780 19116 25789
rect 16488 25644 16540 25696
rect 18512 25712 18564 25764
rect 18972 25712 19024 25764
rect 19800 25823 19852 25832
rect 19800 25789 19809 25823
rect 19809 25789 19843 25823
rect 19843 25789 19852 25823
rect 19800 25780 19852 25789
rect 27896 25823 27948 25832
rect 27896 25789 27905 25823
rect 27905 25789 27939 25823
rect 27939 25789 27948 25823
rect 27896 25780 27948 25789
rect 28080 25780 28132 25832
rect 18144 25687 18196 25696
rect 18144 25653 18153 25687
rect 18153 25653 18187 25687
rect 18187 25653 18196 25687
rect 18144 25644 18196 25653
rect 18328 25644 18380 25696
rect 21364 25644 21416 25696
rect 23204 25644 23256 25696
rect 27528 25644 27580 25696
rect 28172 25644 28224 25696
rect 4322 25542 4374 25594
rect 4386 25542 4438 25594
rect 4450 25542 4502 25594
rect 4514 25542 4566 25594
rect 4578 25542 4630 25594
rect 12096 25542 12148 25594
rect 12160 25542 12212 25594
rect 12224 25542 12276 25594
rect 12288 25542 12340 25594
rect 12352 25542 12404 25594
rect 19870 25542 19922 25594
rect 19934 25542 19986 25594
rect 19998 25542 20050 25594
rect 20062 25542 20114 25594
rect 20126 25542 20178 25594
rect 27644 25542 27696 25594
rect 27708 25542 27760 25594
rect 27772 25542 27824 25594
rect 27836 25542 27888 25594
rect 27900 25542 27952 25594
rect 13176 25440 13228 25492
rect 11888 25347 11940 25356
rect 11888 25313 11897 25347
rect 11897 25313 11931 25347
rect 11931 25313 11940 25347
rect 11888 25304 11940 25313
rect 13084 25304 13136 25356
rect 17960 25440 18012 25492
rect 24860 25440 24912 25492
rect 26424 25440 26476 25492
rect 14188 25372 14240 25424
rect 15200 25372 15252 25424
rect 16948 25372 17000 25424
rect 18696 25372 18748 25424
rect 21640 25372 21692 25424
rect 23388 25415 23440 25424
rect 23388 25381 23397 25415
rect 23397 25381 23431 25415
rect 23431 25381 23440 25415
rect 23388 25372 23440 25381
rect 16212 25304 16264 25356
rect 16488 25347 16540 25356
rect 16488 25313 16497 25347
rect 16497 25313 16531 25347
rect 16531 25313 16540 25347
rect 16488 25304 16540 25313
rect 18328 25347 18380 25356
rect 18328 25313 18337 25347
rect 18337 25313 18371 25347
rect 18371 25313 18380 25347
rect 18328 25304 18380 25313
rect 20352 25304 20404 25356
rect 22284 25304 22336 25356
rect 15384 25236 15436 25288
rect 16028 25236 16080 25288
rect 21456 25236 21508 25288
rect 14004 25168 14056 25220
rect 14648 25100 14700 25152
rect 15568 25100 15620 25152
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 19064 25100 19116 25152
rect 20260 25100 20312 25152
rect 22100 25143 22152 25152
rect 22100 25109 22109 25143
rect 22109 25109 22143 25143
rect 22143 25109 22152 25143
rect 22100 25100 22152 25109
rect 22376 25143 22428 25152
rect 22376 25109 22385 25143
rect 22385 25109 22419 25143
rect 22419 25109 22428 25143
rect 22376 25100 22428 25109
rect 22836 25347 22888 25356
rect 22836 25313 22871 25347
rect 22871 25313 22888 25347
rect 22836 25304 22888 25313
rect 23480 25347 23532 25356
rect 23480 25313 23489 25347
rect 23489 25313 23523 25347
rect 23523 25313 23532 25347
rect 23480 25304 23532 25313
rect 23572 25347 23624 25356
rect 23572 25313 23581 25347
rect 23581 25313 23615 25347
rect 23615 25313 23624 25347
rect 23572 25304 23624 25313
rect 24124 25372 24176 25424
rect 25228 25372 25280 25424
rect 26148 25372 26200 25424
rect 23020 25279 23072 25288
rect 23020 25245 23029 25279
rect 23029 25245 23063 25279
rect 23063 25245 23072 25279
rect 23020 25236 23072 25245
rect 25320 25236 25372 25288
rect 22928 25168 22980 25220
rect 23204 25168 23256 25220
rect 24492 25168 24544 25220
rect 24676 25168 24728 25220
rect 27988 25304 28040 25356
rect 28632 25304 28684 25356
rect 23572 25100 23624 25152
rect 23756 25143 23808 25152
rect 23756 25109 23765 25143
rect 23765 25109 23799 25143
rect 23799 25109 23808 25143
rect 23756 25100 23808 25109
rect 24032 25143 24084 25152
rect 24032 25109 24041 25143
rect 24041 25109 24075 25143
rect 24075 25109 24084 25143
rect 24032 25100 24084 25109
rect 24860 25100 24912 25152
rect 27620 25143 27672 25152
rect 27620 25109 27629 25143
rect 27629 25109 27663 25143
rect 27663 25109 27672 25143
rect 27620 25100 27672 25109
rect 3662 24998 3714 25050
rect 3726 24998 3778 25050
rect 3790 24998 3842 25050
rect 3854 24998 3906 25050
rect 3918 24998 3970 25050
rect 11436 24998 11488 25050
rect 11500 24998 11552 25050
rect 11564 24998 11616 25050
rect 11628 24998 11680 25050
rect 11692 24998 11744 25050
rect 19210 24998 19262 25050
rect 19274 24998 19326 25050
rect 19338 24998 19390 25050
rect 19402 24998 19454 25050
rect 19466 24998 19518 25050
rect 26984 24998 27036 25050
rect 27048 24998 27100 25050
rect 27112 24998 27164 25050
rect 27176 24998 27228 25050
rect 27240 24998 27292 25050
rect 12992 24939 13044 24948
rect 12992 24905 13001 24939
rect 13001 24905 13035 24939
rect 13035 24905 13044 24939
rect 12992 24896 13044 24905
rect 16028 24939 16080 24948
rect 16028 24905 16037 24939
rect 16037 24905 16071 24939
rect 16071 24905 16080 24939
rect 16028 24896 16080 24905
rect 21732 24896 21784 24948
rect 22836 24896 22888 24948
rect 22928 24896 22980 24948
rect 24032 24896 24084 24948
rect 27436 24896 27488 24948
rect 28816 24939 28868 24948
rect 28816 24905 28825 24939
rect 28825 24905 28859 24939
rect 28859 24905 28868 24939
rect 28816 24896 28868 24905
rect 11336 24735 11388 24744
rect 11336 24701 11345 24735
rect 11345 24701 11379 24735
rect 11379 24701 11388 24735
rect 11336 24692 11388 24701
rect 13820 24735 13872 24744
rect 13820 24701 13829 24735
rect 13829 24701 13863 24735
rect 13863 24701 13872 24735
rect 13820 24692 13872 24701
rect 13912 24735 13964 24744
rect 13912 24701 13921 24735
rect 13921 24701 13955 24735
rect 13955 24701 13964 24735
rect 13912 24692 13964 24701
rect 14004 24735 14056 24744
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 14004 24692 14056 24701
rect 13728 24556 13780 24608
rect 14372 24735 14424 24744
rect 14372 24701 14381 24735
rect 14381 24701 14415 24735
rect 14415 24701 14424 24735
rect 14372 24692 14424 24701
rect 17684 24803 17736 24812
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 17960 24828 18012 24880
rect 26608 24828 26660 24880
rect 15016 24624 15068 24676
rect 17960 24692 18012 24744
rect 18512 24760 18564 24812
rect 18972 24760 19024 24812
rect 19064 24735 19116 24744
rect 19064 24701 19073 24735
rect 19073 24701 19107 24735
rect 19107 24701 19116 24735
rect 19064 24692 19116 24701
rect 20260 24803 20312 24812
rect 20260 24769 20269 24803
rect 20269 24769 20303 24803
rect 20303 24769 20312 24803
rect 20260 24760 20312 24769
rect 24492 24803 24544 24812
rect 24492 24769 24501 24803
rect 24501 24769 24535 24803
rect 24535 24769 24544 24803
rect 24492 24760 24544 24769
rect 19800 24735 19852 24744
rect 19800 24701 19809 24735
rect 19809 24701 19843 24735
rect 19843 24701 19852 24735
rect 19800 24692 19852 24701
rect 22008 24692 22060 24744
rect 23112 24692 23164 24744
rect 23756 24692 23808 24744
rect 20260 24624 20312 24676
rect 20352 24624 20404 24676
rect 15292 24556 15344 24608
rect 16212 24556 16264 24608
rect 21732 24624 21784 24676
rect 22284 24624 22336 24676
rect 23664 24624 23716 24676
rect 25044 24735 25096 24744
rect 25044 24701 25053 24735
rect 25053 24701 25087 24735
rect 25087 24701 25096 24735
rect 25044 24692 25096 24701
rect 25228 24735 25280 24744
rect 25228 24701 25237 24735
rect 25237 24701 25271 24735
rect 25271 24701 25280 24735
rect 25228 24692 25280 24701
rect 25320 24735 25372 24744
rect 25320 24701 25329 24735
rect 25329 24701 25363 24735
rect 25363 24701 25372 24735
rect 25320 24692 25372 24701
rect 25504 24692 25556 24744
rect 25596 24735 25648 24744
rect 25596 24701 25605 24735
rect 25605 24701 25639 24735
rect 25639 24701 25648 24735
rect 25596 24692 25648 24701
rect 24676 24624 24728 24676
rect 26056 24735 26108 24744
rect 26056 24701 26065 24735
rect 26065 24701 26099 24735
rect 26099 24701 26108 24735
rect 26056 24692 26108 24701
rect 25780 24624 25832 24676
rect 21640 24599 21692 24608
rect 21640 24565 21649 24599
rect 21649 24565 21683 24599
rect 21683 24565 21692 24599
rect 21640 24556 21692 24565
rect 22468 24556 22520 24608
rect 23020 24556 23072 24608
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 23756 24556 23808 24608
rect 25412 24556 25464 24608
rect 26792 24692 26844 24744
rect 27528 24692 27580 24744
rect 26332 24624 26384 24676
rect 26700 24667 26752 24676
rect 26700 24633 26709 24667
rect 26709 24633 26743 24667
rect 26743 24633 26752 24667
rect 26700 24624 26752 24633
rect 26424 24556 26476 24608
rect 27068 24599 27120 24608
rect 27068 24565 27077 24599
rect 27077 24565 27111 24599
rect 27111 24565 27120 24599
rect 27068 24556 27120 24565
rect 27528 24556 27580 24608
rect 4322 24454 4374 24506
rect 4386 24454 4438 24506
rect 4450 24454 4502 24506
rect 4514 24454 4566 24506
rect 4578 24454 4630 24506
rect 12096 24454 12148 24506
rect 12160 24454 12212 24506
rect 12224 24454 12276 24506
rect 12288 24454 12340 24506
rect 12352 24454 12404 24506
rect 19870 24454 19922 24506
rect 19934 24454 19986 24506
rect 19998 24454 20050 24506
rect 20062 24454 20114 24506
rect 20126 24454 20178 24506
rect 27644 24454 27696 24506
rect 27708 24454 27760 24506
rect 27772 24454 27824 24506
rect 27836 24454 27888 24506
rect 27900 24454 27952 24506
rect 13084 24395 13136 24404
rect 13084 24361 13093 24395
rect 13093 24361 13127 24395
rect 13127 24361 13136 24395
rect 13084 24352 13136 24361
rect 14648 24327 14700 24336
rect 14648 24293 14657 24327
rect 14657 24293 14691 24327
rect 14691 24293 14700 24327
rect 14648 24284 14700 24293
rect 13728 24259 13780 24268
rect 13728 24225 13737 24259
rect 13737 24225 13771 24259
rect 13771 24225 13780 24259
rect 13728 24216 13780 24225
rect 14280 24216 14332 24268
rect 15844 24284 15896 24336
rect 20352 24395 20404 24404
rect 20352 24361 20361 24395
rect 20361 24361 20395 24395
rect 20395 24361 20404 24395
rect 20352 24352 20404 24361
rect 20996 24284 21048 24336
rect 21640 24352 21692 24404
rect 22284 24352 22336 24404
rect 23572 24352 23624 24404
rect 24676 24395 24728 24404
rect 24676 24361 24685 24395
rect 24685 24361 24719 24395
rect 24719 24361 24728 24395
rect 24676 24352 24728 24361
rect 25044 24352 25096 24404
rect 25504 24352 25556 24404
rect 27528 24395 27580 24404
rect 27528 24361 27537 24395
rect 27537 24361 27571 24395
rect 27571 24361 27580 24395
rect 27528 24352 27580 24361
rect 28264 24352 28316 24404
rect 28540 24352 28592 24404
rect 13912 24148 13964 24200
rect 12992 24080 13044 24132
rect 15568 24259 15620 24268
rect 15568 24225 15577 24259
rect 15577 24225 15611 24259
rect 15611 24225 15620 24259
rect 15568 24216 15620 24225
rect 16212 24216 16264 24268
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 16488 24216 16540 24268
rect 18972 24148 19024 24200
rect 21732 24327 21784 24336
rect 21732 24293 21767 24327
rect 21767 24293 21784 24327
rect 21732 24284 21784 24293
rect 21456 24259 21508 24268
rect 21456 24225 21465 24259
rect 21465 24225 21499 24259
rect 21499 24225 21508 24259
rect 21456 24216 21508 24225
rect 21640 24259 21692 24268
rect 21640 24225 21649 24259
rect 21649 24225 21683 24259
rect 21683 24225 21692 24259
rect 21640 24216 21692 24225
rect 22376 24284 22428 24336
rect 23480 24284 23532 24336
rect 23756 24259 23808 24268
rect 26148 24284 26200 24336
rect 27344 24284 27396 24336
rect 27620 24284 27672 24336
rect 28448 24284 28500 24336
rect 23756 24225 23774 24259
rect 23774 24225 23808 24259
rect 23756 24216 23808 24225
rect 24308 24259 24360 24268
rect 24308 24225 24317 24259
rect 24317 24225 24351 24259
rect 24351 24225 24360 24259
rect 24308 24216 24360 24225
rect 15200 24080 15252 24132
rect 16488 24080 16540 24132
rect 21732 24148 21784 24200
rect 21364 24080 21416 24132
rect 24124 24148 24176 24200
rect 24860 24191 24912 24200
rect 24860 24157 24869 24191
rect 24869 24157 24903 24191
rect 24903 24157 24912 24191
rect 24860 24148 24912 24157
rect 25412 24259 25464 24268
rect 25412 24225 25421 24259
rect 25421 24225 25455 24259
rect 25455 24225 25464 24259
rect 25412 24216 25464 24225
rect 25596 24216 25648 24268
rect 25780 24259 25832 24268
rect 25780 24225 25789 24259
rect 25789 24225 25823 24259
rect 25823 24225 25832 24259
rect 25780 24216 25832 24225
rect 26056 24216 26108 24268
rect 26424 24216 26476 24268
rect 26608 24259 26660 24268
rect 26608 24225 26617 24259
rect 26617 24225 26651 24259
rect 26651 24225 26660 24259
rect 26608 24216 26660 24225
rect 27528 24216 27580 24268
rect 27344 24148 27396 24200
rect 28356 24259 28408 24268
rect 28356 24225 28365 24259
rect 28365 24225 28399 24259
rect 28399 24225 28408 24259
rect 28356 24216 28408 24225
rect 28724 24216 28776 24268
rect 14004 24055 14056 24064
rect 14004 24021 14013 24055
rect 14013 24021 14047 24055
rect 14047 24021 14056 24055
rect 14004 24012 14056 24021
rect 15016 24012 15068 24064
rect 16304 24012 16356 24064
rect 26240 24080 26292 24132
rect 28080 24123 28132 24132
rect 28080 24089 28089 24123
rect 28089 24089 28123 24123
rect 28123 24089 28132 24123
rect 28080 24080 28132 24089
rect 23664 24012 23716 24064
rect 27068 24012 27120 24064
rect 28172 24012 28224 24064
rect 28356 24012 28408 24064
rect 3662 23910 3714 23962
rect 3726 23910 3778 23962
rect 3790 23910 3842 23962
rect 3854 23910 3906 23962
rect 3918 23910 3970 23962
rect 11436 23910 11488 23962
rect 11500 23910 11552 23962
rect 11564 23910 11616 23962
rect 11628 23910 11680 23962
rect 11692 23910 11744 23962
rect 19210 23910 19262 23962
rect 19274 23910 19326 23962
rect 19338 23910 19390 23962
rect 19402 23910 19454 23962
rect 19466 23910 19518 23962
rect 26984 23910 27036 23962
rect 27048 23910 27100 23962
rect 27112 23910 27164 23962
rect 27176 23910 27228 23962
rect 27240 23910 27292 23962
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 13636 23740 13688 23792
rect 14188 23672 14240 23724
rect 11336 23604 11388 23656
rect 14372 23604 14424 23656
rect 16120 23740 16172 23792
rect 19708 23808 19760 23860
rect 20352 23851 20404 23860
rect 20352 23817 20361 23851
rect 20361 23817 20395 23851
rect 20395 23817 20404 23851
rect 20352 23808 20404 23817
rect 20812 23808 20864 23860
rect 25964 23808 26016 23860
rect 28080 23808 28132 23860
rect 28356 23851 28408 23860
rect 28356 23817 28365 23851
rect 28365 23817 28399 23851
rect 28399 23817 28408 23851
rect 28356 23808 28408 23817
rect 28724 23808 28776 23860
rect 17040 23740 17092 23792
rect 17868 23672 17920 23724
rect 12992 23579 13044 23588
rect 12992 23545 13001 23579
rect 13001 23545 13035 23579
rect 13035 23545 13044 23579
rect 12992 23536 13044 23545
rect 12440 23511 12492 23520
rect 12440 23477 12449 23511
rect 12449 23477 12483 23511
rect 12483 23477 12492 23511
rect 12440 23468 12492 23477
rect 14648 23579 14700 23588
rect 14648 23545 14657 23579
rect 14657 23545 14691 23579
rect 14691 23545 14700 23579
rect 14648 23536 14700 23545
rect 15200 23468 15252 23520
rect 15844 23647 15896 23656
rect 15844 23613 15853 23647
rect 15853 23613 15887 23647
rect 15887 23613 15896 23647
rect 15844 23604 15896 23613
rect 15936 23647 15988 23656
rect 15936 23613 15945 23647
rect 15945 23613 15979 23647
rect 15979 23613 15988 23647
rect 15936 23604 15988 23613
rect 16120 23647 16172 23656
rect 16120 23613 16129 23647
rect 16129 23613 16163 23647
rect 16163 23613 16172 23647
rect 16120 23604 16172 23613
rect 16212 23604 16264 23656
rect 17132 23647 17184 23656
rect 17132 23613 17141 23647
rect 17141 23613 17175 23647
rect 17175 23613 17184 23647
rect 17132 23604 17184 23613
rect 18788 23604 18840 23656
rect 19064 23647 19116 23656
rect 19064 23613 19073 23647
rect 19073 23613 19107 23647
rect 19107 23613 19116 23647
rect 19064 23604 19116 23613
rect 16488 23536 16540 23588
rect 17960 23536 18012 23588
rect 18144 23536 18196 23588
rect 24584 23604 24636 23656
rect 28448 23740 28500 23792
rect 27620 23672 27672 23724
rect 28264 23672 28316 23724
rect 17040 23468 17092 23520
rect 17592 23468 17644 23520
rect 18788 23468 18840 23520
rect 19248 23536 19300 23588
rect 19800 23536 19852 23588
rect 28172 23604 28224 23656
rect 28632 23647 28684 23656
rect 28632 23613 28641 23647
rect 28641 23613 28675 23647
rect 28675 23613 28684 23647
rect 28632 23604 28684 23613
rect 19156 23511 19208 23520
rect 19156 23477 19165 23511
rect 19165 23477 19199 23511
rect 19199 23477 19208 23511
rect 19156 23468 19208 23477
rect 28080 23468 28132 23520
rect 28356 23511 28408 23520
rect 28356 23477 28365 23511
rect 28365 23477 28399 23511
rect 28399 23477 28408 23511
rect 28356 23468 28408 23477
rect 4322 23366 4374 23418
rect 4386 23366 4438 23418
rect 4450 23366 4502 23418
rect 4514 23366 4566 23418
rect 4578 23366 4630 23418
rect 12096 23366 12148 23418
rect 12160 23366 12212 23418
rect 12224 23366 12276 23418
rect 12288 23366 12340 23418
rect 12352 23366 12404 23418
rect 19870 23366 19922 23418
rect 19934 23366 19986 23418
rect 19998 23366 20050 23418
rect 20062 23366 20114 23418
rect 20126 23366 20178 23418
rect 27644 23366 27696 23418
rect 27708 23366 27760 23418
rect 27772 23366 27824 23418
rect 27836 23366 27888 23418
rect 27900 23366 27952 23418
rect 12624 23264 12676 23316
rect 13636 23307 13688 23316
rect 13636 23273 13645 23307
rect 13645 23273 13679 23307
rect 13679 23273 13688 23307
rect 13636 23264 13688 23273
rect 13912 23196 13964 23248
rect 14372 23264 14424 23316
rect 12348 23128 12400 23180
rect 14188 23171 14240 23180
rect 14188 23137 14197 23171
rect 14197 23137 14231 23171
rect 14231 23137 14240 23171
rect 14188 23128 14240 23137
rect 15292 23196 15344 23248
rect 15752 23264 15804 23316
rect 16212 23307 16264 23316
rect 16212 23273 16221 23307
rect 16221 23273 16255 23307
rect 16255 23273 16264 23307
rect 16212 23264 16264 23273
rect 17868 23264 17920 23316
rect 22192 23264 22244 23316
rect 16488 23196 16540 23248
rect 17132 23196 17184 23248
rect 17684 23196 17736 23248
rect 14648 23171 14700 23180
rect 14648 23137 14657 23171
rect 14657 23137 14691 23171
rect 14691 23137 14700 23171
rect 14648 23128 14700 23137
rect 16856 23128 16908 23180
rect 17592 23171 17644 23180
rect 17592 23137 17601 23171
rect 17601 23137 17635 23171
rect 17635 23137 17644 23171
rect 17592 23128 17644 23137
rect 18696 23128 18748 23180
rect 18880 23171 18932 23180
rect 18880 23137 18889 23171
rect 18889 23137 18923 23171
rect 18923 23137 18932 23171
rect 18880 23128 18932 23137
rect 19156 23171 19208 23180
rect 19156 23137 19165 23171
rect 19165 23137 19199 23171
rect 19199 23137 19208 23171
rect 19156 23128 19208 23137
rect 19708 23128 19760 23180
rect 14832 23060 14884 23112
rect 22008 23196 22060 23248
rect 23388 23264 23440 23316
rect 23112 23239 23164 23248
rect 23112 23205 23121 23239
rect 23121 23205 23155 23239
rect 23155 23205 23164 23239
rect 26792 23264 26844 23316
rect 27436 23264 27488 23316
rect 23112 23196 23164 23205
rect 20720 23171 20772 23180
rect 20720 23137 20729 23171
rect 20729 23137 20763 23171
rect 20763 23137 20772 23171
rect 20720 23128 20772 23137
rect 20996 23171 21048 23180
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 21272 23171 21324 23180
rect 21272 23137 21281 23171
rect 21281 23137 21315 23171
rect 21315 23137 21324 23171
rect 21272 23128 21324 23137
rect 21364 23128 21416 23180
rect 21456 23060 21508 23112
rect 21640 23060 21692 23112
rect 22100 23171 22152 23180
rect 22100 23137 22109 23171
rect 22109 23137 22143 23171
rect 22143 23137 22152 23171
rect 22100 23128 22152 23137
rect 22560 23128 22612 23180
rect 25412 23196 25464 23248
rect 24032 23171 24084 23180
rect 24032 23137 24041 23171
rect 24041 23137 24075 23171
rect 24075 23137 24084 23171
rect 24032 23128 24084 23137
rect 24216 23171 24268 23180
rect 24216 23137 24225 23171
rect 24225 23137 24259 23171
rect 24259 23137 24268 23171
rect 24216 23128 24268 23137
rect 24676 23128 24728 23180
rect 27988 23196 28040 23248
rect 28080 23196 28132 23248
rect 28724 23264 28776 23316
rect 28540 23239 28592 23248
rect 28540 23205 28549 23239
rect 28549 23205 28583 23239
rect 28583 23205 28592 23239
rect 28540 23196 28592 23205
rect 24492 23103 24544 23112
rect 24492 23069 24501 23103
rect 24501 23069 24535 23103
rect 24535 23069 24544 23103
rect 24492 23060 24544 23069
rect 26332 23060 26384 23112
rect 27620 23171 27672 23180
rect 27620 23137 27629 23171
rect 27629 23137 27663 23171
rect 27663 23137 27672 23171
rect 27620 23128 27672 23137
rect 28908 23128 28960 23180
rect 28816 23060 28868 23112
rect 16580 22924 16632 22976
rect 19616 22992 19668 23044
rect 20352 22992 20404 23044
rect 22284 22992 22336 23044
rect 26884 22992 26936 23044
rect 27436 22992 27488 23044
rect 28264 22992 28316 23044
rect 28356 22992 28408 23044
rect 28724 23035 28776 23044
rect 28724 23001 28733 23035
rect 28733 23001 28767 23035
rect 28767 23001 28776 23035
rect 28724 22992 28776 23001
rect 18880 22924 18932 22976
rect 19708 22967 19760 22976
rect 19708 22933 19717 22967
rect 19717 22933 19751 22967
rect 19751 22933 19760 22967
rect 19708 22924 19760 22933
rect 19984 22967 20036 22976
rect 19984 22933 19993 22967
rect 19993 22933 20027 22967
rect 20027 22933 20036 22967
rect 19984 22924 20036 22933
rect 21180 22924 21232 22976
rect 23112 22924 23164 22976
rect 25320 22924 25372 22976
rect 26608 22924 26660 22976
rect 28080 22924 28132 22976
rect 28172 22967 28224 22976
rect 28172 22933 28181 22967
rect 28181 22933 28215 22967
rect 28215 22933 28224 22967
rect 28172 22924 28224 22933
rect 28816 22924 28868 22976
rect 3662 22822 3714 22874
rect 3726 22822 3778 22874
rect 3790 22822 3842 22874
rect 3854 22822 3906 22874
rect 3918 22822 3970 22874
rect 11436 22822 11488 22874
rect 11500 22822 11552 22874
rect 11564 22822 11616 22874
rect 11628 22822 11680 22874
rect 11692 22822 11744 22874
rect 19210 22822 19262 22874
rect 19274 22822 19326 22874
rect 19338 22822 19390 22874
rect 19402 22822 19454 22874
rect 19466 22822 19518 22874
rect 26984 22822 27036 22874
rect 27048 22822 27100 22874
rect 27112 22822 27164 22874
rect 27176 22822 27228 22874
rect 27240 22822 27292 22874
rect 14096 22652 14148 22704
rect 16120 22720 16172 22772
rect 16856 22763 16908 22772
rect 16856 22729 16865 22763
rect 16865 22729 16899 22763
rect 16899 22729 16908 22763
rect 16856 22720 16908 22729
rect 12992 22491 13044 22500
rect 12992 22457 13001 22491
rect 13001 22457 13035 22491
rect 13035 22457 13044 22491
rect 12992 22448 13044 22457
rect 14004 22559 14056 22568
rect 14004 22525 14013 22559
rect 14013 22525 14047 22559
rect 14047 22525 14056 22559
rect 14004 22516 14056 22525
rect 12716 22423 12768 22432
rect 12716 22389 12725 22423
rect 12725 22389 12759 22423
rect 12759 22389 12768 22423
rect 12716 22380 12768 22389
rect 12808 22380 12860 22432
rect 13912 22448 13964 22500
rect 14556 22559 14608 22568
rect 14556 22525 14565 22559
rect 14565 22525 14599 22559
rect 14599 22525 14608 22559
rect 14556 22516 14608 22525
rect 17684 22584 17736 22636
rect 17960 22584 18012 22636
rect 19708 22720 19760 22772
rect 21272 22720 21324 22772
rect 21456 22763 21508 22772
rect 21456 22729 21465 22763
rect 21465 22729 21499 22763
rect 21499 22729 21508 22763
rect 21456 22720 21508 22729
rect 20996 22652 21048 22704
rect 21824 22720 21876 22772
rect 14372 22448 14424 22500
rect 15200 22516 15252 22568
rect 15292 22516 15344 22568
rect 16304 22516 16356 22568
rect 16488 22559 16540 22568
rect 16488 22525 16497 22559
rect 16497 22525 16531 22559
rect 16531 22525 16540 22559
rect 16488 22516 16540 22525
rect 16580 22559 16632 22568
rect 16580 22525 16589 22559
rect 16589 22525 16623 22559
rect 16623 22525 16632 22559
rect 16580 22516 16632 22525
rect 17776 22516 17828 22568
rect 18144 22559 18196 22568
rect 18144 22525 18153 22559
rect 18153 22525 18187 22559
rect 18187 22525 18196 22559
rect 18144 22516 18196 22525
rect 20352 22584 20404 22636
rect 18420 22516 18472 22568
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 18788 22516 18840 22568
rect 19984 22516 20036 22568
rect 20812 22559 20864 22568
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 20812 22516 20864 22525
rect 21088 22559 21140 22568
rect 21088 22525 21097 22559
rect 21097 22525 21131 22559
rect 21131 22525 21140 22559
rect 21088 22516 21140 22525
rect 21180 22559 21232 22568
rect 21180 22525 21189 22559
rect 21189 22525 21223 22559
rect 21223 22525 21232 22559
rect 21180 22516 21232 22525
rect 22100 22652 22152 22704
rect 22192 22652 22244 22704
rect 22744 22652 22796 22704
rect 24492 22652 24544 22704
rect 22008 22559 22060 22568
rect 22008 22525 22043 22559
rect 22043 22525 22060 22559
rect 22008 22516 22060 22525
rect 22192 22559 22244 22568
rect 22192 22525 22201 22559
rect 22201 22525 22235 22559
rect 22235 22525 22244 22559
rect 22192 22516 22244 22525
rect 23020 22516 23072 22568
rect 17408 22448 17460 22500
rect 20720 22448 20772 22500
rect 24400 22559 24452 22568
rect 24400 22525 24409 22559
rect 24409 22525 24443 22559
rect 24443 22525 24452 22559
rect 24400 22516 24452 22525
rect 27436 22652 27488 22704
rect 26332 22584 26384 22636
rect 24676 22516 24728 22568
rect 27160 22584 27212 22636
rect 14004 22380 14056 22432
rect 14464 22423 14516 22432
rect 14464 22389 14473 22423
rect 14473 22389 14507 22423
rect 14507 22389 14516 22423
rect 14464 22380 14516 22389
rect 15476 22380 15528 22432
rect 16212 22380 16264 22432
rect 16304 22380 16356 22432
rect 20444 22380 20496 22432
rect 21548 22423 21600 22432
rect 21548 22389 21557 22423
rect 21557 22389 21591 22423
rect 21591 22389 21600 22423
rect 21548 22380 21600 22389
rect 23204 22380 23256 22432
rect 23664 22380 23716 22432
rect 24032 22380 24084 22432
rect 24768 22380 24820 22432
rect 25136 22448 25188 22500
rect 27160 22448 27212 22500
rect 27436 22516 27488 22568
rect 28632 22516 28684 22568
rect 29000 22516 29052 22568
rect 26792 22380 26844 22432
rect 27988 22380 28040 22432
rect 28448 22380 28500 22432
rect 4322 22278 4374 22330
rect 4386 22278 4438 22330
rect 4450 22278 4502 22330
rect 4514 22278 4566 22330
rect 4578 22278 4630 22330
rect 12096 22278 12148 22330
rect 12160 22278 12212 22330
rect 12224 22278 12276 22330
rect 12288 22278 12340 22330
rect 12352 22278 12404 22330
rect 19870 22278 19922 22330
rect 19934 22278 19986 22330
rect 19998 22278 20050 22330
rect 20062 22278 20114 22330
rect 20126 22278 20178 22330
rect 27644 22278 27696 22330
rect 27708 22278 27760 22330
rect 27772 22278 27824 22330
rect 27836 22278 27888 22330
rect 27900 22278 27952 22330
rect 12808 22176 12860 22228
rect 13912 22176 13964 22228
rect 14648 22176 14700 22228
rect 12716 22108 12768 22160
rect 13636 22083 13688 22092
rect 14464 22108 14516 22160
rect 16304 22108 16356 22160
rect 18788 22176 18840 22228
rect 13636 22049 13654 22083
rect 13654 22049 13688 22083
rect 13636 22040 13688 22049
rect 14004 22083 14056 22092
rect 14004 22049 14013 22083
rect 14013 22049 14047 22083
rect 14047 22049 14056 22083
rect 14004 22040 14056 22049
rect 16212 22040 16264 22092
rect 17316 22083 17368 22092
rect 17316 22049 17325 22083
rect 17325 22049 17359 22083
rect 17359 22049 17368 22083
rect 17316 22040 17368 22049
rect 15936 21972 15988 22024
rect 17592 22040 17644 22092
rect 15568 21904 15620 21956
rect 16488 21904 16540 21956
rect 14280 21836 14332 21888
rect 17132 21836 17184 21888
rect 18972 22108 19024 22160
rect 20444 22176 20496 22228
rect 23480 22176 23532 22228
rect 24676 22176 24728 22228
rect 25136 22219 25188 22228
rect 25136 22185 25145 22219
rect 25145 22185 25179 22219
rect 25179 22185 25188 22219
rect 25136 22176 25188 22185
rect 25320 22219 25372 22228
rect 25320 22185 25329 22219
rect 25329 22185 25363 22219
rect 25363 22185 25372 22219
rect 25320 22176 25372 22185
rect 18420 22083 18472 22092
rect 18420 22049 18429 22083
rect 18429 22049 18463 22083
rect 18463 22049 18472 22083
rect 18420 22040 18472 22049
rect 18880 22040 18932 22092
rect 19064 22083 19116 22092
rect 19064 22049 19098 22083
rect 19098 22049 19116 22083
rect 19064 22040 19116 22049
rect 21548 22151 21600 22160
rect 20168 22040 20220 22092
rect 20444 22083 20496 22092
rect 20444 22049 20453 22083
rect 20453 22049 20487 22083
rect 20487 22049 20496 22083
rect 20444 22040 20496 22049
rect 17960 21904 18012 21956
rect 19984 21836 20036 21888
rect 20260 21879 20312 21888
rect 20260 21845 20269 21879
rect 20269 21845 20303 21879
rect 20303 21845 20312 21879
rect 20260 21836 20312 21845
rect 20444 21904 20496 21956
rect 20720 22083 20772 22092
rect 20720 22049 20755 22083
rect 20755 22049 20772 22083
rect 21548 22117 21582 22151
rect 21582 22117 21600 22151
rect 21548 22108 21600 22117
rect 23204 22108 23256 22160
rect 25964 22151 26016 22160
rect 25964 22117 25973 22151
rect 25973 22117 26007 22151
rect 26007 22117 26016 22151
rect 25964 22108 26016 22117
rect 27436 22176 27488 22228
rect 26608 22108 26660 22160
rect 20720 22040 20772 22049
rect 22836 22040 22888 22092
rect 23112 22083 23164 22092
rect 23112 22049 23121 22083
rect 23121 22049 23155 22083
rect 23155 22049 23164 22083
rect 23112 22040 23164 22049
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 24400 22040 24452 22092
rect 25504 22040 25556 22092
rect 26056 22083 26108 22092
rect 26056 22049 26065 22083
rect 26065 22049 26099 22083
rect 26099 22049 26108 22083
rect 26056 22040 26108 22049
rect 26332 22040 26384 22092
rect 27160 22108 27212 22160
rect 27804 22151 27856 22160
rect 27804 22117 27813 22151
rect 27813 22117 27847 22151
rect 27847 22117 27856 22151
rect 28172 22176 28224 22228
rect 27804 22108 27856 22117
rect 26792 22083 26844 22092
rect 26792 22049 26801 22083
rect 26801 22049 26835 22083
rect 26835 22049 26844 22083
rect 26792 22040 26844 22049
rect 26976 22040 27028 22092
rect 27528 22040 27580 22092
rect 27896 22040 27948 22092
rect 27988 22040 28040 22092
rect 28448 22083 28500 22092
rect 28448 22049 28457 22083
rect 28457 22049 28491 22083
rect 28491 22049 28500 22083
rect 28448 22040 28500 22049
rect 28724 22083 28776 22092
rect 28724 22049 28758 22083
rect 28758 22049 28776 22083
rect 28724 22040 28776 22049
rect 26424 21972 26476 22024
rect 27436 22015 27488 22024
rect 27436 21981 27445 22015
rect 27445 21981 27479 22015
rect 27479 21981 27488 22015
rect 27436 21972 27488 21981
rect 22744 21836 22796 21888
rect 22836 21836 22888 21888
rect 25412 21904 25464 21956
rect 24860 21836 24912 21888
rect 25596 21879 25648 21888
rect 25596 21845 25605 21879
rect 25605 21845 25639 21879
rect 25639 21845 25648 21879
rect 25596 21836 25648 21845
rect 26700 21904 26752 21956
rect 26424 21836 26476 21888
rect 28080 21836 28132 21888
rect 28356 21836 28408 21888
rect 28448 21836 28500 21888
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 11436 21734 11488 21786
rect 11500 21734 11552 21786
rect 11564 21734 11616 21786
rect 11628 21734 11680 21786
rect 11692 21734 11744 21786
rect 19210 21734 19262 21786
rect 19274 21734 19326 21786
rect 19338 21734 19390 21786
rect 19402 21734 19454 21786
rect 19466 21734 19518 21786
rect 26984 21734 27036 21786
rect 27048 21734 27100 21786
rect 27112 21734 27164 21786
rect 27176 21734 27228 21786
rect 27240 21734 27292 21786
rect 13636 21632 13688 21684
rect 14556 21632 14608 21684
rect 14372 21496 14424 21548
rect 14096 21428 14148 21480
rect 15384 21496 15436 21548
rect 17776 21632 17828 21684
rect 19064 21632 19116 21684
rect 20076 21632 20128 21684
rect 20444 21675 20496 21684
rect 20444 21641 20453 21675
rect 20453 21641 20487 21675
rect 20487 21641 20496 21675
rect 20444 21632 20496 21641
rect 21272 21632 21324 21684
rect 20260 21564 20312 21616
rect 14648 21428 14700 21480
rect 17132 21471 17184 21480
rect 17132 21437 17166 21471
rect 17166 21437 17184 21471
rect 17132 21428 17184 21437
rect 15660 21360 15712 21412
rect 20812 21428 20864 21480
rect 22100 21632 22152 21684
rect 23020 21632 23072 21684
rect 23204 21675 23256 21684
rect 23204 21641 23213 21675
rect 23213 21641 23247 21675
rect 23247 21641 23256 21675
rect 23204 21632 23256 21641
rect 24216 21632 24268 21684
rect 25688 21632 25740 21684
rect 27252 21632 27304 21684
rect 27620 21632 27672 21684
rect 28724 21675 28776 21684
rect 28724 21641 28733 21675
rect 28733 21641 28767 21675
rect 28767 21641 28776 21675
rect 28724 21632 28776 21641
rect 23572 21539 23624 21548
rect 23572 21505 23581 21539
rect 23581 21505 23615 21539
rect 23615 21505 23624 21539
rect 23572 21496 23624 21505
rect 24584 21539 24636 21548
rect 24584 21505 24593 21539
rect 24593 21505 24627 21539
rect 24627 21505 24636 21539
rect 24584 21496 24636 21505
rect 24768 21496 24820 21548
rect 25504 21564 25556 21616
rect 21732 21471 21784 21480
rect 21732 21437 21741 21471
rect 21741 21437 21775 21471
rect 21775 21437 21784 21471
rect 21732 21428 21784 21437
rect 22284 21428 22336 21480
rect 23204 21428 23256 21480
rect 19984 21403 20036 21412
rect 19984 21369 19993 21403
rect 19993 21369 20027 21403
rect 20027 21369 20036 21403
rect 19984 21360 20036 21369
rect 16120 21292 16172 21344
rect 18420 21292 18472 21344
rect 18696 21335 18748 21344
rect 18696 21301 18705 21335
rect 18705 21301 18739 21335
rect 18739 21301 18748 21335
rect 18696 21292 18748 21301
rect 19800 21292 19852 21344
rect 20168 21292 20220 21344
rect 20628 21292 20680 21344
rect 21640 21360 21692 21412
rect 24952 21471 25004 21480
rect 24952 21437 24961 21471
rect 24961 21437 24995 21471
rect 24995 21437 25004 21471
rect 24952 21428 25004 21437
rect 25136 21428 25188 21480
rect 25504 21428 25556 21480
rect 25688 21539 25740 21548
rect 25688 21505 25697 21539
rect 25697 21505 25731 21539
rect 25731 21505 25740 21539
rect 25688 21496 25740 21505
rect 25964 21564 26016 21616
rect 26424 21607 26476 21616
rect 26424 21573 26433 21607
rect 26433 21573 26467 21607
rect 26467 21573 26476 21607
rect 26424 21564 26476 21573
rect 28172 21564 28224 21616
rect 28448 21564 28500 21616
rect 24676 21360 24728 21412
rect 25320 21360 25372 21412
rect 26516 21471 26568 21480
rect 26516 21437 26525 21471
rect 26525 21437 26559 21471
rect 26559 21437 26568 21471
rect 26516 21428 26568 21437
rect 26792 21428 26844 21480
rect 27804 21471 27856 21480
rect 27804 21437 27813 21471
rect 27813 21437 27847 21471
rect 27847 21437 27856 21471
rect 27804 21428 27856 21437
rect 27988 21360 28040 21412
rect 28356 21471 28408 21480
rect 28356 21437 28365 21471
rect 28365 21437 28399 21471
rect 28399 21437 28408 21471
rect 28356 21428 28408 21437
rect 29000 21471 29052 21480
rect 29000 21437 29009 21471
rect 29009 21437 29043 21471
rect 29043 21437 29052 21471
rect 29000 21428 29052 21437
rect 28540 21360 28592 21412
rect 22376 21292 22428 21344
rect 23572 21292 23624 21344
rect 23756 21292 23808 21344
rect 25688 21292 25740 21344
rect 25872 21292 25924 21344
rect 26148 21335 26200 21344
rect 26148 21301 26157 21335
rect 26157 21301 26191 21335
rect 26191 21301 26200 21335
rect 26148 21292 26200 21301
rect 28080 21292 28132 21344
rect 28816 21292 28868 21344
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 12096 21190 12148 21242
rect 12160 21190 12212 21242
rect 12224 21190 12276 21242
rect 12288 21190 12340 21242
rect 12352 21190 12404 21242
rect 19870 21190 19922 21242
rect 19934 21190 19986 21242
rect 19998 21190 20050 21242
rect 20062 21190 20114 21242
rect 20126 21190 20178 21242
rect 27644 21190 27696 21242
rect 27708 21190 27760 21242
rect 27772 21190 27824 21242
rect 27836 21190 27888 21242
rect 27900 21190 27952 21242
rect 17592 21131 17644 21140
rect 17592 21097 17601 21131
rect 17601 21097 17635 21131
rect 17635 21097 17644 21131
rect 17592 21088 17644 21097
rect 21732 21088 21784 21140
rect 22744 21088 22796 21140
rect 23940 21088 23992 21140
rect 25136 21131 25188 21140
rect 25136 21097 25145 21131
rect 25145 21097 25179 21131
rect 25179 21097 25188 21131
rect 25136 21088 25188 21097
rect 25412 21088 25464 21140
rect 26332 21088 26384 21140
rect 27252 21088 27304 21140
rect 27712 21131 27764 21140
rect 27712 21097 27721 21131
rect 27721 21097 27755 21131
rect 27755 21097 27764 21131
rect 27712 21088 27764 21097
rect 27988 21131 28040 21140
rect 27988 21097 27997 21131
rect 27997 21097 28031 21131
rect 28031 21097 28040 21131
rect 27988 21088 28040 21097
rect 18696 21020 18748 21072
rect 15384 20952 15436 21004
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 15568 20995 15620 21004
rect 15568 20961 15577 20995
rect 15577 20961 15611 20995
rect 15611 20961 15620 20995
rect 15568 20952 15620 20961
rect 15660 20995 15712 21004
rect 15660 20961 15669 20995
rect 15669 20961 15703 20995
rect 15703 20961 15712 20995
rect 15660 20952 15712 20961
rect 16120 20995 16172 21004
rect 16120 20961 16129 20995
rect 16129 20961 16163 20995
rect 16163 20961 16172 20995
rect 16120 20952 16172 20961
rect 17592 20952 17644 21004
rect 17960 20995 18012 21004
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 22100 20952 22152 21004
rect 27344 20952 27396 21004
rect 18604 20884 18656 20936
rect 24860 20927 24912 20936
rect 24860 20893 24869 20927
rect 24869 20893 24903 20927
rect 24903 20893 24912 20927
rect 24860 20884 24912 20893
rect 27804 20995 27856 21004
rect 27804 20961 27813 20995
rect 27813 20961 27847 20995
rect 27847 20961 27856 20995
rect 27804 20952 27856 20961
rect 28080 20995 28132 21004
rect 28080 20961 28089 20995
rect 28089 20961 28123 20995
rect 28123 20961 28132 20995
rect 28080 20952 28132 20961
rect 27988 20884 28040 20936
rect 17500 20791 17552 20800
rect 17500 20757 17509 20791
rect 17509 20757 17543 20791
rect 17543 20757 17552 20791
rect 17500 20748 17552 20757
rect 23940 20748 23992 20800
rect 24584 20748 24636 20800
rect 28816 20995 28868 21004
rect 28816 20961 28825 20995
rect 28825 20961 28859 20995
rect 28859 20961 28868 20995
rect 28816 20952 28868 20961
rect 28448 20816 28500 20868
rect 28632 20748 28684 20800
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 11436 20646 11488 20698
rect 11500 20646 11552 20698
rect 11564 20646 11616 20698
rect 11628 20646 11680 20698
rect 11692 20646 11744 20698
rect 19210 20646 19262 20698
rect 19274 20646 19326 20698
rect 19338 20646 19390 20698
rect 19402 20646 19454 20698
rect 19466 20646 19518 20698
rect 26984 20646 27036 20698
rect 27048 20646 27100 20698
rect 27112 20646 27164 20698
rect 27176 20646 27228 20698
rect 27240 20646 27292 20698
rect 15476 20544 15528 20596
rect 18236 20476 18288 20528
rect 16672 20340 16724 20392
rect 17500 20340 17552 20392
rect 17592 20340 17644 20392
rect 18880 20340 18932 20392
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 20260 20408 20312 20460
rect 20628 20408 20680 20460
rect 25596 20544 25648 20596
rect 25780 20544 25832 20596
rect 28080 20544 28132 20596
rect 24952 20476 25004 20528
rect 27804 20476 27856 20528
rect 28724 20476 28776 20528
rect 20812 20340 20864 20392
rect 21640 20340 21692 20392
rect 22008 20383 22060 20392
rect 22008 20349 22017 20383
rect 22017 20349 22051 20383
rect 22051 20349 22060 20383
rect 22008 20340 22060 20349
rect 16580 20272 16632 20324
rect 18052 20204 18104 20256
rect 18328 20247 18380 20256
rect 18328 20213 18337 20247
rect 18337 20213 18371 20247
rect 18371 20213 18380 20247
rect 18328 20204 18380 20213
rect 19156 20204 19208 20256
rect 19708 20247 19760 20256
rect 19708 20213 19717 20247
rect 19717 20213 19751 20247
rect 19751 20213 19760 20247
rect 19708 20204 19760 20213
rect 20720 20272 20772 20324
rect 21732 20272 21784 20324
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 23296 20408 23348 20460
rect 23480 20340 23532 20392
rect 24032 20340 24084 20392
rect 23940 20272 23992 20324
rect 20536 20204 20588 20256
rect 22100 20247 22152 20256
rect 22100 20213 22109 20247
rect 22109 20213 22143 20247
rect 22143 20213 22152 20247
rect 22100 20204 22152 20213
rect 22192 20204 22244 20256
rect 22560 20204 22612 20256
rect 24216 20340 24268 20392
rect 26608 20408 26660 20460
rect 25504 20383 25556 20392
rect 25504 20349 25518 20383
rect 25518 20349 25552 20383
rect 25552 20349 25556 20383
rect 25504 20340 25556 20349
rect 27988 20340 28040 20392
rect 28356 20340 28408 20392
rect 25688 20272 25740 20324
rect 25872 20272 25924 20324
rect 27436 20272 27488 20324
rect 26056 20204 26108 20256
rect 27712 20204 27764 20256
rect 28080 20204 28132 20256
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 12096 20102 12148 20154
rect 12160 20102 12212 20154
rect 12224 20102 12276 20154
rect 12288 20102 12340 20154
rect 12352 20102 12404 20154
rect 19870 20102 19922 20154
rect 19934 20102 19986 20154
rect 19998 20102 20050 20154
rect 20062 20102 20114 20154
rect 20126 20102 20178 20154
rect 27644 20102 27696 20154
rect 27708 20102 27760 20154
rect 27772 20102 27824 20154
rect 27836 20102 27888 20154
rect 27900 20102 27952 20154
rect 14832 20000 14884 20052
rect 18236 20000 18288 20052
rect 18512 20000 18564 20052
rect 19248 20000 19300 20052
rect 22100 20000 22152 20052
rect 14832 19907 14884 19916
rect 14832 19873 14841 19907
rect 14841 19873 14875 19907
rect 14875 19873 14884 19907
rect 14832 19864 14884 19873
rect 16488 19932 16540 19984
rect 15384 19864 15436 19916
rect 18328 19932 18380 19984
rect 19616 19932 19668 19984
rect 20260 19932 20312 19984
rect 17960 19907 18012 19916
rect 17960 19873 17994 19907
rect 17994 19873 18012 19907
rect 17960 19864 18012 19873
rect 19156 19907 19208 19916
rect 19156 19873 19165 19907
rect 19165 19873 19199 19907
rect 19199 19873 19208 19907
rect 19156 19864 19208 19873
rect 22008 19932 22060 19984
rect 23388 19932 23440 19984
rect 25320 19932 25372 19984
rect 26240 20000 26292 20052
rect 21640 19907 21692 19916
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 21732 19907 21784 19916
rect 21732 19873 21767 19907
rect 21767 19873 21784 19907
rect 21732 19864 21784 19873
rect 15844 19796 15896 19848
rect 14648 19660 14700 19712
rect 19800 19660 19852 19712
rect 21088 19796 21140 19848
rect 23664 19864 23716 19916
rect 24124 19864 24176 19916
rect 24308 19864 24360 19916
rect 24952 19907 25004 19916
rect 24952 19873 24961 19907
rect 24961 19873 24995 19907
rect 24995 19873 25004 19907
rect 24952 19864 25004 19873
rect 22284 19839 22336 19848
rect 22284 19805 22293 19839
rect 22293 19805 22327 19839
rect 22327 19805 22336 19839
rect 22284 19796 22336 19805
rect 23756 19839 23808 19848
rect 23756 19805 23765 19839
rect 23765 19805 23799 19839
rect 23799 19805 23808 19839
rect 23756 19796 23808 19805
rect 24216 19839 24268 19848
rect 24216 19805 24225 19839
rect 24225 19805 24259 19839
rect 24259 19805 24268 19839
rect 24216 19796 24268 19805
rect 20536 19771 20588 19780
rect 20536 19737 20545 19771
rect 20545 19737 20579 19771
rect 20579 19737 20588 19771
rect 25780 19907 25832 19916
rect 25780 19873 25789 19907
rect 25789 19873 25823 19907
rect 25823 19873 25832 19907
rect 25780 19864 25832 19873
rect 25688 19796 25740 19848
rect 26608 19907 26660 19916
rect 26608 19873 26617 19907
rect 26617 19873 26651 19907
rect 26651 19873 26660 19907
rect 26608 19864 26660 19873
rect 28908 19932 28960 19984
rect 28172 19864 28224 19916
rect 26240 19839 26292 19848
rect 26240 19805 26249 19839
rect 26249 19805 26283 19839
rect 26283 19805 26292 19839
rect 26240 19796 26292 19805
rect 20536 19728 20588 19737
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 25872 19660 25924 19712
rect 26056 19660 26108 19712
rect 27436 19796 27488 19848
rect 26700 19660 26752 19712
rect 27344 19660 27396 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 11436 19558 11488 19610
rect 11500 19558 11552 19610
rect 11564 19558 11616 19610
rect 11628 19558 11680 19610
rect 11692 19558 11744 19610
rect 19210 19558 19262 19610
rect 19274 19558 19326 19610
rect 19338 19558 19390 19610
rect 19402 19558 19454 19610
rect 19466 19558 19518 19610
rect 26984 19558 27036 19610
rect 27048 19558 27100 19610
rect 27112 19558 27164 19610
rect 27176 19558 27228 19610
rect 27240 19558 27292 19610
rect 19616 19456 19668 19508
rect 13820 19252 13872 19304
rect 14648 19295 14700 19304
rect 14648 19261 14682 19295
rect 14682 19261 14700 19295
rect 14648 19252 14700 19261
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 16580 19388 16632 19440
rect 17408 19388 17460 19440
rect 21088 19456 21140 19508
rect 22008 19456 22060 19508
rect 22560 19456 22612 19508
rect 26516 19456 26568 19508
rect 28080 19456 28132 19508
rect 15200 19184 15252 19236
rect 16488 19252 16540 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 25228 19431 25280 19440
rect 25228 19397 25237 19431
rect 25237 19397 25271 19431
rect 25271 19397 25280 19431
rect 25228 19388 25280 19397
rect 27436 19388 27488 19440
rect 15660 19116 15712 19168
rect 17776 19184 17828 19236
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 19708 19320 19760 19372
rect 16488 19159 16540 19168
rect 16488 19125 16497 19159
rect 16497 19125 16531 19159
rect 16531 19125 16540 19159
rect 16488 19116 16540 19125
rect 16580 19116 16632 19168
rect 17960 19116 18012 19168
rect 18236 19116 18288 19168
rect 19800 19252 19852 19304
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 26700 19363 26752 19372
rect 26700 19329 26709 19363
rect 26709 19329 26743 19363
rect 26743 19329 26752 19363
rect 26700 19320 26752 19329
rect 21456 19252 21508 19304
rect 21548 19252 21600 19304
rect 23572 19252 23624 19304
rect 24400 19252 24452 19304
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 26332 19295 26384 19304
rect 26332 19261 26341 19295
rect 26341 19261 26375 19295
rect 26375 19261 26384 19295
rect 26332 19252 26384 19261
rect 26976 19295 27028 19304
rect 26976 19261 26985 19295
rect 26985 19261 27019 19295
rect 27019 19261 27028 19295
rect 26976 19252 27028 19261
rect 27344 19252 27396 19304
rect 27988 19252 28040 19304
rect 20628 19227 20680 19236
rect 20628 19193 20662 19227
rect 20662 19193 20680 19227
rect 20628 19184 20680 19193
rect 22100 19227 22152 19236
rect 22100 19193 22134 19227
rect 22134 19193 22152 19227
rect 22100 19184 22152 19193
rect 24492 19184 24544 19236
rect 26148 19184 26200 19236
rect 28540 19252 28592 19304
rect 22376 19116 22428 19168
rect 23296 19116 23348 19168
rect 28264 19227 28316 19236
rect 28264 19193 28289 19227
rect 28289 19193 28316 19227
rect 28264 19184 28316 19193
rect 28448 19159 28500 19168
rect 28448 19125 28457 19159
rect 28457 19125 28491 19159
rect 28491 19125 28500 19159
rect 28448 19116 28500 19125
rect 28632 19116 28684 19168
rect 29368 19116 29420 19168
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 12096 19014 12148 19066
rect 12160 19014 12212 19066
rect 12224 19014 12276 19066
rect 12288 19014 12340 19066
rect 12352 19014 12404 19066
rect 19870 19014 19922 19066
rect 19934 19014 19986 19066
rect 19998 19014 20050 19066
rect 20062 19014 20114 19066
rect 20126 19014 20178 19066
rect 27644 19014 27696 19066
rect 27708 19014 27760 19066
rect 27772 19014 27824 19066
rect 27836 19014 27888 19066
rect 27900 19014 27952 19066
rect 16488 18912 16540 18964
rect 16856 18912 16908 18964
rect 21272 18912 21324 18964
rect 21548 18955 21600 18964
rect 21548 18921 21557 18955
rect 21557 18921 21591 18955
rect 21591 18921 21600 18955
rect 21548 18912 21600 18921
rect 22100 18955 22152 18964
rect 22100 18921 22109 18955
rect 22109 18921 22143 18955
rect 22143 18921 22152 18955
rect 22100 18912 22152 18921
rect 23572 18955 23624 18964
rect 23572 18921 23581 18955
rect 23581 18921 23615 18955
rect 23615 18921 23624 18955
rect 23572 18912 23624 18921
rect 17868 18844 17920 18896
rect 22284 18844 22336 18896
rect 15200 18776 15252 18828
rect 16304 18776 16356 18828
rect 16580 18776 16632 18828
rect 21548 18776 21600 18828
rect 22192 18776 22244 18828
rect 23020 18776 23072 18828
rect 23664 18776 23716 18828
rect 23940 18912 23992 18964
rect 24400 18955 24452 18964
rect 24400 18921 24409 18955
rect 24409 18921 24443 18955
rect 24443 18921 24452 18955
rect 24400 18912 24452 18921
rect 26056 18912 26108 18964
rect 25228 18844 25280 18896
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 23296 18708 23348 18760
rect 17776 18640 17828 18692
rect 19800 18640 19852 18692
rect 21640 18640 21692 18692
rect 24032 18819 24084 18828
rect 24032 18785 24067 18819
rect 24067 18785 24084 18819
rect 24032 18776 24084 18785
rect 24492 18819 24544 18828
rect 24492 18785 24501 18819
rect 24501 18785 24535 18819
rect 24535 18785 24544 18819
rect 24492 18776 24544 18785
rect 25136 18776 25188 18828
rect 26884 18776 26936 18828
rect 28540 18844 28592 18896
rect 24768 18708 24820 18760
rect 26516 18751 26568 18760
rect 26516 18717 26525 18751
rect 26525 18717 26559 18751
rect 26559 18717 26568 18751
rect 26516 18708 26568 18717
rect 26976 18751 27028 18760
rect 26976 18717 26985 18751
rect 26985 18717 27019 18751
rect 27019 18717 27028 18751
rect 26976 18708 27028 18717
rect 27436 18751 27488 18760
rect 27436 18717 27445 18751
rect 27445 18717 27479 18751
rect 27479 18717 27488 18751
rect 27436 18708 27488 18717
rect 15844 18572 15896 18624
rect 17500 18572 17552 18624
rect 19616 18572 19668 18624
rect 23940 18640 23992 18692
rect 24032 18572 24084 18624
rect 24860 18572 24912 18624
rect 27436 18572 27488 18624
rect 28448 18776 28500 18828
rect 29368 18887 29420 18896
rect 29368 18853 29377 18887
rect 29377 18853 29411 18887
rect 29411 18853 29420 18887
rect 29368 18844 29420 18853
rect 30380 18776 30432 18828
rect 28080 18708 28132 18760
rect 28264 18708 28316 18760
rect 28724 18640 28776 18692
rect 28632 18572 28684 18624
rect 29552 18615 29604 18624
rect 29552 18581 29561 18615
rect 29561 18581 29595 18615
rect 29595 18581 29604 18615
rect 29552 18572 29604 18581
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 11436 18470 11488 18522
rect 11500 18470 11552 18522
rect 11564 18470 11616 18522
rect 11628 18470 11680 18522
rect 11692 18470 11744 18522
rect 19210 18470 19262 18522
rect 19274 18470 19326 18522
rect 19338 18470 19390 18522
rect 19402 18470 19454 18522
rect 19466 18470 19518 18522
rect 26984 18470 27036 18522
rect 27048 18470 27100 18522
rect 27112 18470 27164 18522
rect 27176 18470 27228 18522
rect 27240 18470 27292 18522
rect 16304 18368 16356 18420
rect 26056 18368 26108 18420
rect 27988 18368 28040 18420
rect 30380 18411 30432 18420
rect 30380 18377 30389 18411
rect 30389 18377 30423 18411
rect 30423 18377 30432 18411
rect 30380 18368 30432 18377
rect 13820 18164 13872 18216
rect 17868 18164 17920 18216
rect 18972 18232 19024 18284
rect 20260 18232 20312 18284
rect 18236 18207 18288 18216
rect 18236 18173 18245 18207
rect 18245 18173 18279 18207
rect 18279 18173 18288 18207
rect 18236 18164 18288 18173
rect 18328 18207 18380 18216
rect 18328 18173 18337 18207
rect 18337 18173 18371 18207
rect 18371 18173 18380 18207
rect 18328 18164 18380 18173
rect 14832 18071 14884 18080
rect 14832 18037 14841 18071
rect 14841 18037 14875 18071
rect 14875 18037 14884 18071
rect 14832 18028 14884 18037
rect 15200 18139 15252 18148
rect 15200 18105 15209 18139
rect 15209 18105 15243 18139
rect 15243 18105 15252 18139
rect 15200 18096 15252 18105
rect 15476 18096 15528 18148
rect 16580 18096 16632 18148
rect 17224 18096 17276 18148
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 20536 18232 20588 18284
rect 20628 18232 20680 18284
rect 20720 18232 20772 18284
rect 21824 18232 21876 18284
rect 22008 18232 22060 18284
rect 15292 18028 15344 18080
rect 16396 18028 16448 18080
rect 19800 18096 19852 18148
rect 21640 18164 21692 18216
rect 24492 18164 24544 18216
rect 18052 18028 18104 18080
rect 19708 18028 19760 18080
rect 21732 18096 21784 18148
rect 20812 18028 20864 18080
rect 27436 18164 27488 18216
rect 29000 18207 29052 18216
rect 29000 18173 29009 18207
rect 29009 18173 29043 18207
rect 29043 18173 29052 18207
rect 29000 18164 29052 18173
rect 29552 18164 29604 18216
rect 27988 18028 28040 18080
rect 28724 18071 28776 18080
rect 28724 18037 28733 18071
rect 28733 18037 28767 18071
rect 28767 18037 28776 18071
rect 28724 18028 28776 18037
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 12096 17926 12148 17978
rect 12160 17926 12212 17978
rect 12224 17926 12276 17978
rect 12288 17926 12340 17978
rect 12352 17926 12404 17978
rect 19870 17926 19922 17978
rect 19934 17926 19986 17978
rect 19998 17926 20050 17978
rect 20062 17926 20114 17978
rect 20126 17926 20178 17978
rect 27644 17926 27696 17978
rect 27708 17926 27760 17978
rect 27772 17926 27824 17978
rect 27836 17926 27888 17978
rect 27900 17926 27952 17978
rect 15292 17824 15344 17876
rect 16948 17824 17000 17876
rect 19616 17824 19668 17876
rect 20812 17824 20864 17876
rect 13912 17688 13964 17740
rect 15752 17756 15804 17808
rect 16396 17756 16448 17808
rect 17500 17799 17552 17808
rect 17500 17765 17509 17799
rect 17509 17765 17543 17799
rect 17543 17765 17552 17799
rect 17500 17756 17552 17765
rect 17868 17756 17920 17808
rect 21916 17824 21968 17876
rect 26516 17824 26568 17876
rect 29000 17824 29052 17876
rect 14832 17731 14884 17740
rect 14832 17697 14841 17731
rect 14841 17697 14875 17731
rect 14875 17697 14884 17731
rect 14832 17688 14884 17697
rect 15384 17688 15436 17740
rect 16028 17688 16080 17740
rect 16580 17731 16632 17740
rect 16580 17697 16589 17731
rect 16589 17697 16623 17731
rect 16623 17697 16632 17731
rect 16580 17688 16632 17697
rect 17592 17688 17644 17740
rect 18052 17731 18104 17740
rect 18052 17697 18086 17731
rect 18086 17697 18104 17731
rect 18052 17688 18104 17697
rect 21640 17799 21692 17808
rect 21640 17765 21649 17799
rect 21649 17765 21683 17799
rect 21683 17765 21692 17799
rect 21640 17756 21692 17765
rect 23756 17756 23808 17808
rect 25780 17756 25832 17808
rect 19616 17731 19668 17740
rect 19616 17697 19650 17731
rect 19650 17697 19668 17731
rect 19616 17688 19668 17697
rect 20536 17688 20588 17740
rect 21364 17688 21416 17740
rect 21732 17731 21784 17740
rect 21732 17697 21767 17731
rect 21767 17697 21784 17731
rect 21732 17688 21784 17697
rect 22008 17688 22060 17740
rect 15292 17620 15344 17672
rect 17776 17663 17828 17672
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 21272 17620 21324 17672
rect 22100 17620 22152 17672
rect 23020 17688 23072 17740
rect 23112 17731 23164 17740
rect 23112 17697 23121 17731
rect 23121 17697 23155 17731
rect 23155 17697 23164 17731
rect 23112 17688 23164 17697
rect 22560 17620 22612 17672
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 24492 17731 24544 17740
rect 24492 17697 24501 17731
rect 24501 17697 24535 17731
rect 24535 17697 24544 17731
rect 24492 17688 24544 17697
rect 24676 17731 24728 17740
rect 24676 17697 24685 17731
rect 24685 17697 24719 17731
rect 24719 17697 24728 17731
rect 24676 17688 24728 17697
rect 24400 17620 24452 17672
rect 24768 17620 24820 17672
rect 23020 17552 23072 17604
rect 25688 17688 25740 17740
rect 26056 17731 26108 17740
rect 26056 17697 26065 17731
rect 26065 17697 26099 17731
rect 26099 17697 26108 17731
rect 26056 17688 26108 17697
rect 27988 17688 28040 17740
rect 28724 17620 28776 17672
rect 25504 17552 25556 17604
rect 14188 17484 14240 17536
rect 19064 17484 19116 17536
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 21824 17484 21876 17536
rect 22928 17527 22980 17536
rect 22928 17493 22937 17527
rect 22937 17493 22971 17527
rect 22971 17493 22980 17527
rect 22928 17484 22980 17493
rect 24216 17484 24268 17536
rect 26240 17484 26292 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 11436 17382 11488 17434
rect 11500 17382 11552 17434
rect 11564 17382 11616 17434
rect 11628 17382 11680 17434
rect 11692 17382 11744 17434
rect 19210 17382 19262 17434
rect 19274 17382 19326 17434
rect 19338 17382 19390 17434
rect 19402 17382 19454 17434
rect 19466 17382 19518 17434
rect 26984 17382 27036 17434
rect 27048 17382 27100 17434
rect 27112 17382 27164 17434
rect 27176 17382 27228 17434
rect 27240 17382 27292 17434
rect 15292 17323 15344 17332
rect 15292 17289 15301 17323
rect 15301 17289 15335 17323
rect 15335 17289 15344 17323
rect 15292 17280 15344 17289
rect 15476 17280 15528 17332
rect 17776 17280 17828 17332
rect 19616 17280 19668 17332
rect 18328 17212 18380 17264
rect 20720 17280 20772 17332
rect 21916 17280 21968 17332
rect 22836 17280 22888 17332
rect 24676 17280 24728 17332
rect 26332 17280 26384 17332
rect 26608 17280 26660 17332
rect 24032 17212 24084 17264
rect 24308 17212 24360 17264
rect 13636 17119 13688 17128
rect 13636 17085 13645 17119
rect 13645 17085 13679 17119
rect 13679 17085 13688 17119
rect 13636 17076 13688 17085
rect 14188 17119 14240 17128
rect 14188 17085 14222 17119
rect 14222 17085 14240 17119
rect 14188 17076 14240 17085
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 15844 17119 15896 17128
rect 15844 17085 15853 17119
rect 15853 17085 15887 17119
rect 15887 17085 15896 17119
rect 15844 17076 15896 17085
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 17592 17076 17644 17128
rect 18880 17076 18932 17128
rect 19708 17076 19760 17128
rect 19800 17119 19852 17128
rect 19800 17085 19809 17119
rect 19809 17085 19843 17119
rect 19843 17085 19852 17119
rect 19800 17076 19852 17085
rect 21548 17076 21600 17128
rect 22928 17076 22980 17128
rect 23664 17076 23716 17128
rect 24584 17187 24636 17196
rect 24584 17153 24593 17187
rect 24593 17153 24627 17187
rect 24627 17153 24636 17187
rect 24584 17144 24636 17153
rect 24400 17076 24452 17128
rect 24860 17119 24912 17128
rect 24860 17085 24869 17119
rect 24869 17085 24903 17119
rect 24903 17085 24912 17119
rect 24860 17076 24912 17085
rect 25596 17144 25648 17196
rect 25044 17119 25096 17128
rect 25044 17085 25053 17119
rect 25053 17085 25087 17119
rect 25087 17085 25096 17119
rect 25044 17076 25096 17085
rect 25504 17119 25556 17128
rect 25504 17085 25513 17119
rect 25513 17085 25547 17119
rect 25547 17085 25556 17119
rect 25504 17076 25556 17085
rect 19064 17008 19116 17060
rect 19616 16940 19668 16992
rect 20536 17008 20588 17060
rect 24768 17051 24820 17060
rect 24768 17017 24785 17051
rect 24785 17017 24820 17051
rect 23664 16940 23716 16992
rect 24768 17008 24820 17017
rect 25964 17076 26016 17128
rect 26240 17076 26292 17128
rect 26424 17119 26476 17128
rect 26424 17085 26434 17119
rect 26434 17085 26468 17119
rect 26468 17085 26476 17119
rect 26424 17076 26476 17085
rect 27528 17280 27580 17332
rect 27252 17119 27304 17128
rect 27252 17085 27261 17119
rect 27261 17085 27295 17119
rect 27295 17085 27304 17119
rect 27252 17076 27304 17085
rect 25136 16940 25188 16992
rect 25872 16940 25924 16992
rect 25964 16940 26016 16992
rect 26424 16940 26476 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 12096 16838 12148 16890
rect 12160 16838 12212 16890
rect 12224 16838 12276 16890
rect 12288 16838 12340 16890
rect 12352 16838 12404 16890
rect 19870 16838 19922 16890
rect 19934 16838 19986 16890
rect 19998 16838 20050 16890
rect 20062 16838 20114 16890
rect 20126 16838 20178 16890
rect 27644 16838 27696 16890
rect 27708 16838 27760 16890
rect 27772 16838 27824 16890
rect 27836 16838 27888 16890
rect 27900 16838 27952 16890
rect 18328 16736 18380 16788
rect 20536 16779 20588 16788
rect 20536 16745 20545 16779
rect 20545 16745 20579 16779
rect 20579 16745 20588 16779
rect 20536 16736 20588 16745
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15476 16643 15528 16652
rect 15476 16609 15489 16643
rect 15489 16609 15528 16643
rect 15476 16600 15528 16609
rect 15660 16600 15712 16652
rect 16672 16668 16724 16720
rect 17040 16668 17092 16720
rect 18236 16668 18288 16720
rect 23020 16736 23072 16788
rect 23112 16779 23164 16788
rect 23112 16745 23121 16779
rect 23121 16745 23155 16779
rect 23155 16745 23164 16779
rect 23112 16736 23164 16745
rect 23480 16736 23532 16788
rect 25044 16736 25096 16788
rect 25596 16779 25648 16788
rect 25596 16745 25605 16779
rect 25605 16745 25639 16779
rect 25639 16745 25648 16779
rect 25596 16736 25648 16745
rect 27252 16736 27304 16788
rect 16488 16643 16540 16652
rect 16488 16609 16497 16643
rect 16497 16609 16531 16643
rect 16531 16609 16540 16643
rect 16488 16600 16540 16609
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 17408 16643 17460 16652
rect 17408 16609 17417 16643
rect 17417 16609 17451 16643
rect 17451 16609 17460 16643
rect 17408 16600 17460 16609
rect 18512 16643 18564 16652
rect 18512 16609 18521 16643
rect 18521 16609 18555 16643
rect 18555 16609 18564 16643
rect 18512 16600 18564 16609
rect 21640 16711 21692 16720
rect 21640 16677 21649 16711
rect 21649 16677 21683 16711
rect 21683 16677 21692 16711
rect 21640 16668 21692 16677
rect 21732 16668 21784 16720
rect 22560 16668 22612 16720
rect 22836 16711 22888 16720
rect 22836 16677 22845 16711
rect 22845 16677 22879 16711
rect 22879 16677 22888 16711
rect 22836 16668 22888 16677
rect 23296 16668 23348 16720
rect 18880 16600 18932 16652
rect 19708 16600 19760 16652
rect 21272 16600 21324 16652
rect 21364 16600 21416 16652
rect 16120 16464 16172 16516
rect 19616 16532 19668 16584
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 23480 16600 23532 16652
rect 23664 16643 23716 16652
rect 23664 16609 23673 16643
rect 23673 16609 23707 16643
rect 23707 16609 23716 16643
rect 23664 16600 23716 16609
rect 24216 16643 24268 16652
rect 24216 16609 24225 16643
rect 24225 16609 24259 16643
rect 24259 16609 24268 16643
rect 24216 16600 24268 16609
rect 25872 16643 25924 16652
rect 25872 16609 25881 16643
rect 25881 16609 25915 16643
rect 25915 16609 25924 16643
rect 25872 16600 25924 16609
rect 26792 16668 26844 16720
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 27344 16600 27396 16652
rect 27436 16643 27488 16652
rect 27436 16609 27445 16643
rect 27445 16609 27479 16643
rect 27479 16609 27488 16643
rect 27436 16600 27488 16609
rect 27988 16643 28040 16652
rect 27988 16609 27997 16643
rect 27997 16609 28031 16643
rect 28031 16609 28040 16643
rect 27988 16600 28040 16609
rect 29000 16600 29052 16652
rect 18972 16464 19024 16516
rect 15384 16396 15436 16448
rect 16672 16439 16724 16448
rect 16672 16405 16681 16439
rect 16681 16405 16715 16439
rect 16715 16405 16724 16439
rect 16672 16396 16724 16405
rect 16948 16439 17000 16448
rect 16948 16405 16957 16439
rect 16957 16405 16991 16439
rect 16991 16405 17000 16439
rect 16948 16396 17000 16405
rect 17316 16396 17368 16448
rect 17868 16396 17920 16448
rect 18604 16396 18656 16448
rect 20904 16396 20956 16448
rect 23940 16396 23992 16448
rect 26424 16396 26476 16448
rect 27988 16396 28040 16448
rect 28724 16396 28776 16448
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 11436 16294 11488 16346
rect 11500 16294 11552 16346
rect 11564 16294 11616 16346
rect 11628 16294 11680 16346
rect 11692 16294 11744 16346
rect 19210 16294 19262 16346
rect 19274 16294 19326 16346
rect 19338 16294 19390 16346
rect 19402 16294 19454 16346
rect 19466 16294 19518 16346
rect 26984 16294 27036 16346
rect 27048 16294 27100 16346
rect 27112 16294 27164 16346
rect 27176 16294 27228 16346
rect 27240 16294 27292 16346
rect 17132 16192 17184 16244
rect 17408 16235 17460 16244
rect 17408 16201 17417 16235
rect 17417 16201 17451 16235
rect 17451 16201 17460 16235
rect 17408 16192 17460 16201
rect 16948 16124 17000 16176
rect 15384 16031 15436 16040
rect 15384 15997 15393 16031
rect 15393 15997 15427 16031
rect 15427 15997 15436 16031
rect 15384 15988 15436 15997
rect 15660 15988 15712 16040
rect 16672 16056 16724 16108
rect 17776 16192 17828 16244
rect 18328 16192 18380 16244
rect 19524 16235 19576 16244
rect 19524 16201 19533 16235
rect 19533 16201 19567 16235
rect 19567 16201 19576 16235
rect 19524 16192 19576 16201
rect 20352 16192 20404 16244
rect 25136 16192 25188 16244
rect 27436 16192 27488 16244
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16396 15988 16448 16040
rect 16488 15988 16540 16040
rect 17040 16031 17092 16040
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 17316 16031 17368 16040
rect 17316 15997 17325 16031
rect 17325 15997 17359 16031
rect 17359 15997 17368 16031
rect 17316 15988 17368 15997
rect 18512 16124 18564 16176
rect 17776 16056 17828 16108
rect 16212 15963 16264 15972
rect 16212 15929 16221 15963
rect 16221 15929 16255 15963
rect 16255 15929 16264 15963
rect 16212 15920 16264 15929
rect 17592 15852 17644 15904
rect 17960 16031 18012 16040
rect 17960 15997 17969 16031
rect 17969 15997 18003 16031
rect 18003 15997 18012 16031
rect 17960 15988 18012 15997
rect 18144 16031 18196 16040
rect 18144 15997 18154 16031
rect 18154 15997 18188 16031
rect 18188 15997 18196 16031
rect 18144 15988 18196 15997
rect 18604 15988 18656 16040
rect 18972 16031 19024 16040
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 26516 16124 26568 16176
rect 26700 16124 26752 16176
rect 19340 15988 19392 16040
rect 20444 16056 20496 16108
rect 21180 16056 21232 16108
rect 19616 16031 19668 16040
rect 19616 15997 19625 16031
rect 19625 15997 19659 16031
rect 19659 15997 19668 16031
rect 19616 15988 19668 15997
rect 20904 16031 20956 16040
rect 20904 15997 20913 16031
rect 20913 15997 20947 16031
rect 20947 15997 20956 16031
rect 20904 15988 20956 15997
rect 21548 16031 21600 16040
rect 21548 15997 21557 16031
rect 21557 15997 21591 16031
rect 21591 15997 21600 16031
rect 21548 15988 21600 15997
rect 23940 15988 23992 16040
rect 26792 15988 26844 16040
rect 27344 16031 27396 16040
rect 27344 15997 27353 16031
rect 27353 15997 27387 16031
rect 27387 15997 27396 16031
rect 27344 15988 27396 15997
rect 27988 15988 28040 16040
rect 29000 16031 29052 16040
rect 29000 15997 29009 16031
rect 29009 15997 29043 16031
rect 29043 15997 29052 16031
rect 29000 15988 29052 15997
rect 18420 15920 18472 15972
rect 19064 15963 19116 15972
rect 19064 15929 19073 15963
rect 19073 15929 19107 15963
rect 19107 15929 19116 15963
rect 19064 15920 19116 15929
rect 26884 15963 26936 15972
rect 26884 15929 26893 15963
rect 26893 15929 26927 15963
rect 26927 15929 26936 15963
rect 26884 15920 26936 15929
rect 21088 15895 21140 15904
rect 21088 15861 21097 15895
rect 21097 15861 21131 15895
rect 21131 15861 21140 15895
rect 21088 15852 21140 15861
rect 21272 15852 21324 15904
rect 26240 15852 26292 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 12096 15750 12148 15802
rect 12160 15750 12212 15802
rect 12224 15750 12276 15802
rect 12288 15750 12340 15802
rect 12352 15750 12404 15802
rect 19870 15750 19922 15802
rect 19934 15750 19986 15802
rect 19998 15750 20050 15802
rect 20062 15750 20114 15802
rect 20126 15750 20178 15802
rect 27644 15750 27696 15802
rect 27708 15750 27760 15802
rect 27772 15750 27824 15802
rect 27836 15750 27888 15802
rect 27900 15750 27952 15802
rect 15844 15648 15896 15700
rect 16488 15648 16540 15700
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 23020 15648 23072 15700
rect 15476 15580 15528 15632
rect 16856 15512 16908 15564
rect 18052 15512 18104 15564
rect 21088 15580 21140 15632
rect 19708 15512 19760 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 26424 15555 26476 15564
rect 26424 15521 26433 15555
rect 26433 15521 26467 15555
rect 26467 15521 26476 15555
rect 26424 15512 26476 15521
rect 19524 15487 19576 15496
rect 19524 15453 19533 15487
rect 19533 15453 19567 15487
rect 19567 15453 19576 15487
rect 19524 15444 19576 15453
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 27344 15512 27396 15564
rect 28724 15555 28776 15564
rect 28724 15521 28733 15555
rect 28733 15521 28767 15555
rect 28767 15521 28776 15555
rect 28724 15512 28776 15521
rect 27436 15444 27488 15496
rect 15292 15376 15344 15428
rect 19616 15376 19668 15428
rect 19708 15351 19760 15360
rect 19708 15317 19717 15351
rect 19717 15317 19751 15351
rect 19751 15317 19760 15351
rect 19708 15308 19760 15317
rect 26608 15351 26660 15360
rect 26608 15317 26617 15351
rect 26617 15317 26651 15351
rect 26651 15317 26660 15351
rect 26884 15376 26936 15428
rect 26608 15308 26660 15317
rect 26792 15308 26844 15360
rect 27528 15308 27580 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 11436 15206 11488 15258
rect 11500 15206 11552 15258
rect 11564 15206 11616 15258
rect 11628 15206 11680 15258
rect 11692 15206 11744 15258
rect 19210 15206 19262 15258
rect 19274 15206 19326 15258
rect 19338 15206 19390 15258
rect 19402 15206 19454 15258
rect 19466 15206 19518 15258
rect 26984 15206 27036 15258
rect 27048 15206 27100 15258
rect 27112 15206 27164 15258
rect 27176 15206 27228 15258
rect 27240 15206 27292 15258
rect 16948 15147 17000 15156
rect 16948 15113 16957 15147
rect 16957 15113 16991 15147
rect 16991 15113 17000 15147
rect 16948 15104 17000 15113
rect 20904 15104 20956 15156
rect 17224 15036 17276 15088
rect 16488 15011 16540 15020
rect 16488 14977 16497 15011
rect 16497 14977 16531 15011
rect 16531 14977 16540 15011
rect 16488 14968 16540 14977
rect 13636 14900 13688 14952
rect 16120 14900 16172 14952
rect 16212 14900 16264 14952
rect 16672 14943 16724 14952
rect 16672 14909 16681 14943
rect 16681 14909 16715 14943
rect 16715 14909 16724 14943
rect 16672 14900 16724 14909
rect 17776 14900 17828 14952
rect 18236 14900 18288 14952
rect 18328 14900 18380 14952
rect 18972 14943 19024 14952
rect 18972 14909 18981 14943
rect 18981 14909 19015 14943
rect 19015 14909 19024 14943
rect 18972 14900 19024 14909
rect 19616 15011 19668 15020
rect 19616 14977 19625 15011
rect 19625 14977 19659 15011
rect 19659 14977 19668 15011
rect 19616 14968 19668 14977
rect 23296 15104 23348 15156
rect 23756 15104 23808 15156
rect 16580 14832 16632 14884
rect 18144 14875 18196 14884
rect 18144 14841 18153 14875
rect 18153 14841 18187 14875
rect 18187 14841 18196 14875
rect 19708 14900 19760 14952
rect 21824 14943 21876 14952
rect 21824 14909 21833 14943
rect 21833 14909 21867 14943
rect 21867 14909 21876 14943
rect 21824 14900 21876 14909
rect 22100 14943 22152 14952
rect 22100 14909 22109 14943
rect 22109 14909 22143 14943
rect 22143 14909 22152 14943
rect 22100 14900 22152 14909
rect 25044 14900 25096 14952
rect 26608 15104 26660 15156
rect 26700 15104 26752 15156
rect 27344 15104 27396 15156
rect 18144 14832 18196 14841
rect 20904 14832 20956 14884
rect 14188 14764 14240 14816
rect 15384 14764 15436 14816
rect 18328 14764 18380 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 18972 14764 19024 14816
rect 25688 14943 25740 14952
rect 25688 14909 25697 14943
rect 25697 14909 25731 14943
rect 25731 14909 25740 14943
rect 25688 14900 25740 14909
rect 26424 14900 26476 14952
rect 27436 14900 27488 14952
rect 26700 14832 26752 14884
rect 26148 14764 26200 14816
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 12096 14662 12148 14714
rect 12160 14662 12212 14714
rect 12224 14662 12276 14714
rect 12288 14662 12340 14714
rect 12352 14662 12404 14714
rect 19870 14662 19922 14714
rect 19934 14662 19986 14714
rect 19998 14662 20050 14714
rect 20062 14662 20114 14714
rect 20126 14662 20178 14714
rect 27644 14662 27696 14714
rect 27708 14662 27760 14714
rect 27772 14662 27824 14714
rect 27836 14662 27888 14714
rect 27900 14662 27952 14714
rect 15568 14560 15620 14612
rect 16120 14603 16172 14612
rect 16120 14569 16129 14603
rect 16129 14569 16163 14603
rect 16163 14569 16172 14603
rect 16120 14560 16172 14569
rect 16672 14560 16724 14612
rect 17776 14560 17828 14612
rect 22100 14560 22152 14612
rect 15476 14492 15528 14544
rect 15384 14424 15436 14476
rect 16488 14424 16540 14476
rect 16856 14467 16908 14476
rect 16856 14433 16865 14467
rect 16865 14433 16899 14467
rect 16899 14433 16908 14467
rect 16856 14424 16908 14433
rect 14004 14220 14056 14272
rect 15016 14220 15068 14272
rect 15292 14288 15344 14340
rect 16396 14220 16448 14272
rect 18144 14492 18196 14544
rect 24952 14492 25004 14544
rect 25412 14492 25464 14544
rect 25688 14560 25740 14612
rect 26148 14603 26200 14612
rect 26148 14569 26157 14603
rect 26157 14569 26191 14603
rect 26191 14569 26200 14603
rect 26148 14560 26200 14569
rect 17500 14424 17552 14476
rect 18052 14467 18104 14476
rect 18052 14433 18061 14467
rect 18061 14433 18095 14467
rect 18095 14433 18104 14467
rect 18052 14424 18104 14433
rect 19708 14467 19760 14476
rect 19708 14433 19726 14467
rect 19726 14433 19760 14467
rect 19708 14424 19760 14433
rect 21548 14424 21600 14476
rect 24032 14424 24084 14476
rect 24216 14424 24268 14476
rect 24768 14424 24820 14476
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 26240 14467 26292 14476
rect 26240 14433 26249 14467
rect 26249 14433 26283 14467
rect 26283 14433 26292 14467
rect 26240 14424 26292 14433
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 23572 14288 23624 14340
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 23480 14220 23532 14272
rect 25044 14356 25096 14408
rect 26332 14356 26384 14408
rect 26792 14356 26844 14408
rect 24768 14288 24820 14340
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 25228 14220 25280 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 11436 14118 11488 14170
rect 11500 14118 11552 14170
rect 11564 14118 11616 14170
rect 11628 14118 11680 14170
rect 11692 14118 11744 14170
rect 19210 14118 19262 14170
rect 19274 14118 19326 14170
rect 19338 14118 19390 14170
rect 19402 14118 19454 14170
rect 19466 14118 19518 14170
rect 26984 14118 27036 14170
rect 27048 14118 27100 14170
rect 27112 14118 27164 14170
rect 27176 14118 27228 14170
rect 27240 14118 27292 14170
rect 15292 14059 15344 14068
rect 15292 14025 15301 14059
rect 15301 14025 15335 14059
rect 15335 14025 15344 14059
rect 15292 14016 15344 14025
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 19708 14016 19760 14068
rect 23572 14016 23624 14068
rect 24032 14016 24084 14068
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 18972 13991 19024 14000
rect 18972 13957 18981 13991
rect 18981 13957 19015 13991
rect 19015 13957 19024 13991
rect 18972 13948 19024 13957
rect 24952 14016 25004 14068
rect 25688 13948 25740 14000
rect 18420 13880 18472 13932
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 14004 13812 14056 13864
rect 16672 13812 16724 13864
rect 24492 13812 24544 13864
rect 25964 13880 26016 13932
rect 25504 13855 25556 13864
rect 25504 13821 25513 13855
rect 25513 13821 25547 13855
rect 25547 13821 25556 13855
rect 25504 13812 25556 13821
rect 25780 13855 25832 13864
rect 25780 13821 25789 13855
rect 25789 13821 25823 13855
rect 25823 13821 25832 13855
rect 27988 13880 28040 13932
rect 25780 13812 25832 13821
rect 16396 13787 16448 13796
rect 16396 13753 16430 13787
rect 16430 13753 16448 13787
rect 16396 13744 16448 13753
rect 23296 13787 23348 13796
rect 23296 13753 23305 13787
rect 23305 13753 23339 13787
rect 23339 13753 23348 13787
rect 23296 13744 23348 13753
rect 23480 13787 23532 13796
rect 23480 13753 23505 13787
rect 23505 13753 23532 13787
rect 23480 13744 23532 13753
rect 16028 13719 16080 13728
rect 16028 13685 16037 13719
rect 16037 13685 16071 13719
rect 16071 13685 16080 13719
rect 16028 13676 16080 13685
rect 17592 13719 17644 13728
rect 17592 13685 17601 13719
rect 17601 13685 17635 13719
rect 17635 13685 17644 13719
rect 17592 13676 17644 13685
rect 25228 13744 25280 13796
rect 25688 13787 25740 13796
rect 25688 13753 25697 13787
rect 25697 13753 25731 13787
rect 25731 13753 25740 13787
rect 25688 13744 25740 13753
rect 26148 13744 26200 13796
rect 26240 13744 26292 13796
rect 25872 13676 25924 13728
rect 26424 13676 26476 13728
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 12096 13574 12148 13626
rect 12160 13574 12212 13626
rect 12224 13574 12276 13626
rect 12288 13574 12340 13626
rect 12352 13574 12404 13626
rect 19870 13574 19922 13626
rect 19934 13574 19986 13626
rect 19998 13574 20050 13626
rect 20062 13574 20114 13626
rect 20126 13574 20178 13626
rect 27644 13574 27696 13626
rect 27708 13574 27760 13626
rect 27772 13574 27824 13626
rect 27836 13574 27888 13626
rect 27900 13574 27952 13626
rect 15292 13472 15344 13524
rect 16488 13472 16540 13524
rect 16028 13404 16080 13456
rect 14188 13379 14240 13388
rect 14188 13345 14197 13379
rect 14197 13345 14231 13379
rect 14231 13345 14240 13379
rect 14188 13336 14240 13345
rect 14924 13336 14976 13388
rect 15568 13336 15620 13388
rect 17592 13336 17644 13388
rect 18512 13472 18564 13524
rect 23296 13472 23348 13524
rect 25504 13472 25556 13524
rect 27988 13472 28040 13524
rect 24032 13447 24084 13456
rect 24032 13413 24041 13447
rect 24041 13413 24075 13447
rect 24075 13413 24084 13447
rect 24032 13404 24084 13413
rect 24216 13447 24268 13456
rect 24216 13413 24225 13447
rect 24225 13413 24259 13447
rect 24259 13413 24268 13447
rect 24216 13404 24268 13413
rect 24860 13404 24912 13456
rect 25780 13379 25832 13388
rect 25780 13345 25789 13379
rect 25789 13345 25823 13379
rect 25823 13345 25832 13379
rect 25780 13336 25832 13345
rect 26240 13336 26292 13388
rect 26424 13379 26476 13388
rect 26424 13345 26433 13379
rect 26433 13345 26467 13379
rect 26467 13345 26476 13379
rect 26424 13336 26476 13345
rect 26516 13336 26568 13388
rect 15476 13200 15528 13252
rect 18420 13268 18472 13320
rect 18512 13200 18564 13252
rect 18972 13200 19024 13252
rect 25872 13268 25924 13320
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 25780 13132 25832 13184
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 11436 13030 11488 13082
rect 11500 13030 11552 13082
rect 11564 13030 11616 13082
rect 11628 13030 11680 13082
rect 11692 13030 11744 13082
rect 19210 13030 19262 13082
rect 19274 13030 19326 13082
rect 19338 13030 19390 13082
rect 19402 13030 19454 13082
rect 19466 13030 19518 13082
rect 26984 13030 27036 13082
rect 27048 13030 27100 13082
rect 27112 13030 27164 13082
rect 27176 13030 27228 13082
rect 27240 13030 27292 13082
rect 14924 12928 14976 12980
rect 16672 12971 16724 12980
rect 16672 12937 16681 12971
rect 16681 12937 16715 12971
rect 16715 12937 16724 12971
rect 16672 12928 16724 12937
rect 26516 12928 26568 12980
rect 16856 12792 16908 12844
rect 15016 12724 15068 12776
rect 16120 12724 16172 12776
rect 16580 12724 16632 12776
rect 16488 12656 16540 12708
rect 17500 12724 17552 12776
rect 18420 12724 18472 12776
rect 18880 12767 18932 12776
rect 18880 12733 18889 12767
rect 18889 12733 18923 12767
rect 18923 12733 18932 12767
rect 18880 12724 18932 12733
rect 26332 12860 26384 12912
rect 25688 12792 25740 12844
rect 25780 12767 25832 12776
rect 25780 12733 25789 12767
rect 25789 12733 25823 12767
rect 25823 12733 25832 12767
rect 25780 12724 25832 12733
rect 18052 12699 18104 12708
rect 18052 12665 18061 12699
rect 18061 12665 18095 12699
rect 18095 12665 18104 12699
rect 18052 12656 18104 12665
rect 25228 12656 25280 12708
rect 15568 12588 15620 12640
rect 17132 12631 17184 12640
rect 17132 12597 17141 12631
rect 17141 12597 17175 12631
rect 17175 12597 17184 12631
rect 17132 12588 17184 12597
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 18328 12588 18380 12640
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 12096 12486 12148 12538
rect 12160 12486 12212 12538
rect 12224 12486 12276 12538
rect 12288 12486 12340 12538
rect 12352 12486 12404 12538
rect 19870 12486 19922 12538
rect 19934 12486 19986 12538
rect 19998 12486 20050 12538
rect 20062 12486 20114 12538
rect 20126 12486 20178 12538
rect 27644 12486 27696 12538
rect 27708 12486 27760 12538
rect 27772 12486 27824 12538
rect 27836 12486 27888 12538
rect 27900 12486 27952 12538
rect 16488 12384 16540 12436
rect 17500 12384 17552 12436
rect 18052 12384 18104 12436
rect 18512 12359 18564 12368
rect 18512 12325 18546 12359
rect 18546 12325 18564 12359
rect 16856 12291 16908 12300
rect 16856 12257 16865 12291
rect 16865 12257 16899 12291
rect 16899 12257 16908 12291
rect 16856 12248 16908 12257
rect 18512 12316 18564 12325
rect 17960 12248 18012 12300
rect 18328 12248 18380 12300
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 18236 12044 18288 12096
rect 18972 12044 19024 12096
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 11436 11942 11488 11994
rect 11500 11942 11552 11994
rect 11564 11942 11616 11994
rect 11628 11942 11680 11994
rect 11692 11942 11744 11994
rect 19210 11942 19262 11994
rect 19274 11942 19326 11994
rect 19338 11942 19390 11994
rect 19402 11942 19454 11994
rect 19466 11942 19518 11994
rect 26984 11942 27036 11994
rect 27048 11942 27100 11994
rect 27112 11942 27164 11994
rect 27176 11942 27228 11994
rect 27240 11942 27292 11994
rect 16580 11840 16632 11892
rect 17960 11840 18012 11892
rect 16856 11679 16908 11688
rect 16856 11645 16865 11679
rect 16865 11645 16899 11679
rect 16899 11645 16908 11679
rect 16856 11636 16908 11645
rect 17132 11679 17184 11688
rect 17132 11645 17166 11679
rect 17166 11645 17184 11679
rect 17132 11636 17184 11645
rect 15660 11568 15712 11620
rect 16764 11500 16816 11552
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 12096 11398 12148 11450
rect 12160 11398 12212 11450
rect 12224 11398 12276 11450
rect 12288 11398 12340 11450
rect 12352 11398 12404 11450
rect 19870 11398 19922 11450
rect 19934 11398 19986 11450
rect 19998 11398 20050 11450
rect 20062 11398 20114 11450
rect 20126 11398 20178 11450
rect 27644 11398 27696 11450
rect 27708 11398 27760 11450
rect 27772 11398 27824 11450
rect 27836 11398 27888 11450
rect 27900 11398 27952 11450
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 16856 11296 16908 11348
rect 15568 11203 15620 11212
rect 15568 11169 15577 11203
rect 15577 11169 15611 11203
rect 15611 11169 15620 11203
rect 15568 11160 15620 11169
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 18880 11160 18932 11212
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 11436 10854 11488 10906
rect 11500 10854 11552 10906
rect 11564 10854 11616 10906
rect 11628 10854 11680 10906
rect 11692 10854 11744 10906
rect 19210 10854 19262 10906
rect 19274 10854 19326 10906
rect 19338 10854 19390 10906
rect 19402 10854 19454 10906
rect 19466 10854 19518 10906
rect 26984 10854 27036 10906
rect 27048 10854 27100 10906
rect 27112 10854 27164 10906
rect 27176 10854 27228 10906
rect 27240 10854 27292 10906
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 12096 10310 12148 10362
rect 12160 10310 12212 10362
rect 12224 10310 12276 10362
rect 12288 10310 12340 10362
rect 12352 10310 12404 10362
rect 19870 10310 19922 10362
rect 19934 10310 19986 10362
rect 19998 10310 20050 10362
rect 20062 10310 20114 10362
rect 20126 10310 20178 10362
rect 27644 10310 27696 10362
rect 27708 10310 27760 10362
rect 27772 10310 27824 10362
rect 27836 10310 27888 10362
rect 27900 10310 27952 10362
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 11436 9766 11488 9818
rect 11500 9766 11552 9818
rect 11564 9766 11616 9818
rect 11628 9766 11680 9818
rect 11692 9766 11744 9818
rect 19210 9766 19262 9818
rect 19274 9766 19326 9818
rect 19338 9766 19390 9818
rect 19402 9766 19454 9818
rect 19466 9766 19518 9818
rect 26984 9766 27036 9818
rect 27048 9766 27100 9818
rect 27112 9766 27164 9818
rect 27176 9766 27228 9818
rect 27240 9766 27292 9818
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 12096 9222 12148 9274
rect 12160 9222 12212 9274
rect 12224 9222 12276 9274
rect 12288 9222 12340 9274
rect 12352 9222 12404 9274
rect 19870 9222 19922 9274
rect 19934 9222 19986 9274
rect 19998 9222 20050 9274
rect 20062 9222 20114 9274
rect 20126 9222 20178 9274
rect 27644 9222 27696 9274
rect 27708 9222 27760 9274
rect 27772 9222 27824 9274
rect 27836 9222 27888 9274
rect 27900 9222 27952 9274
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 11436 8678 11488 8730
rect 11500 8678 11552 8730
rect 11564 8678 11616 8730
rect 11628 8678 11680 8730
rect 11692 8678 11744 8730
rect 19210 8678 19262 8730
rect 19274 8678 19326 8730
rect 19338 8678 19390 8730
rect 19402 8678 19454 8730
rect 19466 8678 19518 8730
rect 26984 8678 27036 8730
rect 27048 8678 27100 8730
rect 27112 8678 27164 8730
rect 27176 8678 27228 8730
rect 27240 8678 27292 8730
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 12096 8134 12148 8186
rect 12160 8134 12212 8186
rect 12224 8134 12276 8186
rect 12288 8134 12340 8186
rect 12352 8134 12404 8186
rect 19870 8134 19922 8186
rect 19934 8134 19986 8186
rect 19998 8134 20050 8186
rect 20062 8134 20114 8186
rect 20126 8134 20178 8186
rect 27644 8134 27696 8186
rect 27708 8134 27760 8186
rect 27772 8134 27824 8186
rect 27836 8134 27888 8186
rect 27900 8134 27952 8186
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 11436 7590 11488 7642
rect 11500 7590 11552 7642
rect 11564 7590 11616 7642
rect 11628 7590 11680 7642
rect 11692 7590 11744 7642
rect 19210 7590 19262 7642
rect 19274 7590 19326 7642
rect 19338 7590 19390 7642
rect 19402 7590 19454 7642
rect 19466 7590 19518 7642
rect 26984 7590 27036 7642
rect 27048 7590 27100 7642
rect 27112 7590 27164 7642
rect 27176 7590 27228 7642
rect 27240 7590 27292 7642
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 12096 7046 12148 7098
rect 12160 7046 12212 7098
rect 12224 7046 12276 7098
rect 12288 7046 12340 7098
rect 12352 7046 12404 7098
rect 19870 7046 19922 7098
rect 19934 7046 19986 7098
rect 19998 7046 20050 7098
rect 20062 7046 20114 7098
rect 20126 7046 20178 7098
rect 27644 7046 27696 7098
rect 27708 7046 27760 7098
rect 27772 7046 27824 7098
rect 27836 7046 27888 7098
rect 27900 7046 27952 7098
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 11436 6502 11488 6554
rect 11500 6502 11552 6554
rect 11564 6502 11616 6554
rect 11628 6502 11680 6554
rect 11692 6502 11744 6554
rect 19210 6502 19262 6554
rect 19274 6502 19326 6554
rect 19338 6502 19390 6554
rect 19402 6502 19454 6554
rect 19466 6502 19518 6554
rect 26984 6502 27036 6554
rect 27048 6502 27100 6554
rect 27112 6502 27164 6554
rect 27176 6502 27228 6554
rect 27240 6502 27292 6554
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 12096 5958 12148 6010
rect 12160 5958 12212 6010
rect 12224 5958 12276 6010
rect 12288 5958 12340 6010
rect 12352 5958 12404 6010
rect 19870 5958 19922 6010
rect 19934 5958 19986 6010
rect 19998 5958 20050 6010
rect 20062 5958 20114 6010
rect 20126 5958 20178 6010
rect 27644 5958 27696 6010
rect 27708 5958 27760 6010
rect 27772 5958 27824 6010
rect 27836 5958 27888 6010
rect 27900 5958 27952 6010
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 11436 5414 11488 5466
rect 11500 5414 11552 5466
rect 11564 5414 11616 5466
rect 11628 5414 11680 5466
rect 11692 5414 11744 5466
rect 19210 5414 19262 5466
rect 19274 5414 19326 5466
rect 19338 5414 19390 5466
rect 19402 5414 19454 5466
rect 19466 5414 19518 5466
rect 26984 5414 27036 5466
rect 27048 5414 27100 5466
rect 27112 5414 27164 5466
rect 27176 5414 27228 5466
rect 27240 5414 27292 5466
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 12096 4870 12148 4922
rect 12160 4870 12212 4922
rect 12224 4870 12276 4922
rect 12288 4870 12340 4922
rect 12352 4870 12404 4922
rect 19870 4870 19922 4922
rect 19934 4870 19986 4922
rect 19998 4870 20050 4922
rect 20062 4870 20114 4922
rect 20126 4870 20178 4922
rect 27644 4870 27696 4922
rect 27708 4870 27760 4922
rect 27772 4870 27824 4922
rect 27836 4870 27888 4922
rect 27900 4870 27952 4922
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 11436 4326 11488 4378
rect 11500 4326 11552 4378
rect 11564 4326 11616 4378
rect 11628 4326 11680 4378
rect 11692 4326 11744 4378
rect 19210 4326 19262 4378
rect 19274 4326 19326 4378
rect 19338 4326 19390 4378
rect 19402 4326 19454 4378
rect 19466 4326 19518 4378
rect 26984 4326 27036 4378
rect 27048 4326 27100 4378
rect 27112 4326 27164 4378
rect 27176 4326 27228 4378
rect 27240 4326 27292 4378
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 12096 3782 12148 3834
rect 12160 3782 12212 3834
rect 12224 3782 12276 3834
rect 12288 3782 12340 3834
rect 12352 3782 12404 3834
rect 19870 3782 19922 3834
rect 19934 3782 19986 3834
rect 19998 3782 20050 3834
rect 20062 3782 20114 3834
rect 20126 3782 20178 3834
rect 27644 3782 27696 3834
rect 27708 3782 27760 3834
rect 27772 3782 27824 3834
rect 27836 3782 27888 3834
rect 27900 3782 27952 3834
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 11436 3238 11488 3290
rect 11500 3238 11552 3290
rect 11564 3238 11616 3290
rect 11628 3238 11680 3290
rect 11692 3238 11744 3290
rect 19210 3238 19262 3290
rect 19274 3238 19326 3290
rect 19338 3238 19390 3290
rect 19402 3238 19454 3290
rect 19466 3238 19518 3290
rect 26984 3238 27036 3290
rect 27048 3238 27100 3290
rect 27112 3238 27164 3290
rect 27176 3238 27228 3290
rect 27240 3238 27292 3290
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 12096 2694 12148 2746
rect 12160 2694 12212 2746
rect 12224 2694 12276 2746
rect 12288 2694 12340 2746
rect 12352 2694 12404 2746
rect 19870 2694 19922 2746
rect 19934 2694 19986 2746
rect 19998 2694 20050 2746
rect 20062 2694 20114 2746
rect 20126 2694 20178 2746
rect 27644 2694 27696 2746
rect 27708 2694 27760 2746
rect 27772 2694 27824 2746
rect 27836 2694 27888 2746
rect 27900 2694 27952 2746
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 11436 2150 11488 2202
rect 11500 2150 11552 2202
rect 11564 2150 11616 2202
rect 11628 2150 11680 2202
rect 11692 2150 11744 2202
rect 19210 2150 19262 2202
rect 19274 2150 19326 2202
rect 19338 2150 19390 2202
rect 19402 2150 19454 2202
rect 19466 2150 19518 2202
rect 26984 2150 27036 2202
rect 27048 2150 27100 2202
rect 27112 2150 27164 2202
rect 27176 2150 27228 2202
rect 27240 2150 27292 2202
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 12096 1606 12148 1658
rect 12160 1606 12212 1658
rect 12224 1606 12276 1658
rect 12288 1606 12340 1658
rect 12352 1606 12404 1658
rect 19870 1606 19922 1658
rect 19934 1606 19986 1658
rect 19998 1606 20050 1658
rect 20062 1606 20114 1658
rect 20126 1606 20178 1658
rect 27644 1606 27696 1658
rect 27708 1606 27760 1658
rect 27772 1606 27824 1658
rect 27836 1606 27888 1658
rect 27900 1606 27952 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 11436 1062 11488 1114
rect 11500 1062 11552 1114
rect 11564 1062 11616 1114
rect 11628 1062 11680 1114
rect 11692 1062 11744 1114
rect 19210 1062 19262 1114
rect 19274 1062 19326 1114
rect 19338 1062 19390 1114
rect 19402 1062 19454 1114
rect 19466 1062 19518 1114
rect 26984 1062 27036 1114
rect 27048 1062 27100 1114
rect 27112 1062 27164 1114
rect 27176 1062 27228 1114
rect 27240 1062 27292 1114
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 12096 518 12148 570
rect 12160 518 12212 570
rect 12224 518 12276 570
rect 12288 518 12340 570
rect 12352 518 12404 570
rect 19870 518 19922 570
rect 19934 518 19986 570
rect 19998 518 20050 570
rect 20062 518 20114 570
rect 20126 518 20178 570
rect 27644 518 27696 570
rect 27708 518 27760 570
rect 27772 518 27824 570
rect 27836 518 27888 570
rect 27900 518 27952 570
<< metal2 >>
rect 11794 44840 11850 44849
rect 11794 44775 11850 44784
rect 13082 44840 13138 44849
rect 13082 44775 13138 44784
rect 21638 44840 21694 44849
rect 21638 44775 21694 44784
rect 27434 44840 27490 44849
rect 27434 44775 27490 44784
rect 28170 44840 28226 44849
rect 28170 44775 28226 44784
rect 3662 44636 3970 44645
rect 3662 44634 3668 44636
rect 3724 44634 3748 44636
rect 3804 44634 3828 44636
rect 3884 44634 3908 44636
rect 3964 44634 3970 44636
rect 3724 44582 3726 44634
rect 3906 44582 3908 44634
rect 3662 44580 3668 44582
rect 3724 44580 3748 44582
rect 3804 44580 3828 44582
rect 3884 44580 3908 44582
rect 3964 44580 3970 44582
rect 3662 44571 3970 44580
rect 11436 44636 11744 44645
rect 11436 44634 11442 44636
rect 11498 44634 11522 44636
rect 11578 44634 11602 44636
rect 11658 44634 11682 44636
rect 11738 44634 11744 44636
rect 11498 44582 11500 44634
rect 11680 44582 11682 44634
rect 11436 44580 11442 44582
rect 11498 44580 11522 44582
rect 11578 44580 11602 44582
rect 11658 44580 11682 44582
rect 11738 44580 11744 44582
rect 7194 44568 7250 44577
rect 7194 44503 7196 44512
rect 7248 44503 7250 44512
rect 7654 44568 7710 44577
rect 7654 44503 7656 44512
rect 7196 44474 7248 44480
rect 7708 44503 7710 44512
rect 8298 44568 8354 44577
rect 8298 44503 8300 44512
rect 7656 44474 7708 44480
rect 8352 44503 8354 44512
rect 8758 44568 8814 44577
rect 8758 44503 8760 44512
rect 8300 44474 8352 44480
rect 8812 44503 8814 44512
rect 9310 44568 9366 44577
rect 11436 44571 11744 44580
rect 11808 44538 11836 44775
rect 12806 44568 12862 44577
rect 9310 44503 9312 44512
rect 8760 44474 8812 44480
rect 9364 44503 9366 44512
rect 11796 44532 11848 44538
rect 9312 44474 9364 44480
rect 13096 44538 13124 44775
rect 19210 44636 19518 44645
rect 19210 44634 19216 44636
rect 19272 44634 19296 44636
rect 19352 44634 19376 44636
rect 19432 44634 19456 44636
rect 19512 44634 19518 44636
rect 19272 44582 19274 44634
rect 19454 44582 19456 44634
rect 19210 44580 19216 44582
rect 19272 44580 19296 44582
rect 19352 44580 19376 44582
rect 19432 44580 19456 44582
rect 19512 44580 19518 44582
rect 19210 44571 19518 44580
rect 12806 44503 12808 44512
rect 11796 44474 11848 44480
rect 12860 44503 12862 44512
rect 13084 44532 13136 44538
rect 12808 44474 12860 44480
rect 13084 44474 13136 44480
rect 11888 44396 11940 44402
rect 11888 44338 11940 44344
rect 8208 44328 8260 44334
rect 8208 44270 8260 44276
rect 4322 44092 4630 44101
rect 4322 44090 4328 44092
rect 4384 44090 4408 44092
rect 4464 44090 4488 44092
rect 4544 44090 4568 44092
rect 4624 44090 4630 44092
rect 4384 44038 4386 44090
rect 4566 44038 4568 44090
rect 4322 44036 4328 44038
rect 4384 44036 4408 44038
rect 4464 44036 4488 44038
rect 4544 44036 4568 44038
rect 4624 44036 4630 44038
rect 4322 44027 4630 44036
rect 6550 44024 6606 44033
rect 6550 43959 6552 43968
rect 6604 43959 6606 43968
rect 6918 44024 6974 44033
rect 8220 43994 8248 44270
rect 11060 44260 11112 44266
rect 11060 44202 11112 44208
rect 8300 44192 8352 44198
rect 8300 44134 8352 44140
rect 6918 43959 6920 43968
rect 6552 43930 6604 43936
rect 6972 43959 6974 43968
rect 8208 43988 8260 43994
rect 6920 43930 6972 43936
rect 8208 43930 8260 43936
rect 8220 43858 8248 43930
rect 8312 43858 8340 44134
rect 10690 44024 10746 44033
rect 10690 43959 10692 43968
rect 10744 43959 10746 43968
rect 10692 43930 10744 43936
rect 8208 43852 8260 43858
rect 8208 43794 8260 43800
rect 8300 43852 8352 43858
rect 8300 43794 8352 43800
rect 8852 43852 8904 43858
rect 8852 43794 8904 43800
rect 3662 43548 3970 43557
rect 3662 43546 3668 43548
rect 3724 43546 3748 43548
rect 3804 43546 3828 43548
rect 3884 43546 3908 43548
rect 3964 43546 3970 43548
rect 3724 43494 3726 43546
rect 3906 43494 3908 43546
rect 3662 43492 3668 43494
rect 3724 43492 3748 43494
rect 3804 43492 3828 43494
rect 3884 43492 3908 43494
rect 3964 43492 3970 43494
rect 3662 43483 3970 43492
rect 8864 43450 8892 43794
rect 9772 43648 9824 43654
rect 9772 43590 9824 43596
rect 10968 43648 11020 43654
rect 10968 43590 11020 43596
rect 8852 43444 8904 43450
rect 8852 43386 8904 43392
rect 9784 43382 9812 43590
rect 9772 43376 9824 43382
rect 9772 43318 9824 43324
rect 10980 43246 11008 43590
rect 9404 43240 9456 43246
rect 9404 43182 9456 43188
rect 10324 43240 10376 43246
rect 10324 43182 10376 43188
rect 10968 43240 11020 43246
rect 10968 43182 11020 43188
rect 4322 43004 4630 43013
rect 4322 43002 4328 43004
rect 4384 43002 4408 43004
rect 4464 43002 4488 43004
rect 4544 43002 4568 43004
rect 4624 43002 4630 43004
rect 4384 42950 4386 43002
rect 4566 42950 4568 43002
rect 4322 42948 4328 42950
rect 4384 42948 4408 42950
rect 4464 42948 4488 42950
rect 4544 42948 4568 42950
rect 4624 42948 4630 42950
rect 4322 42939 4630 42948
rect 9416 42770 9444 43182
rect 9404 42764 9456 42770
rect 9404 42706 9456 42712
rect 9680 42764 9732 42770
rect 9680 42706 9732 42712
rect 3662 42460 3970 42469
rect 3662 42458 3668 42460
rect 3724 42458 3748 42460
rect 3804 42458 3828 42460
rect 3884 42458 3908 42460
rect 3964 42458 3970 42460
rect 3724 42406 3726 42458
rect 3906 42406 3908 42458
rect 3662 42404 3668 42406
rect 3724 42404 3748 42406
rect 3804 42404 3828 42406
rect 3884 42404 3908 42406
rect 3964 42404 3970 42406
rect 3662 42395 3970 42404
rect 4322 41916 4630 41925
rect 4322 41914 4328 41916
rect 4384 41914 4408 41916
rect 4464 41914 4488 41916
rect 4544 41914 4568 41916
rect 4624 41914 4630 41916
rect 4384 41862 4386 41914
rect 4566 41862 4568 41914
rect 4322 41860 4328 41862
rect 4384 41860 4408 41862
rect 4464 41860 4488 41862
rect 4544 41860 4568 41862
rect 4624 41860 4630 41862
rect 4322 41851 4630 41860
rect 9692 41818 9720 42706
rect 9680 41812 9732 41818
rect 9680 41754 9732 41760
rect 10336 41682 10364 43182
rect 11072 43178 11100 44202
rect 11334 43888 11390 43897
rect 11244 43852 11296 43858
rect 11334 43823 11390 43832
rect 11244 43794 11296 43800
rect 11060 43172 11112 43178
rect 11060 43114 11112 43120
rect 11072 42770 11100 43114
rect 11060 42764 11112 42770
rect 11060 42706 11112 42712
rect 10968 42560 11020 42566
rect 10968 42502 11020 42508
rect 10980 41750 11008 42502
rect 10968 41744 11020 41750
rect 10968 41686 11020 41692
rect 10140 41676 10192 41682
rect 10140 41618 10192 41624
rect 10324 41676 10376 41682
rect 10324 41618 10376 41624
rect 10784 41676 10836 41682
rect 10784 41618 10836 41624
rect 3662 41372 3970 41381
rect 3662 41370 3668 41372
rect 3724 41370 3748 41372
rect 3804 41370 3828 41372
rect 3884 41370 3908 41372
rect 3964 41370 3970 41372
rect 3724 41318 3726 41370
rect 3906 41318 3908 41370
rect 3662 41316 3668 41318
rect 3724 41316 3748 41318
rect 3804 41316 3828 41318
rect 3884 41316 3908 41318
rect 3964 41316 3970 41318
rect 3662 41307 3970 41316
rect 10152 41274 10180 41618
rect 9680 41268 9732 41274
rect 9680 41210 9732 41216
rect 10140 41268 10192 41274
rect 10140 41210 10192 41216
rect 9220 41200 9272 41206
rect 9220 41142 9272 41148
rect 9232 41070 9260 41142
rect 9496 41132 9548 41138
rect 9496 41074 9548 41080
rect 8300 41064 8352 41070
rect 8300 41006 8352 41012
rect 8944 41064 8996 41070
rect 8944 41006 8996 41012
rect 9220 41064 9272 41070
rect 9220 41006 9272 41012
rect 8116 40928 8168 40934
rect 8116 40870 8168 40876
rect 4322 40828 4630 40837
rect 4322 40826 4328 40828
rect 4384 40826 4408 40828
rect 4464 40826 4488 40828
rect 4544 40826 4568 40828
rect 4624 40826 4630 40828
rect 4384 40774 4386 40826
rect 4566 40774 4568 40826
rect 4322 40772 4328 40774
rect 4384 40772 4408 40774
rect 4464 40772 4488 40774
rect 4544 40772 4568 40774
rect 4624 40772 4630 40774
rect 4322 40763 4630 40772
rect 8128 40594 8156 40870
rect 8116 40588 8168 40594
rect 8116 40530 8168 40536
rect 3662 40284 3970 40293
rect 3662 40282 3668 40284
rect 3724 40282 3748 40284
rect 3804 40282 3828 40284
rect 3884 40282 3908 40284
rect 3964 40282 3970 40284
rect 3724 40230 3726 40282
rect 3906 40230 3908 40282
rect 3662 40228 3668 40230
rect 3724 40228 3748 40230
rect 3804 40228 3828 40230
rect 3884 40228 3908 40230
rect 3964 40228 3970 40230
rect 3662 40219 3970 40228
rect 4322 39740 4630 39749
rect 4322 39738 4328 39740
rect 4384 39738 4408 39740
rect 4464 39738 4488 39740
rect 4544 39738 4568 39740
rect 4624 39738 4630 39740
rect 4384 39686 4386 39738
rect 4566 39686 4568 39738
rect 4322 39684 4328 39686
rect 4384 39684 4408 39686
rect 4464 39684 4488 39686
rect 4544 39684 4568 39686
rect 4624 39684 4630 39686
rect 4322 39675 4630 39684
rect 3662 39196 3970 39205
rect 3662 39194 3668 39196
rect 3724 39194 3748 39196
rect 3804 39194 3828 39196
rect 3884 39194 3908 39196
rect 3964 39194 3970 39196
rect 3724 39142 3726 39194
rect 3906 39142 3908 39194
rect 3662 39140 3668 39142
rect 3724 39140 3748 39142
rect 3804 39140 3828 39142
rect 3884 39140 3908 39142
rect 3964 39140 3970 39142
rect 3662 39131 3970 39140
rect 8312 38894 8340 41006
rect 8668 40928 8720 40934
rect 8668 40870 8720 40876
rect 8680 40050 8708 40870
rect 8956 40662 8984 41006
rect 9128 40928 9180 40934
rect 9128 40870 9180 40876
rect 8944 40656 8996 40662
rect 8944 40598 8996 40604
rect 8852 40588 8904 40594
rect 8852 40530 8904 40536
rect 8864 40186 8892 40530
rect 8852 40180 8904 40186
rect 8852 40122 8904 40128
rect 8668 40044 8720 40050
rect 8668 39986 8720 39992
rect 9140 39982 9168 40870
rect 9508 40390 9536 41074
rect 9588 40588 9640 40594
rect 9588 40530 9640 40536
rect 9496 40384 9548 40390
rect 9496 40326 9548 40332
rect 9128 39976 9180 39982
rect 9128 39918 9180 39924
rect 9220 39976 9272 39982
rect 9220 39918 9272 39924
rect 8392 39840 8444 39846
rect 8392 39782 8444 39788
rect 8404 39506 8432 39782
rect 8392 39500 8444 39506
rect 8392 39442 8444 39448
rect 9232 39438 9260 39918
rect 9220 39432 9272 39438
rect 9220 39374 9272 39380
rect 8300 38888 8352 38894
rect 8300 38830 8352 38836
rect 9128 38888 9180 38894
rect 9128 38830 9180 38836
rect 4322 38652 4630 38661
rect 4322 38650 4328 38652
rect 4384 38650 4408 38652
rect 4464 38650 4488 38652
rect 4544 38650 4568 38652
rect 4624 38650 4630 38652
rect 4384 38598 4386 38650
rect 4566 38598 4568 38650
rect 4322 38596 4328 38598
rect 4384 38596 4408 38598
rect 4464 38596 4488 38598
rect 4544 38596 4568 38598
rect 4624 38596 4630 38598
rect 4322 38587 4630 38596
rect 3662 38108 3970 38117
rect 3662 38106 3668 38108
rect 3724 38106 3748 38108
rect 3804 38106 3828 38108
rect 3884 38106 3908 38108
rect 3964 38106 3970 38108
rect 3724 38054 3726 38106
rect 3906 38054 3908 38106
rect 3662 38052 3668 38054
rect 3724 38052 3748 38054
rect 3804 38052 3828 38054
rect 3884 38052 3908 38054
rect 3964 38052 3970 38054
rect 3662 38043 3970 38052
rect 8312 37942 8340 38830
rect 8484 38752 8536 38758
rect 8484 38694 8536 38700
rect 8496 38486 8524 38694
rect 8484 38480 8536 38486
rect 8484 38422 8536 38428
rect 8300 37936 8352 37942
rect 8300 37878 8352 37884
rect 4322 37564 4630 37573
rect 4322 37562 4328 37564
rect 4384 37562 4408 37564
rect 4464 37562 4488 37564
rect 4544 37562 4568 37564
rect 4624 37562 4630 37564
rect 4384 37510 4386 37562
rect 4566 37510 4568 37562
rect 4322 37508 4328 37510
rect 4384 37508 4408 37510
rect 4464 37508 4488 37510
rect 4544 37508 4568 37510
rect 4624 37508 4630 37510
rect 4322 37499 4630 37508
rect 3662 37020 3970 37029
rect 3662 37018 3668 37020
rect 3724 37018 3748 37020
rect 3804 37018 3828 37020
rect 3884 37018 3908 37020
rect 3964 37018 3970 37020
rect 3724 36966 3726 37018
rect 3906 36966 3908 37018
rect 3662 36964 3668 36966
rect 3724 36964 3748 36966
rect 3804 36964 3828 36966
rect 3884 36964 3908 36966
rect 3964 36964 3970 36966
rect 3662 36955 3970 36964
rect 8312 36786 8340 37878
rect 9140 37466 9168 38830
rect 9508 37806 9536 40326
rect 9600 40066 9628 40530
rect 9692 40186 9720 41210
rect 10336 41154 10364 41618
rect 10416 41608 10468 41614
rect 10416 41550 10468 41556
rect 10428 41414 10456 41550
rect 10428 41386 10548 41414
rect 10336 41126 10456 41154
rect 9772 41064 9824 41070
rect 9772 41006 9824 41012
rect 10140 41064 10192 41070
rect 10140 41006 10192 41012
rect 10324 41064 10376 41070
rect 10324 41006 10376 41012
rect 9680 40180 9732 40186
rect 9680 40122 9732 40128
rect 9600 40050 9720 40066
rect 9588 40044 9720 40050
rect 9640 40038 9720 40044
rect 9588 39986 9640 39992
rect 9588 39840 9640 39846
rect 9588 39782 9640 39788
rect 9600 38962 9628 39782
rect 9692 39302 9720 40038
rect 9784 39642 9812 41006
rect 10152 40730 10180 41006
rect 10140 40724 10192 40730
rect 10140 40666 10192 40672
rect 10232 40656 10284 40662
rect 10336 40644 10364 41006
rect 10284 40616 10364 40644
rect 10232 40598 10284 40604
rect 9864 40452 9916 40458
rect 9864 40394 9916 40400
rect 9772 39636 9824 39642
rect 9772 39578 9824 39584
rect 9772 39500 9824 39506
rect 9876 39488 9904 40394
rect 10140 40112 10192 40118
rect 10140 40054 10192 40060
rect 9956 39976 10008 39982
rect 9956 39918 10008 39924
rect 9968 39506 9996 39918
rect 10048 39568 10100 39574
rect 10048 39510 10100 39516
rect 9824 39460 9904 39488
rect 9956 39500 10008 39506
rect 9772 39442 9824 39448
rect 9956 39442 10008 39448
rect 9784 39370 9812 39442
rect 9772 39364 9824 39370
rect 9772 39306 9824 39312
rect 9680 39296 9732 39302
rect 9680 39238 9732 39244
rect 9588 38956 9640 38962
rect 9588 38898 9640 38904
rect 9600 38554 9628 38898
rect 9680 38888 9732 38894
rect 9680 38830 9732 38836
rect 9588 38548 9640 38554
rect 9588 38490 9640 38496
rect 9496 37800 9548 37806
rect 9232 37760 9496 37788
rect 9128 37460 9180 37466
rect 9128 37402 9180 37408
rect 9232 37346 9260 37760
rect 9496 37742 9548 37748
rect 9496 37664 9548 37670
rect 9496 37606 9548 37612
rect 9140 37330 9260 37346
rect 9508 37330 9536 37606
rect 9128 37324 9260 37330
rect 9180 37318 9260 37324
rect 9496 37324 9548 37330
rect 9128 37266 9180 37272
rect 9496 37266 9548 37272
rect 9312 37120 9364 37126
rect 9312 37062 9364 37068
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 4322 36476 4630 36485
rect 4322 36474 4328 36476
rect 4384 36474 4408 36476
rect 4464 36474 4488 36476
rect 4544 36474 4568 36476
rect 4624 36474 4630 36476
rect 4384 36422 4386 36474
rect 4566 36422 4568 36474
rect 4322 36420 4328 36422
rect 4384 36420 4408 36422
rect 4464 36420 4488 36422
rect 4544 36420 4568 36422
rect 4624 36420 4630 36422
rect 4322 36411 4630 36420
rect 3662 35932 3970 35941
rect 3662 35930 3668 35932
rect 3724 35930 3748 35932
rect 3804 35930 3828 35932
rect 3884 35930 3908 35932
rect 3964 35930 3970 35932
rect 3724 35878 3726 35930
rect 3906 35878 3908 35930
rect 3662 35876 3668 35878
rect 3724 35876 3748 35878
rect 3804 35876 3828 35878
rect 3884 35876 3908 35878
rect 3964 35876 3970 35878
rect 3662 35867 3970 35876
rect 8312 35698 8340 36722
rect 9036 36644 9088 36650
rect 9036 36586 9088 36592
rect 9048 36378 9076 36586
rect 9036 36372 9088 36378
rect 9036 36314 9088 36320
rect 9324 36242 9352 37062
rect 9600 36718 9628 38490
rect 9692 38010 9720 38830
rect 9680 38004 9732 38010
rect 9680 37946 9732 37952
rect 9784 37398 9812 39306
rect 10060 38978 10088 39510
rect 9968 38950 10088 38978
rect 9864 38752 9916 38758
rect 9864 38694 9916 38700
rect 9876 38418 9904 38694
rect 9864 38412 9916 38418
rect 9864 38354 9916 38360
rect 9864 38276 9916 38282
rect 9864 38218 9916 38224
rect 9772 37392 9824 37398
rect 9772 37334 9824 37340
rect 9588 36712 9640 36718
rect 9588 36654 9640 36660
rect 9312 36236 9364 36242
rect 9312 36178 9364 36184
rect 9600 36174 9628 36654
rect 9876 36378 9904 38218
rect 9968 37466 9996 38950
rect 10048 38820 10100 38826
rect 10048 38762 10100 38768
rect 10060 38418 10088 38762
rect 10048 38412 10100 38418
rect 10048 38354 10100 38360
rect 10152 38214 10180 40054
rect 10336 39914 10364 40616
rect 10232 39908 10284 39914
rect 10232 39850 10284 39856
rect 10324 39908 10376 39914
rect 10324 39850 10376 39856
rect 10244 39794 10272 39850
rect 10428 39794 10456 41126
rect 10244 39766 10456 39794
rect 10244 38418 10272 39766
rect 10416 39296 10468 39302
rect 10416 39238 10468 39244
rect 10232 38412 10284 38418
rect 10232 38354 10284 38360
rect 10244 38282 10272 38354
rect 10232 38276 10284 38282
rect 10232 38218 10284 38224
rect 10140 38208 10192 38214
rect 10060 38168 10140 38196
rect 9956 37460 10008 37466
rect 9956 37402 10008 37408
rect 9864 36372 9916 36378
rect 9864 36314 9916 36320
rect 9588 36168 9640 36174
rect 9588 36110 9640 36116
rect 8300 35692 8352 35698
rect 9968 35680 9996 37402
rect 10060 35834 10088 38168
rect 10140 38150 10192 38156
rect 10140 37868 10192 37874
rect 10140 37810 10192 37816
rect 10152 37330 10180 37810
rect 10140 37324 10192 37330
rect 10140 37266 10192 37272
rect 10152 36922 10180 37266
rect 10140 36916 10192 36922
rect 10140 36858 10192 36864
rect 10048 35828 10100 35834
rect 10048 35770 10100 35776
rect 8300 35634 8352 35640
rect 9876 35652 9996 35680
rect 9496 35624 9548 35630
rect 9496 35566 9548 35572
rect 9772 35624 9824 35630
rect 9876 35612 9904 35652
rect 9824 35584 9904 35612
rect 9772 35566 9824 35572
rect 4322 35388 4630 35397
rect 4322 35386 4328 35388
rect 4384 35386 4408 35388
rect 4464 35386 4488 35388
rect 4544 35386 4568 35388
rect 4624 35386 4630 35388
rect 4384 35334 4386 35386
rect 4566 35334 4568 35386
rect 4322 35332 4328 35334
rect 4384 35332 4408 35334
rect 4464 35332 4488 35334
rect 4544 35332 4568 35334
rect 4624 35332 4630 35334
rect 4322 35323 4630 35332
rect 3662 34844 3970 34853
rect 3662 34842 3668 34844
rect 3724 34842 3748 34844
rect 3804 34842 3828 34844
rect 3884 34842 3908 34844
rect 3964 34842 3970 34844
rect 3724 34790 3726 34842
rect 3906 34790 3908 34842
rect 3662 34788 3668 34790
rect 3724 34788 3748 34790
rect 3804 34788 3828 34790
rect 3884 34788 3908 34790
rect 3964 34788 3970 34790
rect 3662 34779 3970 34788
rect 9128 34536 9180 34542
rect 9128 34478 9180 34484
rect 8852 34468 8904 34474
rect 8852 34410 8904 34416
rect 4322 34300 4630 34309
rect 4322 34298 4328 34300
rect 4384 34298 4408 34300
rect 4464 34298 4488 34300
rect 4544 34298 4568 34300
rect 4624 34298 4630 34300
rect 4384 34246 4386 34298
rect 4566 34246 4568 34298
rect 4322 34244 4328 34246
rect 4384 34244 4408 34246
rect 4464 34244 4488 34246
rect 4544 34244 4568 34246
rect 4624 34244 4630 34246
rect 4322 34235 4630 34244
rect 8864 34202 8892 34410
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 3662 33756 3970 33765
rect 3662 33754 3668 33756
rect 3724 33754 3748 33756
rect 3804 33754 3828 33756
rect 3884 33754 3908 33756
rect 3964 33754 3970 33756
rect 3724 33702 3726 33754
rect 3906 33702 3908 33754
rect 3662 33700 3668 33702
rect 3724 33700 3748 33702
rect 3804 33700 3828 33702
rect 3884 33700 3908 33702
rect 3964 33700 3970 33702
rect 3662 33691 3970 33700
rect 4322 33212 4630 33221
rect 4322 33210 4328 33212
rect 4384 33210 4408 33212
rect 4464 33210 4488 33212
rect 4544 33210 4568 33212
rect 4624 33210 4630 33212
rect 4384 33158 4386 33210
rect 4566 33158 4568 33210
rect 4322 33156 4328 33158
rect 4384 33156 4408 33158
rect 4464 33156 4488 33158
rect 4544 33156 4568 33158
rect 4624 33156 4630 33158
rect 4322 33147 4630 33156
rect 8852 32972 8904 32978
rect 8852 32914 8904 32920
rect 3662 32668 3970 32677
rect 3662 32666 3668 32668
rect 3724 32666 3748 32668
rect 3804 32666 3828 32668
rect 3884 32666 3908 32668
rect 3964 32666 3970 32668
rect 3724 32614 3726 32666
rect 3906 32614 3908 32666
rect 3662 32612 3668 32614
rect 3724 32612 3748 32614
rect 3804 32612 3828 32614
rect 3884 32612 3908 32614
rect 3964 32612 3970 32614
rect 3662 32603 3970 32612
rect 8864 32570 8892 32914
rect 8852 32564 8904 32570
rect 8852 32506 8904 32512
rect 4322 32124 4630 32133
rect 4322 32122 4328 32124
rect 4384 32122 4408 32124
rect 4464 32122 4488 32124
rect 4544 32122 4568 32124
rect 4624 32122 4630 32124
rect 4384 32070 4386 32122
rect 4566 32070 4568 32122
rect 4322 32068 4328 32070
rect 4384 32068 4408 32070
rect 4464 32068 4488 32070
rect 4544 32068 4568 32070
rect 4624 32068 4630 32070
rect 4322 32059 4630 32068
rect 9140 31890 9168 34478
rect 9312 34400 9364 34406
rect 9312 34342 9364 34348
rect 9324 34066 9352 34342
rect 9508 34202 9536 35566
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 9496 34196 9548 34202
rect 9496 34138 9548 34144
rect 9220 34060 9272 34066
rect 9220 34002 9272 34008
rect 9312 34060 9364 34066
rect 9312 34002 9364 34008
rect 9232 33946 9260 34002
rect 9692 33998 9720 34682
rect 9784 34066 9812 35022
rect 9772 34060 9824 34066
rect 9824 34020 9904 34048
rect 9772 34002 9824 34008
rect 9680 33992 9732 33998
rect 9232 33930 9352 33946
rect 9680 33934 9732 33940
rect 9232 33924 9364 33930
rect 9232 33918 9312 33924
rect 9312 33866 9364 33872
rect 9220 32972 9272 32978
rect 9220 32914 9272 32920
rect 9232 32502 9260 32914
rect 9220 32496 9272 32502
rect 9220 32438 9272 32444
rect 9128 31884 9180 31890
rect 9128 31826 9180 31832
rect 9140 31754 9168 31826
rect 9048 31726 9168 31754
rect 8852 31680 8904 31686
rect 8852 31622 8904 31628
rect 3662 31580 3970 31589
rect 3662 31578 3668 31580
rect 3724 31578 3748 31580
rect 3804 31578 3828 31580
rect 3884 31578 3908 31580
rect 3964 31578 3970 31580
rect 3724 31526 3726 31578
rect 3906 31526 3908 31578
rect 3662 31524 3668 31526
rect 3724 31524 3748 31526
rect 3804 31524 3828 31526
rect 3884 31524 3908 31526
rect 3964 31524 3970 31526
rect 3662 31515 3970 31524
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 4322 31036 4630 31045
rect 4322 31034 4328 31036
rect 4384 31034 4408 31036
rect 4464 31034 4488 31036
rect 4544 31034 4568 31036
rect 4624 31034 4630 31036
rect 4384 30982 4386 31034
rect 4566 30982 4568 31034
rect 4322 30980 4328 30982
rect 4384 30980 4408 30982
rect 4464 30980 4488 30982
rect 4544 30980 4568 30982
rect 4624 30980 4630 30982
rect 4322 30971 4630 30980
rect 8680 30870 8708 31078
rect 8668 30864 8720 30870
rect 8668 30806 8720 30812
rect 8864 30802 8892 31622
rect 8944 31272 8996 31278
rect 8944 31214 8996 31220
rect 8956 30938 8984 31214
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 8852 30796 8904 30802
rect 8852 30738 8904 30744
rect 3662 30492 3970 30501
rect 3662 30490 3668 30492
rect 3724 30490 3748 30492
rect 3804 30490 3828 30492
rect 3884 30490 3908 30492
rect 3964 30490 3970 30492
rect 3724 30438 3726 30490
rect 3906 30438 3908 30490
rect 3662 30436 3668 30438
rect 3724 30436 3748 30438
rect 3804 30436 3828 30438
rect 3884 30436 3908 30438
rect 3964 30436 3970 30438
rect 3662 30427 3970 30436
rect 9048 30190 9076 31726
rect 9324 31686 9352 33866
rect 9692 32994 9720 33934
rect 9876 33522 9904 34020
rect 9864 33516 9916 33522
rect 9864 33458 9916 33464
rect 9968 33402 9996 35652
rect 10060 35154 10088 35770
rect 10152 35630 10180 36858
rect 10244 36242 10272 38218
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 10336 37874 10364 38150
rect 10324 37868 10376 37874
rect 10324 37810 10376 37816
rect 10428 37466 10456 39238
rect 10520 38350 10548 41386
rect 10796 41138 10824 41618
rect 10600 41132 10652 41138
rect 10600 41074 10652 41080
rect 10784 41132 10836 41138
rect 10784 41074 10836 41080
rect 10612 39982 10640 41074
rect 11072 41070 11100 42706
rect 11256 41414 11284 43794
rect 11348 43450 11376 43823
rect 11436 43548 11744 43557
rect 11436 43546 11442 43548
rect 11498 43546 11522 43548
rect 11578 43546 11602 43548
rect 11658 43546 11682 43548
rect 11738 43546 11744 43548
rect 11498 43494 11500 43546
rect 11680 43494 11682 43546
rect 11436 43492 11442 43494
rect 11498 43492 11522 43494
rect 11578 43492 11602 43494
rect 11658 43492 11682 43494
rect 11738 43492 11744 43494
rect 11436 43483 11744 43492
rect 11336 43444 11388 43450
rect 11336 43386 11388 43392
rect 11900 43110 11928 44338
rect 21652 44334 21680 44775
rect 24030 44704 24086 44713
rect 24030 44639 24086 44648
rect 24398 44704 24454 44713
rect 24398 44639 24454 44648
rect 24950 44704 25006 44713
rect 24950 44639 25006 44648
rect 25502 44704 25558 44713
rect 25502 44639 25558 44648
rect 26054 44704 26110 44713
rect 26054 44639 26110 44648
rect 26514 44704 26570 44713
rect 26514 44639 26570 44648
rect 24044 44334 24072 44639
rect 24412 44334 24440 44639
rect 24964 44334 24992 44639
rect 25228 44464 25280 44470
rect 25228 44406 25280 44412
rect 13728 44328 13780 44334
rect 13728 44270 13780 44276
rect 13820 44328 13872 44334
rect 13820 44270 13872 44276
rect 14004 44328 14056 44334
rect 15844 44328 15896 44334
rect 14056 44276 14504 44282
rect 14004 44270 14504 44276
rect 15844 44270 15896 44276
rect 16488 44328 16540 44334
rect 16488 44270 16540 44276
rect 21640 44328 21692 44334
rect 21640 44270 21692 44276
rect 24032 44328 24084 44334
rect 24032 44270 24084 44276
rect 24400 44328 24452 44334
rect 24400 44270 24452 44276
rect 24952 44328 25004 44334
rect 24952 44270 25004 44276
rect 12440 44192 12492 44198
rect 12440 44134 12492 44140
rect 12532 44192 12584 44198
rect 12532 44134 12584 44140
rect 13544 44192 13596 44198
rect 13544 44134 13596 44140
rect 12096 44092 12404 44101
rect 12096 44090 12102 44092
rect 12158 44090 12182 44092
rect 12238 44090 12262 44092
rect 12318 44090 12342 44092
rect 12398 44090 12404 44092
rect 12158 44038 12160 44090
rect 12340 44038 12342 44090
rect 12096 44036 12102 44038
rect 12158 44036 12182 44038
rect 12238 44036 12262 44038
rect 12318 44036 12342 44038
rect 12398 44036 12404 44038
rect 12096 44027 12404 44036
rect 12348 43852 12400 43858
rect 12452 43840 12480 44134
rect 12400 43812 12480 43840
rect 12348 43794 12400 43800
rect 11980 43240 12032 43246
rect 11980 43182 12032 43188
rect 11888 43104 11940 43110
rect 11888 43046 11940 43052
rect 11336 42696 11388 42702
rect 11336 42638 11388 42644
rect 11164 41386 11284 41414
rect 10968 41064 11020 41070
rect 10968 41006 11020 41012
rect 11060 41064 11112 41070
rect 11060 41006 11112 41012
rect 10980 40730 11008 41006
rect 10968 40724 11020 40730
rect 10968 40666 11020 40672
rect 10692 40520 10744 40526
rect 10692 40462 10744 40468
rect 10704 40390 10732 40462
rect 10968 40452 11020 40458
rect 10968 40394 11020 40400
rect 10692 40384 10744 40390
rect 10692 40326 10744 40332
rect 10980 40118 11008 40394
rect 10968 40112 11020 40118
rect 10968 40054 11020 40060
rect 10600 39976 10652 39982
rect 10600 39918 10652 39924
rect 10692 39976 10744 39982
rect 10692 39918 10744 39924
rect 10876 39976 10928 39982
rect 10876 39918 10928 39924
rect 10966 39944 11022 39953
rect 10612 39098 10640 39918
rect 10704 39642 10732 39918
rect 10692 39636 10744 39642
rect 10692 39578 10744 39584
rect 10888 39098 10916 39918
rect 10966 39879 11022 39888
rect 10980 39574 11008 39879
rect 10968 39568 11020 39574
rect 10968 39510 11020 39516
rect 10600 39092 10652 39098
rect 10600 39034 10652 39040
rect 10876 39092 10928 39098
rect 10876 39034 10928 39040
rect 10508 38344 10560 38350
rect 10508 38286 10560 38292
rect 10612 37670 10640 39034
rect 10968 38956 11020 38962
rect 10968 38898 11020 38904
rect 10980 38350 11008 38898
rect 10968 38344 11020 38350
rect 10968 38286 11020 38292
rect 10876 37800 10928 37806
rect 10876 37742 10928 37748
rect 10600 37664 10652 37670
rect 10600 37606 10652 37612
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10888 37398 10916 37742
rect 10876 37392 10928 37398
rect 10876 37334 10928 37340
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 10416 37324 10468 37330
rect 10416 37266 10468 37272
rect 10232 36236 10284 36242
rect 10232 36178 10284 36184
rect 10140 35624 10192 35630
rect 10336 35578 10364 37266
rect 10428 36650 10456 37266
rect 10692 37120 10744 37126
rect 10692 37062 10744 37068
rect 10416 36644 10468 36650
rect 10416 36586 10468 36592
rect 10140 35566 10192 35572
rect 10152 35290 10180 35566
rect 10244 35550 10364 35578
rect 10140 35284 10192 35290
rect 10140 35226 10192 35232
rect 10048 35148 10100 35154
rect 10100 35108 10180 35136
rect 10048 35090 10100 35096
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 10060 34542 10088 34886
rect 10048 34536 10100 34542
rect 10048 34478 10100 34484
rect 9968 33386 10088 33402
rect 9864 33380 9916 33386
rect 9968 33380 10100 33386
rect 9968 33374 10048 33380
rect 9864 33322 9916 33328
rect 10048 33322 10100 33328
rect 9600 32978 9720 32994
rect 9588 32972 9720 32978
rect 9640 32966 9720 32972
rect 9588 32914 9640 32920
rect 9404 32768 9456 32774
rect 9404 32710 9456 32716
rect 9312 31680 9364 31686
rect 9312 31622 9364 31628
rect 9324 31414 9352 31622
rect 9312 31408 9364 31414
rect 9312 31350 9364 31356
rect 9416 31346 9444 32710
rect 9692 32366 9720 32966
rect 9876 32570 9904 33322
rect 9956 33312 10008 33318
rect 9956 33254 10008 33260
rect 9968 32978 9996 33254
rect 10060 33046 10088 33322
rect 10152 33046 10180 35108
rect 10244 34134 10272 35550
rect 10324 35488 10376 35494
rect 10324 35430 10376 35436
rect 10336 34406 10364 35430
rect 10428 34746 10456 36586
rect 10704 36242 10732 37062
rect 11060 36644 11112 36650
rect 11060 36586 11112 36592
rect 10968 36576 11020 36582
rect 10968 36518 11020 36524
rect 10980 36310 11008 36518
rect 10968 36304 11020 36310
rect 10968 36246 11020 36252
rect 10508 36236 10560 36242
rect 10508 36178 10560 36184
rect 10692 36236 10744 36242
rect 10692 36178 10744 36184
rect 10520 35562 10548 36178
rect 10508 35556 10560 35562
rect 10508 35498 10560 35504
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10324 34400 10376 34406
rect 10324 34342 10376 34348
rect 10232 34128 10284 34134
rect 10232 34070 10284 34076
rect 10244 33454 10272 34070
rect 10520 33590 10548 35498
rect 11072 34542 11100 36586
rect 11060 34536 11112 34542
rect 11060 34478 11112 34484
rect 10508 33584 10560 33590
rect 10508 33526 10560 33532
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10232 33448 10284 33454
rect 10232 33390 10284 33396
rect 10048 33040 10100 33046
rect 10048 32982 10100 32988
rect 10140 33040 10192 33046
rect 10140 32982 10192 32988
rect 9956 32972 10008 32978
rect 9956 32914 10008 32920
rect 9864 32564 9916 32570
rect 9864 32506 9916 32512
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9876 32230 9904 32506
rect 10152 32434 10180 32982
rect 10140 32428 10192 32434
rect 10140 32370 10192 32376
rect 10048 32292 10100 32298
rect 10048 32234 10100 32240
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 9864 32224 9916 32230
rect 9864 32166 9916 32172
rect 9956 32224 10008 32230
rect 9956 32166 10008 32172
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9692 31278 9720 32166
rect 9968 31278 9996 32166
rect 9680 31272 9732 31278
rect 9680 31214 9732 31220
rect 9956 31272 10008 31278
rect 9956 31214 10008 31220
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 9600 30122 9628 31078
rect 9692 30394 9720 31214
rect 10060 30802 10088 32234
rect 10244 31958 10272 33390
rect 10428 33114 10456 33458
rect 10416 33108 10468 33114
rect 10336 33068 10416 33096
rect 10232 31952 10284 31958
rect 10232 31894 10284 31900
rect 10336 30938 10364 33068
rect 10416 33050 10468 33056
rect 10520 32910 10548 33526
rect 10968 33448 11020 33454
rect 10968 33390 11020 33396
rect 10692 33312 10744 33318
rect 10692 33254 10744 33260
rect 10508 32904 10560 32910
rect 10508 32846 10560 32852
rect 10416 32768 10468 32774
rect 10416 32710 10468 32716
rect 10508 32768 10560 32774
rect 10508 32710 10560 32716
rect 10428 32366 10456 32710
rect 10520 32366 10548 32710
rect 10704 32366 10732 33254
rect 10876 33040 10928 33046
rect 10876 32982 10928 32988
rect 10784 32972 10836 32978
rect 10784 32914 10836 32920
rect 10796 32570 10824 32914
rect 10784 32564 10836 32570
rect 10784 32506 10836 32512
rect 10416 32360 10468 32366
rect 10416 32302 10468 32308
rect 10508 32360 10560 32366
rect 10508 32302 10560 32308
rect 10692 32360 10744 32366
rect 10692 32302 10744 32308
rect 10888 31958 10916 32982
rect 10980 32026 11008 33390
rect 11060 33312 11112 33318
rect 11060 33254 11112 33260
rect 11072 32366 11100 33254
rect 11060 32360 11112 32366
rect 11060 32302 11112 32308
rect 10968 32020 11020 32026
rect 10968 31962 11020 31968
rect 10876 31952 10928 31958
rect 10876 31894 10928 31900
rect 11060 31680 11112 31686
rect 11060 31622 11112 31628
rect 11072 31278 11100 31622
rect 11164 31482 11192 41386
rect 11348 40050 11376 42638
rect 11436 42460 11744 42469
rect 11436 42458 11442 42460
rect 11498 42458 11522 42460
rect 11578 42458 11602 42460
rect 11658 42458 11682 42460
rect 11738 42458 11744 42460
rect 11498 42406 11500 42458
rect 11680 42406 11682 42458
rect 11436 42404 11442 42406
rect 11498 42404 11522 42406
rect 11578 42404 11602 42406
rect 11658 42404 11682 42406
rect 11738 42404 11744 42406
rect 11436 42395 11744 42404
rect 11436 41372 11744 41381
rect 11436 41370 11442 41372
rect 11498 41370 11522 41372
rect 11578 41370 11602 41372
rect 11658 41370 11682 41372
rect 11738 41370 11744 41372
rect 11498 41318 11500 41370
rect 11680 41318 11682 41370
rect 11436 41316 11442 41318
rect 11498 41316 11522 41318
rect 11578 41316 11602 41318
rect 11658 41316 11682 41318
rect 11738 41316 11744 41318
rect 11436 41307 11744 41316
rect 11796 40996 11848 41002
rect 11796 40938 11848 40944
rect 11808 40730 11836 40938
rect 11796 40724 11848 40730
rect 11796 40666 11848 40672
rect 11796 40452 11848 40458
rect 11796 40394 11848 40400
rect 11436 40284 11744 40293
rect 11436 40282 11442 40284
rect 11498 40282 11522 40284
rect 11578 40282 11602 40284
rect 11658 40282 11682 40284
rect 11738 40282 11744 40284
rect 11498 40230 11500 40282
rect 11680 40230 11682 40282
rect 11436 40228 11442 40230
rect 11498 40228 11522 40230
rect 11578 40228 11602 40230
rect 11658 40228 11682 40230
rect 11738 40228 11744 40230
rect 11436 40219 11744 40228
rect 11808 40168 11836 40394
rect 11716 40140 11836 40168
rect 11336 40044 11388 40050
rect 11336 39986 11388 39992
rect 11336 39908 11388 39914
rect 11336 39850 11388 39856
rect 11348 39438 11376 39850
rect 11612 39840 11664 39846
rect 11612 39782 11664 39788
rect 11624 39642 11652 39782
rect 11612 39636 11664 39642
rect 11612 39578 11664 39584
rect 11716 39506 11744 40140
rect 11900 39930 11928 43046
rect 11992 42906 12020 43182
rect 12096 43004 12404 43013
rect 12096 43002 12102 43004
rect 12158 43002 12182 43004
rect 12238 43002 12262 43004
rect 12318 43002 12342 43004
rect 12398 43002 12404 43004
rect 12158 42950 12160 43002
rect 12340 42950 12342 43002
rect 12096 42948 12102 42950
rect 12158 42948 12182 42950
rect 12238 42948 12262 42950
rect 12318 42948 12342 42950
rect 12398 42948 12404 42950
rect 12096 42939 12404 42948
rect 11980 42900 12032 42906
rect 11980 42842 12032 42848
rect 12544 42770 12572 44134
rect 13266 44024 13322 44033
rect 13266 43959 13268 43968
rect 13320 43959 13322 43968
rect 13268 43930 13320 43936
rect 13556 43246 13584 44134
rect 13544 43240 13596 43246
rect 13544 43182 13596 43188
rect 12532 42764 12584 42770
rect 12532 42706 12584 42712
rect 13544 42764 13596 42770
rect 13544 42706 13596 42712
rect 13556 42362 13584 42706
rect 13740 42378 13768 44270
rect 13832 43994 13860 44270
rect 14016 44254 14504 44270
rect 14280 44192 14332 44198
rect 14280 44134 14332 44140
rect 13820 43988 13872 43994
rect 13820 43930 13872 43936
rect 14292 43858 14320 44134
rect 14004 43852 14056 43858
rect 14004 43794 14056 43800
rect 14280 43852 14332 43858
rect 14280 43794 14332 43800
rect 13818 43752 13874 43761
rect 13818 43687 13874 43696
rect 13832 43654 13860 43687
rect 13820 43648 13872 43654
rect 13820 43590 13872 43596
rect 14016 43246 14044 43794
rect 14188 43784 14240 43790
rect 14188 43726 14240 43732
rect 14200 43382 14228 43726
rect 14370 43480 14426 43489
rect 14370 43415 14372 43424
rect 14424 43415 14426 43424
rect 14372 43386 14424 43392
rect 14188 43376 14240 43382
rect 14188 43318 14240 43324
rect 14200 43246 14228 43318
rect 14004 43240 14056 43246
rect 14004 43182 14056 43188
rect 14188 43240 14240 43246
rect 14188 43182 14240 43188
rect 14016 42906 14044 43182
rect 14188 43104 14240 43110
rect 14188 43046 14240 43052
rect 14004 42900 14056 42906
rect 14004 42842 14056 42848
rect 13544 42356 13596 42362
rect 13740 42350 13860 42378
rect 13544 42298 13596 42304
rect 13728 42152 13780 42158
rect 13728 42094 13780 42100
rect 12096 41916 12404 41925
rect 12096 41914 12102 41916
rect 12158 41914 12182 41916
rect 12238 41914 12262 41916
rect 12318 41914 12342 41916
rect 12398 41914 12404 41916
rect 12158 41862 12160 41914
rect 12340 41862 12342 41914
rect 12096 41860 12102 41862
rect 12158 41860 12182 41862
rect 12238 41860 12262 41862
rect 12318 41860 12342 41862
rect 12398 41860 12404 41862
rect 12096 41851 12404 41860
rect 13740 41857 13768 42094
rect 13726 41848 13782 41857
rect 13832 41818 13860 42350
rect 14200 42158 14228 43046
rect 14280 42696 14332 42702
rect 14280 42638 14332 42644
rect 14292 42362 14320 42638
rect 14280 42356 14332 42362
rect 14280 42298 14332 42304
rect 14004 42152 14056 42158
rect 14004 42094 14056 42100
rect 14188 42152 14240 42158
rect 14188 42094 14240 42100
rect 13726 41783 13782 41792
rect 13820 41812 13872 41818
rect 13820 41754 13872 41760
rect 14016 41682 14044 42094
rect 14280 41812 14332 41818
rect 14280 41754 14332 41760
rect 14004 41676 14056 41682
rect 14004 41618 14056 41624
rect 12716 41608 12768 41614
rect 12716 41550 12768 41556
rect 12440 41472 12492 41478
rect 12440 41414 12492 41420
rect 12096 40828 12404 40837
rect 12096 40826 12102 40828
rect 12158 40826 12182 40828
rect 12238 40826 12262 40828
rect 12318 40826 12342 40828
rect 12398 40826 12404 40828
rect 12158 40774 12160 40826
rect 12340 40774 12342 40826
rect 12096 40772 12102 40774
rect 12158 40772 12182 40774
rect 12238 40772 12262 40774
rect 12318 40772 12342 40774
rect 12398 40772 12404 40774
rect 12096 40763 12404 40772
rect 12452 40730 12480 41414
rect 12624 41268 12676 41274
rect 12624 41210 12676 41216
rect 12532 40928 12584 40934
rect 12532 40870 12584 40876
rect 12440 40724 12492 40730
rect 12440 40666 12492 40672
rect 11980 40656 12032 40662
rect 11980 40598 12032 40604
rect 11808 39902 11928 39930
rect 11704 39500 11756 39506
rect 11704 39442 11756 39448
rect 11336 39432 11388 39438
rect 11336 39374 11388 39380
rect 11348 38486 11376 39374
rect 11436 39196 11744 39205
rect 11436 39194 11442 39196
rect 11498 39194 11522 39196
rect 11578 39194 11602 39196
rect 11658 39194 11682 39196
rect 11738 39194 11744 39196
rect 11498 39142 11500 39194
rect 11680 39142 11682 39194
rect 11436 39140 11442 39142
rect 11498 39140 11522 39142
rect 11578 39140 11602 39142
rect 11658 39140 11682 39142
rect 11738 39140 11744 39142
rect 11436 39131 11744 39140
rect 11336 38480 11388 38486
rect 11336 38422 11388 38428
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 11256 37806 11284 38150
rect 11244 37800 11296 37806
rect 11244 37742 11296 37748
rect 11348 36802 11376 38422
rect 11436 38108 11744 38117
rect 11436 38106 11442 38108
rect 11498 38106 11522 38108
rect 11578 38106 11602 38108
rect 11658 38106 11682 38108
rect 11738 38106 11744 38108
rect 11498 38054 11500 38106
rect 11680 38054 11682 38106
rect 11436 38052 11442 38054
rect 11498 38052 11522 38054
rect 11578 38052 11602 38054
rect 11658 38052 11682 38054
rect 11738 38052 11744 38054
rect 11436 38043 11744 38052
rect 11436 37020 11744 37029
rect 11436 37018 11442 37020
rect 11498 37018 11522 37020
rect 11578 37018 11602 37020
rect 11658 37018 11682 37020
rect 11738 37018 11744 37020
rect 11498 36966 11500 37018
rect 11680 36966 11682 37018
rect 11436 36964 11442 36966
rect 11498 36964 11522 36966
rect 11578 36964 11602 36966
rect 11658 36964 11682 36966
rect 11738 36964 11744 36966
rect 11436 36955 11744 36964
rect 11348 36774 11560 36802
rect 11244 36712 11296 36718
rect 11244 36654 11296 36660
rect 11428 36712 11480 36718
rect 11428 36654 11480 36660
rect 11256 36310 11284 36654
rect 11440 36378 11468 36654
rect 11428 36372 11480 36378
rect 11428 36314 11480 36320
rect 11244 36304 11296 36310
rect 11244 36246 11296 36252
rect 11532 36174 11560 36774
rect 11244 36168 11296 36174
rect 11244 36110 11296 36116
rect 11520 36168 11572 36174
rect 11520 36110 11572 36116
rect 11256 35086 11284 36110
rect 11436 35932 11744 35941
rect 11436 35930 11442 35932
rect 11498 35930 11522 35932
rect 11578 35930 11602 35932
rect 11658 35930 11682 35932
rect 11738 35930 11744 35932
rect 11498 35878 11500 35930
rect 11680 35878 11682 35930
rect 11436 35876 11442 35878
rect 11498 35876 11522 35878
rect 11578 35876 11602 35878
rect 11658 35876 11682 35878
rect 11738 35876 11744 35878
rect 11436 35867 11744 35876
rect 11520 35556 11572 35562
rect 11520 35498 11572 35504
rect 11704 35556 11756 35562
rect 11704 35498 11756 35504
rect 11532 35290 11560 35498
rect 11612 35488 11664 35494
rect 11612 35430 11664 35436
rect 11520 35284 11572 35290
rect 11520 35226 11572 35232
rect 11624 35154 11652 35430
rect 11612 35148 11664 35154
rect 11612 35090 11664 35096
rect 11244 35080 11296 35086
rect 11244 35022 11296 35028
rect 11256 33930 11284 35022
rect 11716 34950 11744 35498
rect 11808 35034 11836 39902
rect 11888 39840 11940 39846
rect 11888 39782 11940 39788
rect 11900 39506 11928 39782
rect 11992 39574 12020 40598
rect 12544 40594 12572 40870
rect 12164 40588 12216 40594
rect 12164 40530 12216 40536
rect 12256 40588 12308 40594
rect 12256 40530 12308 40536
rect 12532 40588 12584 40594
rect 12532 40530 12584 40536
rect 12176 39914 12204 40530
rect 12268 40186 12296 40530
rect 12636 40474 12664 41210
rect 12728 40934 12756 41550
rect 12808 40996 12860 41002
rect 12808 40938 12860 40944
rect 13084 40996 13136 41002
rect 13084 40938 13136 40944
rect 12716 40928 12768 40934
rect 12716 40870 12768 40876
rect 12728 40662 12756 40870
rect 12716 40656 12768 40662
rect 12716 40598 12768 40604
rect 12452 40446 12664 40474
rect 12256 40180 12308 40186
rect 12256 40122 12308 40128
rect 12164 39908 12216 39914
rect 12164 39850 12216 39856
rect 12096 39740 12404 39749
rect 12096 39738 12102 39740
rect 12158 39738 12182 39740
rect 12238 39738 12262 39740
rect 12318 39738 12342 39740
rect 12398 39738 12404 39740
rect 12158 39686 12160 39738
rect 12340 39686 12342 39738
rect 12096 39684 12102 39686
rect 12158 39684 12182 39686
rect 12238 39684 12262 39686
rect 12318 39684 12342 39686
rect 12398 39684 12404 39686
rect 12096 39675 12404 39684
rect 12452 39642 12480 40446
rect 12624 40384 12676 40390
rect 12624 40326 12676 40332
rect 12532 39840 12584 39846
rect 12532 39782 12584 39788
rect 12440 39636 12492 39642
rect 12440 39578 12492 39584
rect 12544 39574 12572 39782
rect 11980 39568 12032 39574
rect 11980 39510 12032 39516
rect 12532 39568 12584 39574
rect 12532 39510 12584 39516
rect 11888 39500 11940 39506
rect 11888 39442 11940 39448
rect 11888 39296 11940 39302
rect 11888 39238 11940 39244
rect 11900 38486 11928 39238
rect 11888 38480 11940 38486
rect 11888 38422 11940 38428
rect 11992 38298 12020 39510
rect 12636 39506 12664 40326
rect 12716 39908 12768 39914
rect 12820 39896 12848 40938
rect 12900 40588 12952 40594
rect 12900 40530 12952 40536
rect 12992 40588 13044 40594
rect 12992 40530 13044 40536
rect 12768 39868 12848 39896
rect 12716 39850 12768 39856
rect 12624 39500 12676 39506
rect 12624 39442 12676 39448
rect 12532 39432 12584 39438
rect 12532 39374 12584 39380
rect 12440 39296 12492 39302
rect 12440 39238 12492 39244
rect 12452 38894 12480 39238
rect 12544 39098 12572 39374
rect 12624 39364 12676 39370
rect 12624 39306 12676 39312
rect 12532 39092 12584 39098
rect 12532 39034 12584 39040
rect 12440 38888 12492 38894
rect 12440 38830 12492 38836
rect 12096 38652 12404 38661
rect 12096 38650 12102 38652
rect 12158 38650 12182 38652
rect 12238 38650 12262 38652
rect 12318 38650 12342 38652
rect 12398 38650 12404 38652
rect 12158 38598 12160 38650
rect 12340 38598 12342 38650
rect 12096 38596 12102 38598
rect 12158 38596 12182 38598
rect 12238 38596 12262 38598
rect 12318 38596 12342 38598
rect 12398 38596 12404 38598
rect 12096 38587 12404 38596
rect 12452 38418 12480 38830
rect 12440 38412 12492 38418
rect 12440 38354 12492 38360
rect 11900 38270 12020 38298
rect 11900 36174 11928 38270
rect 12452 38010 12480 38354
rect 12440 38004 12492 38010
rect 12440 37946 12492 37952
rect 12096 37564 12404 37573
rect 12096 37562 12102 37564
rect 12158 37562 12182 37564
rect 12238 37562 12262 37564
rect 12318 37562 12342 37564
rect 12398 37562 12404 37564
rect 12158 37510 12160 37562
rect 12340 37510 12342 37562
rect 12096 37508 12102 37510
rect 12158 37508 12182 37510
rect 12238 37508 12262 37510
rect 12318 37508 12342 37510
rect 12398 37508 12404 37510
rect 12096 37499 12404 37508
rect 12636 36718 12664 39306
rect 12728 38826 12756 39850
rect 12912 39846 12940 40530
rect 13004 39953 13032 40530
rect 13096 40050 13124 40938
rect 13268 40928 13320 40934
rect 13268 40870 13320 40876
rect 14096 40928 14148 40934
rect 14096 40870 14148 40876
rect 13280 40594 13308 40870
rect 14108 40594 14136 40870
rect 13268 40588 13320 40594
rect 13268 40530 13320 40536
rect 14096 40588 14148 40594
rect 14096 40530 14148 40536
rect 14096 40452 14148 40458
rect 14096 40394 14148 40400
rect 13268 40112 13320 40118
rect 13268 40054 13320 40060
rect 13084 40044 13136 40050
rect 13084 39986 13136 39992
rect 12990 39944 13046 39953
rect 13046 39902 13216 39930
rect 12990 39879 13046 39888
rect 12900 39840 12952 39846
rect 12900 39782 12952 39788
rect 12992 39500 13044 39506
rect 12992 39442 13044 39448
rect 12808 39092 12860 39098
rect 12808 39034 12860 39040
rect 12716 38820 12768 38826
rect 12716 38762 12768 38768
rect 12716 38208 12768 38214
rect 12716 38150 12768 38156
rect 12728 37806 12756 38150
rect 12820 37806 12848 39034
rect 12900 38820 12952 38826
rect 12900 38762 12952 38768
rect 12912 37942 12940 38762
rect 13004 38400 13032 39442
rect 13004 38372 13124 38400
rect 12992 38276 13044 38282
rect 12992 38218 13044 38224
rect 12900 37936 12952 37942
rect 12900 37878 12952 37884
rect 12716 37800 12768 37806
rect 12716 37742 12768 37748
rect 12808 37800 12860 37806
rect 12808 37742 12860 37748
rect 12912 37618 12940 37878
rect 13004 37806 13032 38218
rect 13096 38010 13124 38372
rect 13084 38004 13136 38010
rect 13084 37946 13136 37952
rect 12992 37800 13044 37806
rect 12992 37742 13044 37748
rect 12912 37590 13032 37618
rect 12900 36916 12952 36922
rect 12900 36858 12952 36864
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12096 36476 12404 36485
rect 12096 36474 12102 36476
rect 12158 36474 12182 36476
rect 12238 36474 12262 36476
rect 12318 36474 12342 36476
rect 12398 36474 12404 36476
rect 12158 36422 12160 36474
rect 12340 36422 12342 36474
rect 12096 36420 12102 36422
rect 12158 36420 12182 36422
rect 12238 36420 12262 36422
rect 12318 36420 12342 36422
rect 12398 36420 12404 36422
rect 12096 36411 12404 36420
rect 12636 36242 12664 36654
rect 12912 36242 12940 36858
rect 13004 36582 13032 37590
rect 12992 36576 13044 36582
rect 12992 36518 13044 36524
rect 11980 36236 12032 36242
rect 11980 36178 12032 36184
rect 12164 36236 12216 36242
rect 12624 36236 12676 36242
rect 12216 36196 12296 36224
rect 12164 36178 12216 36184
rect 11888 36168 11940 36174
rect 11888 36110 11940 36116
rect 11888 36032 11940 36038
rect 11888 35974 11940 35980
rect 11900 35154 11928 35974
rect 11992 35290 12020 36178
rect 12268 35766 12296 36196
rect 12624 36178 12676 36184
rect 12808 36236 12860 36242
rect 12808 36178 12860 36184
rect 12900 36236 12952 36242
rect 12900 36178 12952 36184
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12636 35834 12664 35974
rect 12728 35834 12756 36110
rect 12820 35834 12848 36178
rect 12624 35828 12676 35834
rect 12624 35770 12676 35776
rect 12716 35828 12768 35834
rect 12716 35770 12768 35776
rect 12808 35828 12860 35834
rect 12808 35770 12860 35776
rect 12256 35760 12308 35766
rect 12256 35702 12308 35708
rect 12268 35578 12296 35702
rect 12268 35550 12480 35578
rect 12096 35388 12404 35397
rect 12096 35386 12102 35388
rect 12158 35386 12182 35388
rect 12238 35386 12262 35388
rect 12318 35386 12342 35388
rect 12398 35386 12404 35388
rect 12158 35334 12160 35386
rect 12340 35334 12342 35386
rect 12096 35332 12102 35334
rect 12158 35332 12182 35334
rect 12238 35332 12262 35334
rect 12318 35332 12342 35334
rect 12398 35332 12404 35334
rect 12096 35323 12404 35332
rect 11980 35284 12032 35290
rect 11980 35226 12032 35232
rect 11888 35148 11940 35154
rect 11888 35090 11940 35096
rect 12072 35148 12124 35154
rect 12072 35090 12124 35096
rect 12164 35148 12216 35154
rect 12164 35090 12216 35096
rect 11808 35006 12020 35034
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11888 34944 11940 34950
rect 11888 34886 11940 34892
rect 11436 34844 11744 34853
rect 11436 34842 11442 34844
rect 11498 34842 11522 34844
rect 11578 34842 11602 34844
rect 11658 34842 11682 34844
rect 11738 34842 11744 34844
rect 11498 34790 11500 34842
rect 11680 34790 11682 34842
rect 11436 34788 11442 34790
rect 11498 34788 11522 34790
rect 11578 34788 11602 34790
rect 11658 34788 11682 34790
rect 11738 34788 11744 34790
rect 11436 34779 11744 34788
rect 11796 34740 11848 34746
rect 11796 34682 11848 34688
rect 11808 34202 11836 34682
rect 11336 34196 11388 34202
rect 11336 34138 11388 34144
rect 11796 34196 11848 34202
rect 11796 34138 11848 34144
rect 11244 33924 11296 33930
rect 11244 33866 11296 33872
rect 11348 33538 11376 34138
rect 11900 34066 11928 34886
rect 11888 34060 11940 34066
rect 11888 34002 11940 34008
rect 11796 33856 11848 33862
rect 11796 33798 11848 33804
rect 11436 33756 11744 33765
rect 11436 33754 11442 33756
rect 11498 33754 11522 33756
rect 11578 33754 11602 33756
rect 11658 33754 11682 33756
rect 11738 33754 11744 33756
rect 11498 33702 11500 33754
rect 11680 33702 11682 33754
rect 11436 33700 11442 33702
rect 11498 33700 11522 33702
rect 11578 33700 11602 33702
rect 11658 33700 11682 33702
rect 11738 33700 11744 33702
rect 11436 33691 11744 33700
rect 11348 33510 11468 33538
rect 11808 33522 11836 33798
rect 11336 33448 11388 33454
rect 11336 33390 11388 33396
rect 11348 32978 11376 33390
rect 11336 32972 11388 32978
rect 11336 32914 11388 32920
rect 11440 32774 11468 33510
rect 11796 33516 11848 33522
rect 11796 33458 11848 33464
rect 11610 33416 11666 33425
rect 11900 33402 11928 34002
rect 11610 33351 11612 33360
rect 11664 33351 11666 33360
rect 11808 33374 11928 33402
rect 11612 33322 11664 33328
rect 11808 32978 11836 33374
rect 11796 32972 11848 32978
rect 11796 32914 11848 32920
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11428 32768 11480 32774
rect 11428 32710 11480 32716
rect 11244 32564 11296 32570
rect 11244 32506 11296 32512
rect 11256 32366 11284 32506
rect 11348 32366 11376 32710
rect 11436 32668 11744 32677
rect 11436 32666 11442 32668
rect 11498 32666 11522 32668
rect 11578 32666 11602 32668
rect 11658 32666 11682 32668
rect 11738 32666 11744 32668
rect 11498 32614 11500 32666
rect 11680 32614 11682 32666
rect 11436 32612 11442 32614
rect 11498 32612 11522 32614
rect 11578 32612 11602 32614
rect 11658 32612 11682 32614
rect 11738 32612 11744 32614
rect 11436 32603 11744 32612
rect 11808 32434 11836 32914
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11244 32360 11296 32366
rect 11244 32302 11296 32308
rect 11336 32360 11388 32366
rect 11336 32302 11388 32308
rect 11244 32224 11296 32230
rect 11244 32166 11296 32172
rect 11888 32224 11940 32230
rect 11888 32166 11940 32172
rect 11152 31476 11204 31482
rect 11152 31418 11204 31424
rect 11256 31346 11284 32166
rect 11336 31952 11388 31958
rect 11336 31894 11388 31900
rect 11244 31340 11296 31346
rect 11244 31282 11296 31288
rect 11348 31278 11376 31894
rect 11436 31580 11744 31589
rect 11436 31578 11442 31580
rect 11498 31578 11522 31580
rect 11578 31578 11602 31580
rect 11658 31578 11682 31580
rect 11738 31578 11744 31580
rect 11498 31526 11500 31578
rect 11680 31526 11682 31578
rect 11436 31524 11442 31526
rect 11498 31524 11522 31526
rect 11578 31524 11602 31526
rect 11658 31524 11682 31526
rect 11738 31524 11744 31526
rect 11436 31515 11744 31524
rect 11900 31414 11928 32166
rect 11888 31408 11940 31414
rect 11888 31350 11940 31356
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 11888 31272 11940 31278
rect 11888 31214 11940 31220
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 10324 30932 10376 30938
rect 10324 30874 10376 30880
rect 10048 30796 10100 30802
rect 10048 30738 10100 30744
rect 10336 30734 10364 30874
rect 10324 30728 10376 30734
rect 10324 30670 10376 30676
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 11348 30190 11376 31078
rect 11612 30932 11664 30938
rect 11612 30874 11664 30880
rect 11624 30734 11652 30874
rect 11900 30802 11928 31214
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 11612 30728 11664 30734
rect 11612 30670 11664 30676
rect 11900 30598 11928 30738
rect 11888 30592 11940 30598
rect 11888 30534 11940 30540
rect 11436 30492 11744 30501
rect 11436 30490 11442 30492
rect 11498 30490 11522 30492
rect 11578 30490 11602 30492
rect 11658 30490 11682 30492
rect 11738 30490 11744 30492
rect 11498 30438 11500 30490
rect 11680 30438 11682 30490
rect 11436 30436 11442 30438
rect 11498 30436 11522 30438
rect 11578 30436 11602 30438
rect 11658 30436 11682 30438
rect 11738 30436 11744 30438
rect 11436 30427 11744 30436
rect 11992 30274 12020 35006
rect 12084 34746 12112 35090
rect 12176 34950 12204 35090
rect 12164 34944 12216 34950
rect 12164 34886 12216 34892
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 12452 34678 12480 35550
rect 12636 35222 12664 35770
rect 12808 35692 12860 35698
rect 12808 35634 12860 35640
rect 12624 35216 12676 35222
rect 12624 35158 12676 35164
rect 12716 35080 12768 35086
rect 12714 35048 12716 35057
rect 12768 35048 12770 35057
rect 12714 34983 12770 34992
rect 12440 34672 12492 34678
rect 12440 34614 12492 34620
rect 12820 34542 12848 35634
rect 12912 35494 12940 36178
rect 12900 35488 12952 35494
rect 12900 35430 12952 35436
rect 12808 34536 12860 34542
rect 12808 34478 12860 34484
rect 12900 34536 12952 34542
rect 12900 34478 12952 34484
rect 12096 34300 12404 34309
rect 12096 34298 12102 34300
rect 12158 34298 12182 34300
rect 12238 34298 12262 34300
rect 12318 34298 12342 34300
rect 12398 34298 12404 34300
rect 12158 34246 12160 34298
rect 12340 34246 12342 34298
rect 12096 34244 12102 34246
rect 12158 34244 12182 34246
rect 12238 34244 12262 34246
rect 12318 34244 12342 34246
rect 12398 34244 12404 34246
rect 12096 34235 12404 34244
rect 12440 34128 12492 34134
rect 12440 34070 12492 34076
rect 12072 33924 12124 33930
rect 12072 33866 12124 33872
rect 12084 33454 12112 33866
rect 12348 33584 12400 33590
rect 12348 33526 12400 33532
rect 12360 33454 12388 33526
rect 12072 33448 12124 33454
rect 12072 33390 12124 33396
rect 12348 33448 12400 33454
rect 12348 33390 12400 33396
rect 12452 33318 12480 34070
rect 12716 33924 12768 33930
rect 12716 33866 12768 33872
rect 12532 33448 12584 33454
rect 12530 33416 12532 33425
rect 12624 33448 12676 33454
rect 12584 33416 12586 33425
rect 12624 33390 12676 33396
rect 12530 33351 12586 33360
rect 12440 33312 12492 33318
rect 12440 33254 12492 33260
rect 12096 33212 12404 33221
rect 12096 33210 12102 33212
rect 12158 33210 12182 33212
rect 12238 33210 12262 33212
rect 12318 33210 12342 33212
rect 12398 33210 12404 33212
rect 12158 33158 12160 33210
rect 12340 33158 12342 33210
rect 12096 33156 12102 33158
rect 12158 33156 12182 33158
rect 12238 33156 12262 33158
rect 12318 33156 12342 33158
rect 12398 33156 12404 33158
rect 12096 33147 12404 33156
rect 12636 33046 12664 33390
rect 12624 33040 12676 33046
rect 12624 32982 12676 32988
rect 12728 32910 12756 33866
rect 12820 33862 12848 34478
rect 12912 34202 12940 34478
rect 12900 34196 12952 34202
rect 12900 34138 12952 34144
rect 13004 34066 13032 36518
rect 13188 36378 13216 39902
rect 13280 38350 13308 40054
rect 14108 39982 14136 40394
rect 13544 39976 13596 39982
rect 13544 39918 13596 39924
rect 14096 39976 14148 39982
rect 14096 39918 14148 39924
rect 13452 39908 13504 39914
rect 13452 39850 13504 39856
rect 13464 39642 13492 39850
rect 13556 39642 13584 39918
rect 13636 39840 13688 39846
rect 13688 39800 13768 39828
rect 13636 39782 13688 39788
rect 13452 39636 13504 39642
rect 13452 39578 13504 39584
rect 13544 39636 13596 39642
rect 13544 39578 13596 39584
rect 13740 39370 13768 39800
rect 13636 39364 13688 39370
rect 13636 39306 13688 39312
rect 13728 39364 13780 39370
rect 13728 39306 13780 39312
rect 13360 39296 13412 39302
rect 13360 39238 13412 39244
rect 13268 38344 13320 38350
rect 13268 38286 13320 38292
rect 13280 36922 13308 38286
rect 13268 36916 13320 36922
rect 13268 36858 13320 36864
rect 13176 36372 13228 36378
rect 13176 36314 13228 36320
rect 13084 35624 13136 35630
rect 13188 35612 13216 36314
rect 13136 35584 13216 35612
rect 13084 35566 13136 35572
rect 13188 34474 13216 35584
rect 13268 35556 13320 35562
rect 13268 35498 13320 35504
rect 13280 34542 13308 35498
rect 13372 35154 13400 39238
rect 13648 38962 13676 39306
rect 13636 38956 13688 38962
rect 13636 38898 13688 38904
rect 13452 38480 13504 38486
rect 13452 38422 13504 38428
rect 13464 35698 13492 38422
rect 13648 36106 13676 38898
rect 13740 37126 13768 39306
rect 14096 38752 14148 38758
rect 14096 38694 14148 38700
rect 14108 38418 14136 38694
rect 13820 38412 13872 38418
rect 13820 38354 13872 38360
rect 14096 38412 14148 38418
rect 14096 38354 14148 38360
rect 13728 37120 13780 37126
rect 13728 37062 13780 37068
rect 13832 36854 13860 38354
rect 14188 38208 14240 38214
rect 14188 38150 14240 38156
rect 14200 37738 14228 38150
rect 13912 37732 13964 37738
rect 13912 37674 13964 37680
rect 14188 37732 14240 37738
rect 14188 37674 14240 37680
rect 13820 36848 13872 36854
rect 13820 36790 13872 36796
rect 13832 36242 13860 36790
rect 13820 36236 13872 36242
rect 13820 36178 13872 36184
rect 13636 36100 13688 36106
rect 13636 36042 13688 36048
rect 13924 36038 13952 37674
rect 14188 36644 14240 36650
rect 14188 36586 14240 36592
rect 14004 36100 14056 36106
rect 14004 36042 14056 36048
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13452 35692 13504 35698
rect 13452 35634 13504 35640
rect 13544 35556 13596 35562
rect 13544 35498 13596 35504
rect 13728 35556 13780 35562
rect 13728 35498 13780 35504
rect 13360 35148 13412 35154
rect 13360 35090 13412 35096
rect 13452 34944 13504 34950
rect 13452 34886 13504 34892
rect 13464 34678 13492 34886
rect 13452 34672 13504 34678
rect 13452 34614 13504 34620
rect 13268 34536 13320 34542
rect 13268 34478 13320 34484
rect 13176 34468 13228 34474
rect 13176 34410 13228 34416
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 13280 33930 13308 34478
rect 13268 33924 13320 33930
rect 13268 33866 13320 33872
rect 12808 33856 12860 33862
rect 12808 33798 12860 33804
rect 12820 33590 12848 33798
rect 12808 33584 12860 33590
rect 12808 33526 12860 33532
rect 13464 32978 13492 34614
rect 13556 34134 13584 35498
rect 13740 35154 13768 35498
rect 13636 35148 13688 35154
rect 13636 35090 13688 35096
rect 13728 35148 13780 35154
rect 13728 35090 13780 35096
rect 13648 35018 13676 35090
rect 13740 35057 13768 35090
rect 13726 35048 13782 35057
rect 13636 35012 13688 35018
rect 13726 34983 13782 34992
rect 13636 34954 13688 34960
rect 13544 34128 13596 34134
rect 13544 34070 13596 34076
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13452 32972 13504 32978
rect 13452 32914 13504 32920
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12348 32768 12400 32774
rect 12348 32710 12400 32716
rect 12532 32768 12584 32774
rect 12532 32710 12584 32716
rect 12360 32366 12388 32710
rect 12544 32366 12572 32710
rect 12348 32360 12400 32366
rect 12348 32302 12400 32308
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12440 32292 12492 32298
rect 12440 32234 12492 32240
rect 12096 32124 12404 32133
rect 12096 32122 12102 32124
rect 12158 32122 12182 32124
rect 12238 32122 12262 32124
rect 12318 32122 12342 32124
rect 12398 32122 12404 32124
rect 12158 32070 12160 32122
rect 12340 32070 12342 32122
rect 12096 32068 12102 32070
rect 12158 32068 12182 32070
rect 12238 32068 12262 32070
rect 12318 32068 12342 32070
rect 12398 32068 12404 32070
rect 12096 32059 12404 32068
rect 12452 32008 12480 32234
rect 12360 31980 12480 32008
rect 12360 31686 12388 31980
rect 12728 31890 12756 32846
rect 13464 32570 13492 32914
rect 13452 32564 13504 32570
rect 13452 32506 13504 32512
rect 12808 32360 12860 32366
rect 12808 32302 12860 32308
rect 12716 31884 12768 31890
rect 12716 31826 12768 31832
rect 12820 31822 12848 32302
rect 13556 31890 13584 33934
rect 13648 33658 13676 34954
rect 13740 34474 13768 34983
rect 13912 34944 13964 34950
rect 13912 34886 13964 34892
rect 13924 34542 13952 34886
rect 13912 34536 13964 34542
rect 13912 34478 13964 34484
rect 13728 34468 13780 34474
rect 13728 34410 13780 34416
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13636 33312 13688 33318
rect 13636 33254 13688 33260
rect 13648 32978 13676 33254
rect 13636 32972 13688 32978
rect 13636 32914 13688 32920
rect 13740 31890 13768 34410
rect 13912 34400 13964 34406
rect 13912 34342 13964 34348
rect 13924 33998 13952 34342
rect 13912 33992 13964 33998
rect 13912 33934 13964 33940
rect 14016 33454 14044 36042
rect 14200 34406 14228 36586
rect 14292 36530 14320 41754
rect 14372 40928 14424 40934
rect 14372 40870 14424 40876
rect 14384 40594 14412 40870
rect 14372 40588 14424 40594
rect 14372 40530 14424 40536
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 14384 37466 14412 38150
rect 14372 37460 14424 37466
rect 14372 37402 14424 37408
rect 14292 36502 14412 36530
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14292 36009 14320 36110
rect 14278 36000 14334 36009
rect 14278 35935 14334 35944
rect 14280 35148 14332 35154
rect 14280 35090 14332 35096
rect 14188 34400 14240 34406
rect 14188 34342 14240 34348
rect 14292 34202 14320 35090
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 14188 33448 14240 33454
rect 14188 33390 14240 33396
rect 14200 33046 14228 33390
rect 14188 33040 14240 33046
rect 14188 32982 14240 32988
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 13832 32502 13860 32914
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 13820 32224 13872 32230
rect 13820 32166 13872 32172
rect 13544 31884 13596 31890
rect 13544 31826 13596 31832
rect 13728 31884 13780 31890
rect 13728 31826 13780 31832
rect 12808 31816 12860 31822
rect 12808 31758 12860 31764
rect 12716 31748 12768 31754
rect 12716 31690 12768 31696
rect 12348 31680 12400 31686
rect 12348 31622 12400 31628
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 12360 31278 12388 31350
rect 12348 31272 12400 31278
rect 12348 31214 12400 31220
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12096 31036 12404 31045
rect 12096 31034 12102 31036
rect 12158 31034 12182 31036
rect 12238 31034 12262 31036
rect 12318 31034 12342 31036
rect 12398 31034 12404 31036
rect 12158 30982 12160 31034
rect 12340 30982 12342 31034
rect 12096 30980 12102 30982
rect 12158 30980 12182 30982
rect 12238 30980 12262 30982
rect 12318 30980 12342 30982
rect 12398 30980 12404 30982
rect 12096 30971 12404 30980
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12084 30394 12112 30670
rect 12072 30388 12124 30394
rect 12072 30330 12124 30336
rect 11900 30246 12020 30274
rect 11336 30184 11388 30190
rect 11336 30126 11388 30132
rect 9404 30116 9456 30122
rect 9404 30058 9456 30064
rect 9588 30116 9640 30122
rect 9588 30058 9640 30064
rect 4322 29948 4630 29957
rect 4322 29946 4328 29948
rect 4384 29946 4408 29948
rect 4464 29946 4488 29948
rect 4544 29946 4568 29948
rect 4624 29946 4630 29948
rect 4384 29894 4386 29946
rect 4566 29894 4568 29946
rect 4322 29892 4328 29894
rect 4384 29892 4408 29894
rect 4464 29892 4488 29894
rect 4544 29892 4568 29894
rect 4624 29892 4630 29894
rect 4322 29883 4630 29892
rect 3662 29404 3970 29413
rect 3662 29402 3668 29404
rect 3724 29402 3748 29404
rect 3804 29402 3828 29404
rect 3884 29402 3908 29404
rect 3964 29402 3970 29404
rect 3724 29350 3726 29402
rect 3906 29350 3908 29402
rect 3662 29348 3668 29350
rect 3724 29348 3748 29350
rect 3804 29348 3828 29350
rect 3884 29348 3908 29350
rect 3964 29348 3970 29350
rect 3662 29339 3970 29348
rect 9416 29102 9444 30058
rect 11900 29782 11928 30246
rect 12176 30138 12204 30670
rect 11992 30110 12204 30138
rect 11888 29776 11940 29782
rect 11888 29718 11940 29724
rect 11436 29404 11744 29413
rect 11436 29402 11442 29404
rect 11498 29402 11522 29404
rect 11578 29402 11602 29404
rect 11658 29402 11682 29404
rect 11738 29402 11744 29404
rect 11498 29350 11500 29402
rect 11680 29350 11682 29402
rect 11436 29348 11442 29350
rect 11498 29348 11522 29350
rect 11578 29348 11602 29350
rect 11658 29348 11682 29350
rect 11738 29348 11744 29350
rect 11436 29339 11744 29348
rect 11900 29306 11928 29718
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11336 29232 11388 29238
rect 11336 29174 11388 29180
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 4322 28860 4630 28869
rect 4322 28858 4328 28860
rect 4384 28858 4408 28860
rect 4464 28858 4488 28860
rect 4544 28858 4568 28860
rect 4624 28858 4630 28860
rect 4384 28806 4386 28858
rect 4566 28806 4568 28858
rect 4322 28804 4328 28806
rect 4384 28804 4408 28806
rect 4464 28804 4488 28806
rect 4544 28804 4568 28806
rect 4624 28804 4630 28806
rect 4322 28795 4630 28804
rect 11072 28626 11100 28902
rect 11060 28620 11112 28626
rect 11060 28562 11112 28568
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 3662 28316 3970 28325
rect 3662 28314 3668 28316
rect 3724 28314 3748 28316
rect 3804 28314 3828 28316
rect 3884 28314 3908 28316
rect 3964 28314 3970 28316
rect 3724 28262 3726 28314
rect 3906 28262 3908 28314
rect 3662 28260 3668 28262
rect 3724 28260 3748 28262
rect 3804 28260 3828 28262
rect 3884 28260 3908 28262
rect 3964 28260 3970 28262
rect 3662 28251 3970 28260
rect 11256 28218 11284 28562
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 11348 28014 11376 29174
rect 11532 29102 11560 29242
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11716 29102 11744 29174
rect 11520 29096 11572 29102
rect 11520 29038 11572 29044
rect 11704 29096 11756 29102
rect 11704 29038 11756 29044
rect 11716 28506 11744 29038
rect 11992 29034 12020 30110
rect 12096 29948 12404 29957
rect 12096 29946 12102 29948
rect 12158 29946 12182 29948
rect 12238 29946 12262 29948
rect 12318 29946 12342 29948
rect 12398 29946 12404 29948
rect 12158 29894 12160 29946
rect 12340 29894 12342 29946
rect 12096 29892 12102 29894
rect 12158 29892 12182 29894
rect 12238 29892 12262 29894
rect 12318 29892 12342 29894
rect 12398 29892 12404 29894
rect 12096 29883 12404 29892
rect 12452 29102 12480 31214
rect 12728 30938 12756 31690
rect 12820 31482 12848 31758
rect 12808 31476 12860 31482
rect 12808 31418 12860 31424
rect 13452 31340 13504 31346
rect 13452 31282 13504 31288
rect 12808 31204 12860 31210
rect 12808 31146 12860 31152
rect 12820 30938 12848 31146
rect 13084 31136 13136 31142
rect 13084 31078 13136 31084
rect 12716 30932 12768 30938
rect 12716 30874 12768 30880
rect 12808 30932 12860 30938
rect 12808 30874 12860 30880
rect 12728 30666 12756 30874
rect 13096 30802 13124 31078
rect 13464 30938 13492 31282
rect 13832 31278 13860 32166
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 14200 31210 14228 32982
rect 14188 31204 14240 31210
rect 14240 31164 14320 31192
rect 14188 31146 14240 31152
rect 13452 30932 13504 30938
rect 13452 30874 13504 30880
rect 13084 30796 13136 30802
rect 13084 30738 13136 30744
rect 13268 30796 13320 30802
rect 13268 30738 13320 30744
rect 12716 30660 12768 30666
rect 12716 30602 12768 30608
rect 12532 30592 12584 30598
rect 12532 30534 12584 30540
rect 12544 30326 12572 30534
rect 12532 30320 12584 30326
rect 12532 30262 12584 30268
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 13096 29102 13124 29242
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 13084 29096 13136 29102
rect 13084 29038 13136 29044
rect 13176 29096 13228 29102
rect 13176 29038 13228 29044
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 11992 28762 12020 28970
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 12096 28860 12404 28869
rect 12096 28858 12102 28860
rect 12158 28858 12182 28860
rect 12238 28858 12262 28860
rect 12318 28858 12342 28860
rect 12398 28858 12404 28860
rect 12158 28806 12160 28858
rect 12340 28806 12342 28858
rect 12096 28804 12102 28806
rect 12158 28804 12182 28806
rect 12238 28804 12262 28806
rect 12318 28804 12342 28806
rect 12398 28804 12404 28806
rect 12096 28795 12404 28804
rect 11980 28756 12032 28762
rect 11980 28698 12032 28704
rect 11716 28478 11836 28506
rect 11436 28316 11744 28325
rect 11436 28314 11442 28316
rect 11498 28314 11522 28316
rect 11578 28314 11602 28316
rect 11658 28314 11682 28316
rect 11738 28314 11744 28316
rect 11498 28262 11500 28314
rect 11680 28262 11682 28314
rect 11436 28260 11442 28262
rect 11498 28260 11522 28262
rect 11578 28260 11602 28262
rect 11658 28260 11682 28262
rect 11738 28260 11744 28262
rect 11436 28251 11744 28260
rect 11808 28014 11836 28478
rect 11336 28008 11388 28014
rect 11336 27950 11388 27956
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 4322 27772 4630 27781
rect 4322 27770 4328 27772
rect 4384 27770 4408 27772
rect 4464 27770 4488 27772
rect 4544 27770 4568 27772
rect 4624 27770 4630 27772
rect 4384 27718 4386 27770
rect 4566 27718 4568 27770
rect 4322 27716 4328 27718
rect 4384 27716 4408 27718
rect 4464 27716 4488 27718
rect 4544 27716 4568 27718
rect 4624 27716 4630 27718
rect 4322 27707 4630 27716
rect 11716 27520 11744 27950
rect 11992 27946 12020 28698
rect 12452 28626 12480 28902
rect 12636 28626 12664 28902
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 13188 28558 13216 29038
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 11980 27940 12032 27946
rect 11980 27882 12032 27888
rect 11796 27532 11848 27538
rect 11716 27492 11796 27520
rect 11796 27474 11848 27480
rect 11808 27402 11836 27474
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11992 27334 12020 27882
rect 12096 27772 12404 27781
rect 12096 27770 12102 27772
rect 12158 27770 12182 27772
rect 12238 27770 12262 27772
rect 12318 27770 12342 27772
rect 12398 27770 12404 27772
rect 12158 27718 12160 27770
rect 12340 27718 12342 27770
rect 12096 27716 12102 27718
rect 12158 27716 12182 27718
rect 12238 27716 12262 27718
rect 12318 27716 12342 27718
rect 12398 27716 12404 27718
rect 12096 27707 12404 27716
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 3662 27228 3970 27237
rect 3662 27226 3668 27228
rect 3724 27226 3748 27228
rect 3804 27226 3828 27228
rect 3884 27226 3908 27228
rect 3964 27226 3970 27228
rect 3724 27174 3726 27226
rect 3906 27174 3908 27226
rect 3662 27172 3668 27174
rect 3724 27172 3748 27174
rect 3804 27172 3828 27174
rect 3884 27172 3908 27174
rect 3964 27172 3970 27174
rect 3662 27163 3970 27172
rect 11348 27010 11376 27270
rect 11436 27228 11744 27237
rect 11436 27226 11442 27228
rect 11498 27226 11522 27228
rect 11578 27226 11602 27228
rect 11658 27226 11682 27228
rect 11738 27226 11744 27228
rect 11498 27174 11500 27226
rect 11680 27174 11682 27226
rect 11436 27172 11442 27174
rect 11498 27172 11522 27174
rect 11578 27172 11602 27174
rect 11658 27172 11682 27174
rect 11738 27172 11744 27174
rect 11436 27163 11744 27172
rect 12544 27130 12572 27474
rect 13188 27470 13216 28494
rect 13280 28014 13308 30738
rect 14188 30660 14240 30666
rect 14188 30602 14240 30608
rect 14096 30048 14148 30054
rect 14096 29990 14148 29996
rect 14108 29714 14136 29990
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 14200 29102 14228 30602
rect 14292 30190 14320 31164
rect 14280 30184 14332 30190
rect 14280 30126 14332 30132
rect 14384 29306 14412 36502
rect 14476 31958 14504 44254
rect 15752 44192 15804 44198
rect 15752 44134 15804 44140
rect 15292 43784 15344 43790
rect 15292 43726 15344 43732
rect 15304 43450 15332 43726
rect 15292 43444 15344 43450
rect 15292 43386 15344 43392
rect 15016 43240 15068 43246
rect 15660 43240 15712 43246
rect 15016 43182 15068 43188
rect 15106 43208 15162 43217
rect 15028 42906 15056 43182
rect 15660 43182 15712 43188
rect 15106 43143 15162 43152
rect 15016 42900 15068 42906
rect 15016 42842 15068 42848
rect 14648 42764 14700 42770
rect 14648 42706 14700 42712
rect 14660 42158 14688 42706
rect 15016 42696 15068 42702
rect 15016 42638 15068 42644
rect 15028 42362 15056 42638
rect 15016 42356 15068 42362
rect 15016 42298 15068 42304
rect 14648 42152 14700 42158
rect 14648 42094 14700 42100
rect 14832 41676 14884 41682
rect 14832 41618 14884 41624
rect 14556 37324 14608 37330
rect 14556 37266 14608 37272
rect 14568 36922 14596 37266
rect 14556 36916 14608 36922
rect 14556 36858 14608 36864
rect 14568 36786 14596 36858
rect 14556 36780 14608 36786
rect 14556 36722 14608 36728
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14568 36378 14596 36518
rect 14556 36372 14608 36378
rect 14556 36314 14608 36320
rect 14740 36032 14792 36038
rect 14740 35974 14792 35980
rect 14648 35828 14700 35834
rect 14648 35770 14700 35776
rect 14660 35154 14688 35770
rect 14752 35154 14780 35974
rect 14556 35148 14608 35154
rect 14556 35090 14608 35096
rect 14648 35148 14700 35154
rect 14648 35090 14700 35096
rect 14740 35148 14792 35154
rect 14740 35090 14792 35096
rect 14568 34746 14596 35090
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 14660 32978 14688 35090
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 14752 34066 14780 34682
rect 14740 34060 14792 34066
rect 14740 34002 14792 34008
rect 14648 32972 14700 32978
rect 14648 32914 14700 32920
rect 14464 31952 14516 31958
rect 14464 31894 14516 31900
rect 14556 31816 14608 31822
rect 14556 31758 14608 31764
rect 14464 31680 14516 31686
rect 14464 31622 14516 31628
rect 14476 30870 14504 31622
rect 14464 30864 14516 30870
rect 14464 30806 14516 30812
rect 14568 30802 14596 31758
rect 14556 30796 14608 30802
rect 14556 30738 14608 30744
rect 14648 29776 14700 29782
rect 14648 29718 14700 29724
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14384 29102 14412 29242
rect 14660 29186 14688 29718
rect 14740 29708 14792 29714
rect 14740 29650 14792 29656
rect 14752 29306 14780 29650
rect 14740 29300 14792 29306
rect 14740 29242 14792 29248
rect 14660 29158 14780 29186
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 14372 29096 14424 29102
rect 14372 29038 14424 29044
rect 14200 28694 14228 29038
rect 14278 28792 14334 28801
rect 14278 28727 14280 28736
rect 14332 28727 14334 28736
rect 14280 28698 14332 28704
rect 14188 28688 14240 28694
rect 14188 28630 14240 28636
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 13280 27538 13308 27950
rect 13820 27940 13872 27946
rect 13820 27882 13872 27888
rect 13268 27532 13320 27538
rect 13268 27474 13320 27480
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 11348 26982 11468 27010
rect 11440 26926 11468 26982
rect 13740 26926 13768 27474
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 4322 26684 4630 26693
rect 4322 26682 4328 26684
rect 4384 26682 4408 26684
rect 4464 26682 4488 26684
rect 4544 26682 4568 26684
rect 4624 26682 4630 26684
rect 4384 26630 4386 26682
rect 4566 26630 4568 26682
rect 4322 26628 4328 26630
rect 4384 26628 4408 26630
rect 4464 26628 4488 26630
rect 4544 26628 4568 26630
rect 4624 26628 4630 26630
rect 4322 26619 4630 26628
rect 3662 26140 3970 26149
rect 3662 26138 3668 26140
rect 3724 26138 3748 26140
rect 3804 26138 3828 26140
rect 3884 26138 3908 26140
rect 3964 26138 3970 26140
rect 3724 26086 3726 26138
rect 3906 26086 3908 26138
rect 3662 26084 3668 26086
rect 3724 26084 3748 26086
rect 3804 26084 3828 26086
rect 3884 26084 3908 26086
rect 3964 26084 3970 26086
rect 3662 26075 3970 26084
rect 11256 25820 11284 26862
rect 12096 26684 12404 26693
rect 12096 26682 12102 26684
rect 12158 26682 12182 26684
rect 12238 26682 12262 26684
rect 12318 26682 12342 26684
rect 12398 26682 12404 26684
rect 12158 26630 12160 26682
rect 12340 26630 12342 26682
rect 12096 26628 12102 26630
rect 12158 26628 12182 26630
rect 12238 26628 12262 26630
rect 12318 26628 12342 26630
rect 12398 26628 12404 26630
rect 12096 26619 12404 26628
rect 13832 26586 13860 27882
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14016 27130 14044 27474
rect 14004 27124 14056 27130
rect 14004 27066 14056 27072
rect 14200 26790 14228 28630
rect 14752 28558 14780 29158
rect 14844 28762 14872 41618
rect 15016 41540 15068 41546
rect 15016 41482 15068 41488
rect 15028 40050 15056 41482
rect 15120 41070 15148 43143
rect 15568 43104 15620 43110
rect 15568 43046 15620 43052
rect 15474 42936 15530 42945
rect 15474 42871 15476 42880
rect 15528 42871 15530 42880
rect 15476 42842 15528 42848
rect 15488 42294 15516 42842
rect 15476 42288 15528 42294
rect 15476 42230 15528 42236
rect 15476 42152 15528 42158
rect 15476 42094 15528 42100
rect 15200 42016 15252 42022
rect 15200 41958 15252 41964
rect 15212 41206 15240 41958
rect 15384 41472 15436 41478
rect 15384 41414 15436 41420
rect 15396 41290 15424 41414
rect 15304 41262 15424 41290
rect 15200 41200 15252 41206
rect 15200 41142 15252 41148
rect 15108 41064 15160 41070
rect 15108 41006 15160 41012
rect 15200 41064 15252 41070
rect 15304 41052 15332 41262
rect 15252 41024 15332 41052
rect 15384 41064 15436 41070
rect 15200 41006 15252 41012
rect 15384 41006 15436 41012
rect 15120 40730 15148 41006
rect 15200 40928 15252 40934
rect 15200 40870 15252 40876
rect 15292 40928 15344 40934
rect 15292 40870 15344 40876
rect 15108 40724 15160 40730
rect 15108 40666 15160 40672
rect 15016 40044 15068 40050
rect 15016 39986 15068 39992
rect 14924 39840 14976 39846
rect 14924 39782 14976 39788
rect 14936 39438 14964 39782
rect 14924 39432 14976 39438
rect 14924 39374 14976 39380
rect 15108 38548 15160 38554
rect 15108 38490 15160 38496
rect 14924 38412 14976 38418
rect 14924 38354 14976 38360
rect 14936 38010 14964 38354
rect 14924 38004 14976 38010
rect 14924 37946 14976 37952
rect 15120 37194 15148 38490
rect 15212 38486 15240 40870
rect 15200 38480 15252 38486
rect 15200 38422 15252 38428
rect 15304 37346 15332 40870
rect 15396 40186 15424 41006
rect 15384 40180 15436 40186
rect 15384 40122 15436 40128
rect 15384 40044 15436 40050
rect 15384 39986 15436 39992
rect 15396 39302 15424 39986
rect 15488 39642 15516 42094
rect 15580 41274 15608 43046
rect 15672 42226 15700 43182
rect 15660 42220 15712 42226
rect 15660 42162 15712 42168
rect 15672 41478 15700 42162
rect 15764 42158 15792 44134
rect 15856 43722 15884 44270
rect 16120 43852 16172 43858
rect 16120 43794 16172 43800
rect 15844 43716 15896 43722
rect 15844 43658 15896 43664
rect 15856 43246 15884 43658
rect 15844 43240 15896 43246
rect 15844 43182 15896 43188
rect 16028 43240 16080 43246
rect 16028 43182 16080 43188
rect 15752 42152 15804 42158
rect 15752 42094 15804 42100
rect 15764 42022 15792 42094
rect 15752 42016 15804 42022
rect 15752 41958 15804 41964
rect 15856 41546 15884 43182
rect 16040 42634 16068 43182
rect 16028 42628 16080 42634
rect 16028 42570 16080 42576
rect 16132 41546 16160 43794
rect 16500 43314 16528 44270
rect 16764 44192 16816 44198
rect 16764 44134 16816 44140
rect 19248 44192 19300 44198
rect 19248 44134 19300 44140
rect 21824 44192 21876 44198
rect 21824 44134 21876 44140
rect 22008 44192 22060 44198
rect 22008 44134 22060 44140
rect 24584 44192 24636 44198
rect 24584 44134 24636 44140
rect 25136 44192 25188 44198
rect 25136 44134 25188 44140
rect 16578 44024 16634 44033
rect 16578 43959 16634 43968
rect 16592 43926 16620 43959
rect 16580 43920 16632 43926
rect 16580 43862 16632 43868
rect 16488 43308 16540 43314
rect 16488 43250 16540 43256
rect 16304 43240 16356 43246
rect 16304 43182 16356 43188
rect 16316 42906 16344 43182
rect 16396 43104 16448 43110
rect 16396 43046 16448 43052
rect 16304 42900 16356 42906
rect 16304 42842 16356 42848
rect 16212 42764 16264 42770
rect 16212 42706 16264 42712
rect 16224 41750 16252 42706
rect 16316 42702 16344 42842
rect 16304 42696 16356 42702
rect 16304 42638 16356 42644
rect 16408 42294 16436 43046
rect 16396 42288 16448 42294
rect 16396 42230 16448 42236
rect 16212 41744 16264 41750
rect 16212 41686 16264 41692
rect 15844 41540 15896 41546
rect 15844 41482 15896 41488
rect 16120 41540 16172 41546
rect 16120 41482 16172 41488
rect 15660 41472 15712 41478
rect 15660 41414 15712 41420
rect 15568 41268 15620 41274
rect 15568 41210 15620 41216
rect 15568 41064 15620 41070
rect 15568 41006 15620 41012
rect 15580 39982 15608 41006
rect 15568 39976 15620 39982
rect 15568 39918 15620 39924
rect 15476 39636 15528 39642
rect 15476 39578 15528 39584
rect 15580 39506 15608 39918
rect 15568 39500 15620 39506
rect 15568 39442 15620 39448
rect 15384 39296 15436 39302
rect 15384 39238 15436 39244
rect 15396 37806 15424 39238
rect 15568 39024 15620 39030
rect 15568 38966 15620 38972
rect 15476 38752 15528 38758
rect 15476 38694 15528 38700
rect 15488 37806 15516 38694
rect 15580 37806 15608 38966
rect 15672 38894 15700 41414
rect 15936 41064 15988 41070
rect 15936 41006 15988 41012
rect 16120 41064 16172 41070
rect 16120 41006 16172 41012
rect 15844 40384 15896 40390
rect 15844 40326 15896 40332
rect 15856 39982 15884 40326
rect 15948 39982 15976 41006
rect 16132 40186 16160 41006
rect 16224 40594 16252 41686
rect 16500 41274 16528 43250
rect 16592 43246 16620 43862
rect 16776 43858 16804 44134
rect 17406 44024 17462 44033
rect 17406 43959 17462 43968
rect 18142 44024 18198 44033
rect 18142 43959 18144 43968
rect 16764 43852 16816 43858
rect 16764 43794 16816 43800
rect 17040 43784 17092 43790
rect 17040 43726 17092 43732
rect 16580 43240 16632 43246
rect 16632 43200 16712 43228
rect 16580 43182 16632 43188
rect 16580 43104 16632 43110
rect 16580 43046 16632 43052
rect 16488 41268 16540 41274
rect 16488 41210 16540 41216
rect 16302 41168 16358 41177
rect 16302 41103 16358 41112
rect 16316 41070 16344 41103
rect 16304 41064 16356 41070
rect 16304 41006 16356 41012
rect 16212 40588 16264 40594
rect 16212 40530 16264 40536
rect 16120 40180 16172 40186
rect 16120 40122 16172 40128
rect 15844 39976 15896 39982
rect 15844 39918 15896 39924
rect 15936 39976 15988 39982
rect 15936 39918 15988 39924
rect 15948 39522 15976 39918
rect 15856 39494 15976 39522
rect 15856 39438 15884 39494
rect 15844 39432 15896 39438
rect 15844 39374 15896 39380
rect 15660 38888 15712 38894
rect 15660 38830 15712 38836
rect 15672 38554 15700 38830
rect 15660 38548 15712 38554
rect 15660 38490 15712 38496
rect 15660 38208 15712 38214
rect 15660 38150 15712 38156
rect 15752 38208 15804 38214
rect 15752 38150 15804 38156
rect 15384 37800 15436 37806
rect 15384 37742 15436 37748
rect 15476 37800 15528 37806
rect 15476 37742 15528 37748
rect 15568 37800 15620 37806
rect 15568 37742 15620 37748
rect 15672 37466 15700 38150
rect 15660 37460 15712 37466
rect 15660 37402 15712 37408
rect 15200 37324 15252 37330
rect 15304 37318 15424 37346
rect 15200 37266 15252 37272
rect 15108 37188 15160 37194
rect 15108 37130 15160 37136
rect 15120 36922 15148 37130
rect 15108 36916 15160 36922
rect 15108 36858 15160 36864
rect 15016 35692 15068 35698
rect 15016 35634 15068 35640
rect 15028 35222 15056 35634
rect 15016 35216 15068 35222
rect 15016 35158 15068 35164
rect 15108 35148 15160 35154
rect 15108 35090 15160 35096
rect 15120 34542 15148 35090
rect 15108 34536 15160 34542
rect 15108 34478 15160 34484
rect 15212 33046 15240 37266
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 15304 36174 15332 37198
rect 15292 36168 15344 36174
rect 15292 36110 15344 36116
rect 15292 35624 15344 35630
rect 15292 35566 15344 35572
rect 15304 34950 15332 35566
rect 15292 34944 15344 34950
rect 15292 34886 15344 34892
rect 15396 33862 15424 37318
rect 15660 37256 15712 37262
rect 15660 37198 15712 37204
rect 15568 37120 15620 37126
rect 15568 37062 15620 37068
rect 15580 36786 15608 37062
rect 15672 36854 15700 37198
rect 15660 36848 15712 36854
rect 15660 36790 15712 36796
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15580 36666 15608 36722
rect 15672 36718 15700 36790
rect 15488 36638 15608 36666
rect 15660 36712 15712 36718
rect 15660 36654 15712 36660
rect 15488 36242 15516 36638
rect 15568 36576 15620 36582
rect 15568 36518 15620 36524
rect 15476 36236 15528 36242
rect 15476 36178 15528 36184
rect 15476 35624 15528 35630
rect 15476 35566 15528 35572
rect 15488 35494 15516 35566
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15476 35284 15528 35290
rect 15476 35226 15528 35232
rect 15488 34950 15516 35226
rect 15476 34944 15528 34950
rect 15476 34886 15528 34892
rect 15488 34066 15516 34886
rect 15580 34066 15608 36518
rect 15764 35766 15792 38150
rect 15856 37806 15884 39374
rect 16316 38978 16344 41006
rect 16500 39846 16528 41210
rect 16592 39982 16620 43046
rect 16684 42906 16712 43200
rect 16764 43104 16816 43110
rect 16764 43046 16816 43052
rect 16672 42900 16724 42906
rect 16672 42842 16724 42848
rect 16776 42158 16804 43046
rect 16948 42764 17000 42770
rect 16948 42706 17000 42712
rect 16856 42220 16908 42226
rect 16856 42162 16908 42168
rect 16764 42152 16816 42158
rect 16764 42094 16816 42100
rect 16776 41818 16804 42094
rect 16764 41812 16816 41818
rect 16764 41754 16816 41760
rect 16672 40928 16724 40934
rect 16672 40870 16724 40876
rect 16684 40050 16712 40870
rect 16764 40724 16816 40730
rect 16764 40666 16816 40672
rect 16776 40594 16804 40666
rect 16868 40610 16896 42162
rect 16960 42158 16988 42706
rect 17052 42362 17080 43726
rect 17132 43376 17184 43382
rect 17132 43318 17184 43324
rect 17144 43246 17172 43318
rect 17420 43246 17448 43959
rect 18196 43959 18198 43968
rect 18144 43930 18196 43936
rect 19260 43858 19288 44134
rect 19870 44092 20178 44101
rect 19870 44090 19876 44092
rect 19932 44090 19956 44092
rect 20012 44090 20036 44092
rect 20092 44090 20116 44092
rect 20172 44090 20178 44092
rect 19932 44038 19934 44090
rect 20114 44038 20116 44090
rect 19870 44036 19876 44038
rect 19932 44036 19956 44038
rect 20012 44036 20036 44038
rect 20092 44036 20116 44038
rect 20172 44036 20178 44038
rect 19870 44027 20178 44036
rect 21836 43926 21864 44134
rect 21824 43920 21876 43926
rect 21824 43862 21876 43868
rect 19248 43852 19300 43858
rect 19248 43794 19300 43800
rect 19708 43784 19760 43790
rect 19708 43726 19760 43732
rect 19616 43648 19668 43654
rect 19616 43590 19668 43596
rect 19210 43548 19518 43557
rect 19210 43546 19216 43548
rect 19272 43546 19296 43548
rect 19352 43546 19376 43548
rect 19432 43546 19456 43548
rect 19512 43546 19518 43548
rect 19272 43494 19274 43546
rect 19454 43494 19456 43546
rect 19210 43492 19216 43494
rect 19272 43492 19296 43494
rect 19352 43492 19376 43494
rect 19432 43492 19456 43494
rect 19512 43492 19518 43494
rect 19210 43483 19518 43492
rect 19628 43353 19656 43590
rect 19614 43344 19670 43353
rect 17604 43302 17816 43330
rect 17132 43240 17184 43246
rect 17132 43182 17184 43188
rect 17408 43240 17460 43246
rect 17408 43182 17460 43188
rect 17500 43240 17552 43246
rect 17500 43182 17552 43188
rect 17144 42838 17172 43182
rect 17224 43104 17276 43110
rect 17512 43092 17540 43182
rect 17604 43110 17632 43302
rect 17788 43246 17816 43302
rect 19524 43308 19576 43314
rect 19614 43279 19670 43288
rect 19524 43250 19576 43256
rect 17776 43240 17828 43246
rect 18880 43240 18932 43246
rect 17776 43182 17828 43188
rect 18800 43200 18880 43228
rect 18144 43172 18196 43178
rect 18196 43132 18552 43160
rect 18144 43114 18196 43120
rect 17224 43046 17276 43052
rect 17420 43064 17540 43092
rect 17592 43104 17644 43110
rect 17132 42832 17184 42838
rect 17132 42774 17184 42780
rect 17040 42356 17092 42362
rect 17040 42298 17092 42304
rect 17144 42242 17172 42774
rect 17052 42214 17172 42242
rect 16948 42152 17000 42158
rect 16948 42094 17000 42100
rect 17052 41070 17080 42214
rect 17236 42090 17264 43046
rect 17420 42770 17448 43064
rect 17592 43046 17644 43052
rect 17776 43104 17828 43110
rect 17776 43046 17828 43052
rect 17960 43104 18012 43110
rect 17960 43046 18012 43052
rect 17408 42764 17460 42770
rect 17408 42706 17460 42712
rect 17316 42356 17368 42362
rect 17316 42298 17368 42304
rect 17224 42084 17276 42090
rect 17224 42026 17276 42032
rect 17132 41812 17184 41818
rect 17132 41754 17184 41760
rect 17144 41138 17172 41754
rect 17328 41274 17356 42298
rect 17420 42265 17448 42706
rect 17500 42560 17552 42566
rect 17500 42502 17552 42508
rect 17406 42256 17462 42265
rect 17406 42191 17462 42200
rect 17316 41268 17368 41274
rect 17316 41210 17368 41216
rect 17132 41132 17184 41138
rect 17132 41074 17184 41080
rect 17040 41064 17092 41070
rect 17040 41006 17092 41012
rect 16764 40588 16816 40594
rect 16868 40582 16988 40610
rect 16764 40530 16816 40536
rect 16856 40520 16908 40526
rect 16856 40462 16908 40468
rect 16764 40452 16816 40458
rect 16764 40394 16816 40400
rect 16776 40118 16804 40394
rect 16868 40186 16896 40462
rect 16856 40180 16908 40186
rect 16856 40122 16908 40128
rect 16764 40112 16816 40118
rect 16764 40054 16816 40060
rect 16672 40044 16724 40050
rect 16672 39986 16724 39992
rect 16960 39982 16988 40582
rect 16580 39976 16632 39982
rect 16580 39918 16632 39924
rect 16948 39976 17000 39982
rect 16948 39918 17000 39924
rect 16396 39840 16448 39846
rect 16396 39782 16448 39788
rect 16488 39840 16540 39846
rect 16488 39782 16540 39788
rect 16672 39840 16724 39846
rect 16672 39782 16724 39788
rect 16224 38950 16344 38978
rect 16224 38894 16252 38950
rect 16212 38888 16264 38894
rect 16212 38830 16264 38836
rect 16212 38752 16264 38758
rect 16212 38694 16264 38700
rect 16224 38418 16252 38694
rect 16316 38536 16344 38950
rect 16408 38706 16436 39782
rect 16500 39574 16528 39782
rect 16488 39568 16540 39574
rect 16488 39510 16540 39516
rect 16500 38894 16528 39510
rect 16488 38888 16540 38894
rect 16488 38830 16540 38836
rect 16684 38758 16712 39782
rect 16960 39098 16988 39918
rect 16948 39092 17000 39098
rect 16948 39034 17000 39040
rect 16960 38962 16988 39034
rect 16948 38956 17000 38962
rect 16948 38898 17000 38904
rect 16948 38820 17000 38826
rect 16948 38762 17000 38768
rect 16672 38752 16724 38758
rect 16408 38678 16528 38706
rect 16672 38694 16724 38700
rect 16856 38752 16908 38758
rect 16856 38694 16908 38700
rect 16396 38548 16448 38554
rect 16316 38508 16396 38536
rect 16396 38490 16448 38496
rect 16028 38412 16080 38418
rect 16028 38354 16080 38360
rect 16212 38412 16264 38418
rect 16212 38354 16264 38360
rect 15936 38344 15988 38350
rect 15936 38286 15988 38292
rect 15948 38010 15976 38286
rect 15936 38004 15988 38010
rect 15936 37946 15988 37952
rect 15844 37800 15896 37806
rect 15844 37742 15896 37748
rect 16040 36718 16068 38354
rect 16120 38276 16172 38282
rect 16120 38218 16172 38224
rect 16132 36854 16160 38218
rect 16212 37800 16264 37806
rect 16212 37742 16264 37748
rect 16224 36922 16252 37742
rect 16408 37738 16436 38490
rect 16500 37942 16528 38678
rect 16488 37936 16540 37942
rect 16488 37878 16540 37884
rect 16396 37732 16448 37738
rect 16396 37674 16448 37680
rect 16500 37618 16528 37878
rect 16408 37590 16528 37618
rect 16408 37330 16436 37590
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16396 37324 16448 37330
rect 16396 37266 16448 37272
rect 16212 36916 16264 36922
rect 16212 36858 16264 36864
rect 16120 36848 16172 36854
rect 16120 36790 16172 36796
rect 16028 36712 16080 36718
rect 16028 36654 16080 36660
rect 16040 36378 16068 36654
rect 16132 36582 16160 36790
rect 16396 36780 16448 36786
rect 16396 36722 16448 36728
rect 16212 36644 16264 36650
rect 16212 36586 16264 36592
rect 16120 36576 16172 36582
rect 16120 36518 16172 36524
rect 16028 36372 16080 36378
rect 16028 36314 16080 36320
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 16040 35698 16068 36314
rect 16224 36242 16252 36586
rect 16408 36394 16436 36722
rect 16500 36718 16528 37402
rect 16488 36712 16540 36718
rect 16488 36654 16540 36660
rect 16408 36366 16528 36394
rect 16212 36236 16264 36242
rect 16396 36236 16448 36242
rect 16264 36196 16396 36224
rect 16212 36178 16264 36184
rect 16028 35692 16080 35698
rect 16028 35634 16080 35640
rect 15660 35624 15712 35630
rect 15660 35566 15712 35572
rect 16212 35624 16264 35630
rect 16212 35566 16264 35572
rect 15476 34060 15528 34066
rect 15476 34002 15528 34008
rect 15568 34060 15620 34066
rect 15568 34002 15620 34008
rect 15384 33856 15436 33862
rect 15384 33798 15436 33804
rect 15580 33590 15608 34002
rect 15568 33584 15620 33590
rect 15568 33526 15620 33532
rect 15292 33516 15344 33522
rect 15292 33458 15344 33464
rect 15200 33040 15252 33046
rect 15200 32982 15252 32988
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 14924 32292 14976 32298
rect 14924 32234 14976 32240
rect 14936 32026 14964 32234
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 15212 31890 15240 32778
rect 15304 31890 15332 33458
rect 15384 32972 15436 32978
rect 15384 32914 15436 32920
rect 15396 32570 15424 32914
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15672 32230 15700 35566
rect 16224 35290 16252 35566
rect 16212 35284 16264 35290
rect 16212 35226 16264 35232
rect 16028 35012 16080 35018
rect 16028 34954 16080 34960
rect 16040 34542 16068 34954
rect 16028 34536 16080 34542
rect 16028 34478 16080 34484
rect 16316 34066 16344 36196
rect 16396 36178 16448 36184
rect 16500 36174 16528 36366
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16396 36032 16448 36038
rect 16396 35974 16448 35980
rect 16488 36032 16540 36038
rect 16488 35974 16540 35980
rect 16408 35154 16436 35974
rect 16500 35766 16528 35974
rect 16488 35760 16540 35766
rect 16488 35702 16540 35708
rect 16488 35624 16540 35630
rect 16488 35566 16540 35572
rect 16500 35494 16528 35566
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 16396 35148 16448 35154
rect 16396 35090 16448 35096
rect 16500 34746 16528 35430
rect 16488 34740 16540 34746
rect 16488 34682 16540 34688
rect 16684 34610 16712 38694
rect 16868 38010 16896 38694
rect 16856 38004 16908 38010
rect 16856 37946 16908 37952
rect 16960 37806 16988 38762
rect 16948 37800 17000 37806
rect 16948 37742 17000 37748
rect 16856 37664 16908 37670
rect 16856 37606 16908 37612
rect 16868 36242 16896 37606
rect 16960 37330 16988 37742
rect 16948 37324 17000 37330
rect 16948 37266 17000 37272
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 16764 35624 16816 35630
rect 16764 35566 16816 35572
rect 16776 35290 16804 35566
rect 16764 35284 16816 35290
rect 16764 35226 16816 35232
rect 16960 35154 16988 37266
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 16500 34190 16804 34218
rect 16304 34060 16356 34066
rect 16304 34002 16356 34008
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 16028 32972 16080 32978
rect 16028 32914 16080 32920
rect 15844 32564 15896 32570
rect 15844 32506 15896 32512
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15672 31890 15700 32166
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15292 31884 15344 31890
rect 15292 31826 15344 31832
rect 15660 31884 15712 31890
rect 15660 31826 15712 31832
rect 15752 31884 15804 31890
rect 15752 31826 15804 31832
rect 15212 31278 15240 31826
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15304 30870 15332 31826
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15292 30864 15344 30870
rect 15292 30806 15344 30812
rect 15304 29238 15332 30806
rect 15396 30258 15424 31214
rect 15568 30796 15620 30802
rect 15568 30738 15620 30744
rect 15580 30394 15608 30738
rect 15568 30388 15620 30394
rect 15568 30330 15620 30336
rect 15384 30252 15436 30258
rect 15384 30194 15436 30200
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 15672 29102 15700 31826
rect 15764 31142 15792 31826
rect 15856 31754 15884 32506
rect 16040 32366 16068 32914
rect 16132 32570 16160 33798
rect 16500 33046 16528 34190
rect 16776 34134 16804 34190
rect 16764 34128 16816 34134
rect 16764 34070 16816 34076
rect 16580 34060 16632 34066
rect 16580 34002 16632 34008
rect 16592 33046 16620 34002
rect 16948 33924 17000 33930
rect 16948 33866 17000 33872
rect 16856 33856 16908 33862
rect 16856 33798 16908 33804
rect 16764 33584 16816 33590
rect 16764 33526 16816 33532
rect 16672 33448 16724 33454
rect 16672 33390 16724 33396
rect 16684 33114 16712 33390
rect 16776 33130 16804 33526
rect 16868 33522 16896 33798
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16776 33114 16896 33130
rect 16672 33108 16724 33114
rect 16776 33108 16908 33114
rect 16776 33102 16856 33108
rect 16672 33050 16724 33056
rect 16856 33050 16908 33056
rect 16488 33040 16540 33046
rect 16488 32982 16540 32988
rect 16580 33040 16632 33046
rect 16580 32982 16632 32988
rect 16960 32910 16988 33866
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 16120 32564 16172 32570
rect 16120 32506 16172 32512
rect 16132 32434 16160 32506
rect 16120 32428 16172 32434
rect 16120 32370 16172 32376
rect 16028 32360 16080 32366
rect 16028 32302 16080 32308
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15948 31958 15976 32166
rect 15936 31952 15988 31958
rect 15936 31894 15988 31900
rect 15856 31726 15976 31754
rect 15948 31278 15976 31726
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15936 31272 15988 31278
rect 15936 31214 15988 31220
rect 16120 31272 16172 31278
rect 16120 31214 16172 31220
rect 15752 31136 15804 31142
rect 15752 31078 15804 31084
rect 15856 30938 15884 31214
rect 15844 30932 15896 30938
rect 15844 30874 15896 30880
rect 16132 30054 16160 31214
rect 16316 30938 16344 32846
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16408 30818 16436 32370
rect 16684 31958 16712 32506
rect 16776 32298 16804 32778
rect 17052 32774 17080 41006
rect 17144 40594 17172 41074
rect 17408 40996 17460 41002
rect 17408 40938 17460 40944
rect 17316 40928 17368 40934
rect 17316 40870 17368 40876
rect 17224 40724 17276 40730
rect 17224 40666 17276 40672
rect 17132 40588 17184 40594
rect 17132 40530 17184 40536
rect 17132 39976 17184 39982
rect 17132 39918 17184 39924
rect 17144 39574 17172 39918
rect 17132 39568 17184 39574
rect 17132 39510 17184 39516
rect 17236 38978 17264 40666
rect 17328 40610 17356 40870
rect 17420 40730 17448 40938
rect 17408 40724 17460 40730
rect 17408 40666 17460 40672
rect 17328 40582 17448 40610
rect 17316 40520 17368 40526
rect 17316 40462 17368 40468
rect 17328 39846 17356 40462
rect 17420 40390 17448 40582
rect 17512 40390 17540 42502
rect 17604 41478 17632 43046
rect 17592 41472 17644 41478
rect 17592 41414 17644 41420
rect 17604 41138 17632 41414
rect 17592 41132 17644 41138
rect 17592 41074 17644 41080
rect 17592 40996 17644 41002
rect 17592 40938 17644 40944
rect 17604 40662 17632 40938
rect 17788 40662 17816 43046
rect 17972 42945 18000 43046
rect 17958 42936 18014 42945
rect 17958 42871 18014 42880
rect 17972 42770 18000 42871
rect 18156 42838 18184 43114
rect 18144 42832 18196 42838
rect 18144 42774 18196 42780
rect 17960 42764 18012 42770
rect 17960 42706 18012 42712
rect 18326 42256 18382 42265
rect 18326 42191 18382 42200
rect 18340 42022 18368 42191
rect 18524 42158 18552 43132
rect 18696 42356 18748 42362
rect 18696 42298 18748 42304
rect 18708 42158 18736 42298
rect 18512 42152 18564 42158
rect 18512 42094 18564 42100
rect 18696 42152 18748 42158
rect 18696 42094 18748 42100
rect 18144 42016 18196 42022
rect 18144 41958 18196 41964
rect 18328 42016 18380 42022
rect 18328 41958 18380 41964
rect 17868 41676 17920 41682
rect 17868 41618 17920 41624
rect 17880 41070 17908 41618
rect 18156 41274 18184 41958
rect 18524 41818 18552 42094
rect 18512 41812 18564 41818
rect 18512 41754 18564 41760
rect 18800 41414 18828 43200
rect 18880 43182 18932 43188
rect 19154 43208 19210 43217
rect 19154 43143 19156 43152
rect 19208 43143 19210 43152
rect 19156 43114 19208 43120
rect 19168 43058 19196 43114
rect 18616 41386 18828 41414
rect 18892 43030 19196 43058
rect 18144 41268 18196 41274
rect 18144 41210 18196 41216
rect 17868 41064 17920 41070
rect 17868 41006 17920 41012
rect 17960 41064 18012 41070
rect 17960 41006 18012 41012
rect 17972 40882 18000 41006
rect 17880 40854 18000 40882
rect 18052 40928 18104 40934
rect 18052 40870 18104 40876
rect 17592 40656 17644 40662
rect 17592 40598 17644 40604
rect 17776 40656 17828 40662
rect 17776 40598 17828 40604
rect 17684 40452 17736 40458
rect 17684 40394 17736 40400
rect 17408 40384 17460 40390
rect 17408 40326 17460 40332
rect 17500 40384 17552 40390
rect 17500 40326 17552 40332
rect 17420 39982 17448 40326
rect 17408 39976 17460 39982
rect 17408 39918 17460 39924
rect 17316 39840 17368 39846
rect 17316 39782 17368 39788
rect 17144 38950 17264 38978
rect 17144 35834 17172 38950
rect 17328 38894 17356 39782
rect 17224 38888 17276 38894
rect 17224 38830 17276 38836
rect 17316 38888 17368 38894
rect 17316 38830 17368 38836
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 17236 34950 17264 38830
rect 17420 35018 17448 39918
rect 17696 39642 17724 40394
rect 17880 40186 17908 40854
rect 17960 40588 18012 40594
rect 18064 40576 18092 40870
rect 18012 40548 18092 40576
rect 17960 40530 18012 40536
rect 17868 40180 17920 40186
rect 17868 40122 17920 40128
rect 18156 40118 18184 41210
rect 18616 40662 18644 41386
rect 18420 40656 18472 40662
rect 18420 40598 18472 40604
rect 18604 40656 18656 40662
rect 18604 40598 18656 40604
rect 17776 40112 17828 40118
rect 17776 40054 17828 40060
rect 18144 40112 18196 40118
rect 18144 40054 18196 40060
rect 17684 39636 17736 39642
rect 17684 39578 17736 39584
rect 17696 38418 17724 39578
rect 17788 39370 17816 40054
rect 17776 39364 17828 39370
rect 17776 39306 17828 39312
rect 17684 38412 17736 38418
rect 17684 38354 17736 38360
rect 17500 38344 17552 38350
rect 17500 38286 17552 38292
rect 17408 35012 17460 35018
rect 17408 34954 17460 34960
rect 17224 34944 17276 34950
rect 17224 34886 17276 34892
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 17144 33386 17172 33594
rect 17132 33380 17184 33386
rect 17132 33322 17184 33328
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 17512 32366 17540 38286
rect 17696 37942 17724 38354
rect 17684 37936 17736 37942
rect 17684 37878 17736 37884
rect 17788 37754 17816 39306
rect 18432 39302 18460 40598
rect 18892 40594 18920 43030
rect 19536 42770 19564 43250
rect 19628 43246 19656 43279
rect 19616 43240 19668 43246
rect 19616 43182 19668 43188
rect 19616 43104 19668 43110
rect 19616 43046 19668 43052
rect 19628 42786 19656 43046
rect 19720 42906 19748 43726
rect 21456 43648 21508 43654
rect 21456 43590 21508 43596
rect 19800 43240 19852 43246
rect 19800 43182 19852 43188
rect 19708 42900 19760 42906
rect 19708 42842 19760 42848
rect 19524 42764 19576 42770
rect 19628 42758 19748 42786
rect 19524 42706 19576 42712
rect 19616 42628 19668 42634
rect 19616 42570 19668 42576
rect 18972 42560 19024 42566
rect 19156 42560 19208 42566
rect 18972 42502 19024 42508
rect 19076 42520 19156 42548
rect 18984 42294 19012 42502
rect 18972 42288 19024 42294
rect 18972 42230 19024 42236
rect 19076 42158 19104 42520
rect 19156 42502 19208 42508
rect 19210 42460 19518 42469
rect 19210 42458 19216 42460
rect 19272 42458 19296 42460
rect 19352 42458 19376 42460
rect 19432 42458 19456 42460
rect 19512 42458 19518 42460
rect 19272 42406 19274 42458
rect 19454 42406 19456 42458
rect 19210 42404 19216 42406
rect 19272 42404 19296 42406
rect 19352 42404 19376 42406
rect 19432 42404 19456 42406
rect 19512 42404 19518 42406
rect 19210 42395 19518 42404
rect 19628 42362 19656 42570
rect 19432 42356 19484 42362
rect 19432 42298 19484 42304
rect 19616 42356 19668 42362
rect 19616 42298 19668 42304
rect 19154 42256 19210 42265
rect 19154 42191 19210 42200
rect 19168 42158 19196 42191
rect 19064 42152 19116 42158
rect 19064 42094 19116 42100
rect 19156 42152 19208 42158
rect 19444 42106 19472 42298
rect 19720 42242 19748 42758
rect 19536 42214 19748 42242
rect 19536 42158 19564 42214
rect 19156 42094 19208 42100
rect 19076 41274 19104 42094
rect 19352 42090 19472 42106
rect 19524 42152 19576 42158
rect 19708 42152 19760 42158
rect 19524 42094 19576 42100
rect 19628 42112 19708 42140
rect 19340 42084 19472 42090
rect 19392 42078 19472 42084
rect 19340 42026 19392 42032
rect 19628 41614 19656 42112
rect 19708 42094 19760 42100
rect 19812 42090 19840 43182
rect 20260 43104 20312 43110
rect 20260 43046 20312 43052
rect 20352 43104 20404 43110
rect 20352 43046 20404 43052
rect 21088 43104 21140 43110
rect 21088 43046 21140 43052
rect 21272 43104 21324 43110
rect 21272 43046 21324 43052
rect 19870 43004 20178 43013
rect 19870 43002 19876 43004
rect 19932 43002 19956 43004
rect 20012 43002 20036 43004
rect 20092 43002 20116 43004
rect 20172 43002 20178 43004
rect 19932 42950 19934 43002
rect 20114 42950 20116 43002
rect 19870 42948 19876 42950
rect 19932 42948 19956 42950
rect 20012 42948 20036 42950
rect 20092 42948 20116 42950
rect 20172 42948 20178 42950
rect 19870 42939 20178 42948
rect 20272 42770 20300 43046
rect 20364 42770 20392 43046
rect 20536 42832 20588 42838
rect 20536 42774 20588 42780
rect 20076 42764 20128 42770
rect 20076 42706 20128 42712
rect 20260 42764 20312 42770
rect 20260 42706 20312 42712
rect 20352 42764 20404 42770
rect 20352 42706 20404 42712
rect 20088 42294 20116 42706
rect 20076 42288 20128 42294
rect 20076 42230 20128 42236
rect 20260 42152 20312 42158
rect 20260 42094 20312 42100
rect 19800 42084 19852 42090
rect 19800 42026 19852 42032
rect 19616 41608 19668 41614
rect 19616 41550 19668 41556
rect 19210 41372 19518 41381
rect 19210 41370 19216 41372
rect 19272 41370 19296 41372
rect 19352 41370 19376 41372
rect 19432 41370 19456 41372
rect 19512 41370 19518 41372
rect 19272 41318 19274 41370
rect 19454 41318 19456 41370
rect 19210 41316 19216 41318
rect 19272 41316 19296 41318
rect 19352 41316 19376 41318
rect 19432 41316 19456 41318
rect 19512 41316 19518 41318
rect 19210 41307 19518 41316
rect 19064 41268 19116 41274
rect 19064 41210 19116 41216
rect 19340 41064 19392 41070
rect 19340 41006 19392 41012
rect 19524 41064 19576 41070
rect 19628 41052 19656 41550
rect 19576 41024 19656 41052
rect 19708 41064 19760 41070
rect 19524 41006 19576 41012
rect 19708 41006 19760 41012
rect 19248 40996 19300 41002
rect 19248 40938 19300 40944
rect 19260 40730 19288 40938
rect 19248 40724 19300 40730
rect 19248 40666 19300 40672
rect 19352 40594 19380 41006
rect 18880 40588 18932 40594
rect 18880 40530 18932 40536
rect 19340 40588 19392 40594
rect 19340 40530 19392 40536
rect 19616 40588 19668 40594
rect 19616 40530 19668 40536
rect 18696 40384 18748 40390
rect 18696 40326 18748 40332
rect 18708 39506 18736 40326
rect 18892 40050 18920 40530
rect 19064 40452 19116 40458
rect 19064 40394 19116 40400
rect 18880 40044 18932 40050
rect 18880 39986 18932 39992
rect 18972 39976 19024 39982
rect 18972 39918 19024 39924
rect 18984 39642 19012 39918
rect 18972 39636 19024 39642
rect 18972 39578 19024 39584
rect 18512 39500 18564 39506
rect 18512 39442 18564 39448
rect 18696 39500 18748 39506
rect 18696 39442 18748 39448
rect 18880 39500 18932 39506
rect 18880 39442 18932 39448
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18432 38826 18460 39238
rect 18524 39098 18552 39442
rect 18892 39370 18920 39442
rect 18880 39364 18932 39370
rect 18880 39306 18932 39312
rect 18512 39092 18564 39098
rect 18512 39034 18564 39040
rect 18420 38820 18472 38826
rect 18420 38762 18472 38768
rect 18432 38418 18460 38762
rect 19076 38418 19104 40394
rect 19210 40284 19518 40293
rect 19210 40282 19216 40284
rect 19272 40282 19296 40284
rect 19352 40282 19376 40284
rect 19432 40282 19456 40284
rect 19512 40282 19518 40284
rect 19272 40230 19274 40282
rect 19454 40230 19456 40282
rect 19210 40228 19216 40230
rect 19272 40228 19296 40230
rect 19352 40228 19376 40230
rect 19432 40228 19456 40230
rect 19512 40228 19518 40230
rect 19210 40219 19518 40228
rect 19628 39506 19656 40530
rect 19720 39964 19748 41006
rect 19812 40594 19840 42026
rect 19870 41916 20178 41925
rect 19870 41914 19876 41916
rect 19932 41914 19956 41916
rect 20012 41914 20036 41916
rect 20092 41914 20116 41916
rect 20172 41914 20178 41916
rect 19932 41862 19934 41914
rect 20114 41862 20116 41914
rect 19870 41860 19876 41862
rect 19932 41860 19956 41862
rect 20012 41860 20036 41862
rect 20092 41860 20116 41862
rect 20172 41860 20178 41862
rect 19870 41851 20178 41860
rect 20076 41812 20128 41818
rect 20076 41754 20128 41760
rect 20088 41002 20116 41754
rect 20272 41750 20300 42094
rect 20364 42022 20392 42706
rect 20352 42016 20404 42022
rect 20352 41958 20404 41964
rect 20444 42016 20496 42022
rect 20444 41958 20496 41964
rect 20260 41744 20312 41750
rect 20260 41686 20312 41692
rect 20364 41414 20392 41958
rect 20456 41614 20484 41958
rect 20444 41608 20496 41614
rect 20444 41550 20496 41556
rect 20272 41386 20392 41414
rect 20272 41070 20300 41386
rect 20352 41268 20404 41274
rect 20352 41210 20404 41216
rect 20364 41070 20392 41210
rect 20456 41070 20484 41550
rect 20548 41478 20576 42774
rect 21100 42226 21128 43046
rect 21284 42770 21312 43046
rect 21272 42764 21324 42770
rect 21272 42706 21324 42712
rect 21364 42764 21416 42770
rect 21364 42706 21416 42712
rect 21376 42362 21404 42706
rect 21364 42356 21416 42362
rect 21364 42298 21416 42304
rect 21088 42220 21140 42226
rect 21088 42162 21140 42168
rect 20812 42152 20864 42158
rect 20812 42094 20864 42100
rect 20996 42152 21048 42158
rect 20996 42094 21048 42100
rect 20536 41472 20588 41478
rect 20536 41414 20588 41420
rect 20260 41064 20312 41070
rect 20260 41006 20312 41012
rect 20352 41064 20404 41070
rect 20352 41006 20404 41012
rect 20444 41064 20496 41070
rect 20444 41006 20496 41012
rect 20076 40996 20128 41002
rect 20076 40938 20128 40944
rect 19870 40828 20178 40837
rect 19870 40826 19876 40828
rect 19932 40826 19956 40828
rect 20012 40826 20036 40828
rect 20092 40826 20116 40828
rect 20172 40826 20178 40828
rect 19932 40774 19934 40826
rect 20114 40774 20116 40826
rect 19870 40772 19876 40774
rect 19932 40772 19956 40774
rect 20012 40772 20036 40774
rect 20092 40772 20116 40774
rect 20172 40772 20178 40774
rect 19870 40763 20178 40772
rect 19800 40588 19852 40594
rect 19800 40530 19852 40536
rect 19800 39976 19852 39982
rect 19720 39936 19800 39964
rect 19800 39918 19852 39924
rect 19248 39500 19300 39506
rect 19248 39442 19300 39448
rect 19616 39500 19668 39506
rect 19616 39442 19668 39448
rect 19260 39302 19288 39442
rect 19248 39296 19300 39302
rect 19248 39238 19300 39244
rect 19210 39196 19518 39205
rect 19210 39194 19216 39196
rect 19272 39194 19296 39196
rect 19352 39194 19376 39196
rect 19432 39194 19456 39196
rect 19512 39194 19518 39196
rect 19272 39142 19274 39194
rect 19454 39142 19456 39194
rect 19210 39140 19216 39142
rect 19272 39140 19296 39142
rect 19352 39140 19376 39142
rect 19432 39140 19456 39142
rect 19512 39140 19518 39142
rect 19210 39131 19518 39140
rect 19432 39092 19484 39098
rect 19432 39034 19484 39040
rect 18420 38412 18472 38418
rect 18420 38354 18472 38360
rect 19064 38412 19116 38418
rect 19064 38354 19116 38360
rect 18972 38344 19024 38350
rect 18972 38286 19024 38292
rect 17868 38208 17920 38214
rect 17868 38150 17920 38156
rect 17880 37874 17908 38150
rect 18052 38004 18104 38010
rect 18052 37946 18104 37952
rect 18880 38004 18932 38010
rect 18880 37946 18932 37952
rect 17868 37868 17920 37874
rect 17868 37810 17920 37816
rect 17788 37726 17908 37754
rect 17880 37670 17908 37726
rect 17868 37664 17920 37670
rect 17868 37606 17920 37612
rect 17880 36922 17908 37606
rect 17868 36916 17920 36922
rect 17868 36858 17920 36864
rect 17960 36644 18012 36650
rect 17960 36586 18012 36592
rect 17972 36378 18000 36586
rect 17960 36372 18012 36378
rect 17960 36314 18012 36320
rect 17972 36242 18000 36314
rect 17960 36236 18012 36242
rect 17960 36178 18012 36184
rect 18064 35086 18092 37946
rect 18328 37800 18380 37806
rect 18328 37742 18380 37748
rect 18340 37618 18368 37742
rect 18892 37738 18920 37946
rect 18984 37806 19012 38286
rect 18972 37800 19024 37806
rect 18972 37742 19024 37748
rect 18788 37732 18840 37738
rect 18788 37674 18840 37680
rect 18880 37732 18932 37738
rect 18880 37674 18932 37680
rect 18248 37590 18368 37618
rect 18144 36576 18196 36582
rect 18144 36518 18196 36524
rect 18156 36174 18184 36518
rect 18144 36168 18196 36174
rect 18144 36110 18196 36116
rect 18156 35494 18184 36110
rect 18144 35488 18196 35494
rect 18144 35430 18196 35436
rect 18052 35080 18104 35086
rect 18052 35022 18104 35028
rect 18064 34610 18092 35022
rect 18052 34604 18104 34610
rect 18052 34546 18104 34552
rect 18144 34604 18196 34610
rect 18144 34546 18196 34552
rect 17960 34536 18012 34542
rect 17960 34478 18012 34484
rect 17972 33998 18000 34478
rect 18064 34082 18092 34546
rect 18156 34202 18184 34546
rect 18248 34406 18276 37590
rect 18800 37380 18828 37674
rect 18880 37392 18932 37398
rect 18800 37352 18880 37380
rect 18880 37334 18932 37340
rect 18328 37120 18380 37126
rect 18328 37062 18380 37068
rect 18604 37120 18656 37126
rect 18604 37062 18656 37068
rect 18340 36174 18368 37062
rect 18420 36236 18472 36242
rect 18420 36178 18472 36184
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 18236 34400 18288 34406
rect 18236 34342 18288 34348
rect 18248 34202 18276 34342
rect 18144 34196 18196 34202
rect 18144 34138 18196 34144
rect 18236 34196 18288 34202
rect 18236 34138 18288 34144
rect 18064 34054 18184 34082
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 17696 32570 17724 32846
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 17972 32366 18000 33934
rect 18064 33454 18092 33934
rect 18156 33454 18184 34054
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 18144 33448 18196 33454
rect 18144 33390 18196 33396
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17316 32360 17368 32366
rect 17500 32360 17552 32366
rect 17368 32320 17500 32348
rect 17316 32302 17368 32308
rect 17500 32302 17552 32308
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 16764 32292 16816 32298
rect 16764 32234 16816 32240
rect 16948 32292 17000 32298
rect 16948 32234 17000 32240
rect 16776 32026 16804 32234
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 16672 31952 16724 31958
rect 16670 31920 16672 31929
rect 16724 31920 16726 31929
rect 16670 31855 16726 31864
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16224 30790 16436 30818
rect 16500 30802 16528 31078
rect 16592 30870 16620 31214
rect 16580 30864 16632 30870
rect 16580 30806 16632 30812
rect 16488 30796 16540 30802
rect 16224 30326 16252 30790
rect 16488 30738 16540 30744
rect 16304 30660 16356 30666
rect 16304 30602 16356 30608
rect 16212 30320 16264 30326
rect 16212 30262 16264 30268
rect 16212 30184 16264 30190
rect 16316 30138 16344 30602
rect 16396 30592 16448 30598
rect 16396 30534 16448 30540
rect 16408 30190 16436 30534
rect 16488 30320 16540 30326
rect 16488 30262 16540 30268
rect 16264 30132 16344 30138
rect 16212 30126 16344 30132
rect 16396 30184 16448 30190
rect 16396 30126 16448 30132
rect 16224 30110 16344 30126
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 15936 29708 15988 29714
rect 15936 29650 15988 29656
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 15108 28688 15160 28694
rect 15108 28630 15160 28636
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14476 27674 14504 28494
rect 14568 28218 14596 28494
rect 14556 28212 14608 28218
rect 14556 28154 14608 28160
rect 15120 28014 15148 28630
rect 15948 28558 15976 29650
rect 16120 29504 16172 29510
rect 16120 29446 16172 29452
rect 16132 29170 16160 29446
rect 16224 29238 16252 30110
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16212 29232 16264 29238
rect 16212 29174 16264 29180
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16224 28642 16252 29174
rect 16316 28762 16344 29990
rect 16304 28756 16356 28762
rect 16304 28698 16356 28704
rect 16224 28626 16344 28642
rect 16224 28620 16356 28626
rect 16224 28614 16304 28620
rect 16304 28562 16356 28568
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15948 28150 15976 28494
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 16120 28144 16172 28150
rect 16120 28086 16172 28092
rect 16132 28014 16160 28086
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 16120 28008 16172 28014
rect 16120 27950 16172 27956
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 15120 27606 15148 27950
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 15108 27600 15160 27606
rect 15108 27542 15160 27548
rect 14740 27532 14792 27538
rect 14740 27474 14792 27480
rect 14280 27396 14332 27402
rect 14280 27338 14332 27344
rect 14292 26926 14320 27338
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14556 26920 14608 26926
rect 14556 26862 14608 26868
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 13820 26580 13872 26586
rect 13820 26522 13872 26528
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 11436 26140 11744 26149
rect 11436 26138 11442 26140
rect 11498 26138 11522 26140
rect 11578 26138 11602 26140
rect 11658 26138 11682 26140
rect 11738 26138 11744 26140
rect 11498 26086 11500 26138
rect 11680 26086 11682 26138
rect 11436 26084 11442 26086
rect 11498 26084 11522 26086
rect 11578 26084 11602 26086
rect 11658 26084 11682 26086
rect 11738 26084 11744 26086
rect 11436 26075 11744 26084
rect 12636 25906 12664 26318
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 11336 25832 11388 25838
rect 11256 25792 11336 25820
rect 11336 25774 11388 25780
rect 4322 25596 4630 25605
rect 4322 25594 4328 25596
rect 4384 25594 4408 25596
rect 4464 25594 4488 25596
rect 4544 25594 4568 25596
rect 4624 25594 4630 25596
rect 4384 25542 4386 25594
rect 4566 25542 4568 25594
rect 4322 25540 4328 25542
rect 4384 25540 4408 25542
rect 4464 25540 4488 25542
rect 4544 25540 4568 25542
rect 4624 25540 4630 25542
rect 4322 25531 4630 25540
rect 3662 25052 3970 25061
rect 3662 25050 3668 25052
rect 3724 25050 3748 25052
rect 3804 25050 3828 25052
rect 3884 25050 3908 25052
rect 3964 25050 3970 25052
rect 3724 24998 3726 25050
rect 3906 24998 3908 25050
rect 3662 24996 3668 24998
rect 3724 24996 3748 24998
rect 3804 24996 3828 24998
rect 3884 24996 3908 24998
rect 3964 24996 3970 24998
rect 3662 24987 3970 24996
rect 11348 24750 11376 25774
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11900 25362 11928 25638
rect 12096 25596 12404 25605
rect 12096 25594 12102 25596
rect 12158 25594 12182 25596
rect 12238 25594 12262 25596
rect 12318 25594 12342 25596
rect 12398 25594 12404 25596
rect 12158 25542 12160 25594
rect 12340 25542 12342 25594
rect 12096 25540 12102 25542
rect 12158 25540 12182 25542
rect 12238 25540 12262 25542
rect 12318 25540 12342 25542
rect 12398 25540 12404 25542
rect 12096 25531 12404 25540
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11436 25052 11744 25061
rect 11436 25050 11442 25052
rect 11498 25050 11522 25052
rect 11578 25050 11602 25052
rect 11658 25050 11682 25052
rect 11738 25050 11744 25052
rect 11498 24998 11500 25050
rect 11680 24998 11682 25050
rect 11436 24996 11442 24998
rect 11498 24996 11522 24998
rect 11578 24996 11602 24998
rect 11658 24996 11682 24998
rect 11738 24996 11744 24998
rect 11436 24987 11744 24996
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 4322 24508 4630 24517
rect 4322 24506 4328 24508
rect 4384 24506 4408 24508
rect 4464 24506 4488 24508
rect 4544 24506 4568 24508
rect 4624 24506 4630 24508
rect 4384 24454 4386 24506
rect 4566 24454 4568 24506
rect 4322 24452 4328 24454
rect 4384 24452 4408 24454
rect 4464 24452 4488 24454
rect 4544 24452 4568 24454
rect 4624 24452 4630 24454
rect 4322 24443 4630 24452
rect 3662 23964 3970 23973
rect 3662 23962 3668 23964
rect 3724 23962 3748 23964
rect 3804 23962 3828 23964
rect 3884 23962 3908 23964
rect 3964 23962 3970 23964
rect 3724 23910 3726 23962
rect 3906 23910 3908 23962
rect 3662 23908 3668 23910
rect 3724 23908 3748 23910
rect 3804 23908 3828 23910
rect 3884 23908 3908 23910
rect 3964 23908 3970 23910
rect 3662 23899 3970 23908
rect 11348 23662 11376 24686
rect 12096 24508 12404 24517
rect 12096 24506 12102 24508
rect 12158 24506 12182 24508
rect 12238 24506 12262 24508
rect 12318 24506 12342 24508
rect 12398 24506 12404 24508
rect 12158 24454 12160 24506
rect 12340 24454 12342 24506
rect 12096 24452 12102 24454
rect 12158 24452 12182 24454
rect 12238 24452 12262 24454
rect 12318 24452 12342 24454
rect 12398 24452 12404 24454
rect 12096 24443 12404 24452
rect 11436 23964 11744 23973
rect 11436 23962 11442 23964
rect 11498 23962 11522 23964
rect 11578 23962 11602 23964
rect 11658 23962 11682 23964
rect 11738 23962 11744 23964
rect 11498 23910 11500 23962
rect 11680 23910 11682 23962
rect 11436 23908 11442 23910
rect 11498 23908 11522 23910
rect 11578 23908 11602 23910
rect 11658 23908 11682 23910
rect 11738 23908 11744 23910
rect 11436 23899 11744 23908
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 4322 23420 4630 23429
rect 4322 23418 4328 23420
rect 4384 23418 4408 23420
rect 4464 23418 4488 23420
rect 4544 23418 4568 23420
rect 4624 23418 4630 23420
rect 4384 23366 4386 23418
rect 4566 23366 4568 23418
rect 4322 23364 4328 23366
rect 4384 23364 4408 23366
rect 4464 23364 4488 23366
rect 4544 23364 4568 23366
rect 4624 23364 4630 23366
rect 4322 23355 4630 23364
rect 12096 23420 12404 23429
rect 12096 23418 12102 23420
rect 12158 23418 12182 23420
rect 12238 23418 12262 23420
rect 12318 23418 12342 23420
rect 12398 23418 12404 23420
rect 12158 23366 12160 23418
rect 12340 23366 12342 23418
rect 12096 23364 12102 23366
rect 12158 23364 12182 23366
rect 12238 23364 12262 23366
rect 12318 23364 12342 23366
rect 12398 23364 12404 23366
rect 12096 23355 12404 23364
rect 12348 23180 12400 23186
rect 12452 23168 12480 23462
rect 12636 23322 12664 25842
rect 12820 25838 12848 26318
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12400 23140 12480 23168
rect 12348 23122 12400 23128
rect 3662 22876 3970 22885
rect 3662 22874 3668 22876
rect 3724 22874 3748 22876
rect 3804 22874 3828 22876
rect 3884 22874 3908 22876
rect 3964 22874 3970 22876
rect 3724 22822 3726 22874
rect 3906 22822 3908 22874
rect 3662 22820 3668 22822
rect 3724 22820 3748 22822
rect 3804 22820 3828 22822
rect 3884 22820 3908 22822
rect 3964 22820 3970 22822
rect 3662 22811 3970 22820
rect 11436 22876 11744 22885
rect 11436 22874 11442 22876
rect 11498 22874 11522 22876
rect 11578 22874 11602 22876
rect 11658 22874 11682 22876
rect 11738 22874 11744 22876
rect 11498 22822 11500 22874
rect 11680 22822 11682 22874
rect 11436 22820 11442 22822
rect 11498 22820 11522 22822
rect 11578 22820 11602 22822
rect 11658 22820 11682 22822
rect 11738 22820 11744 22822
rect 11436 22811 11744 22820
rect 12820 22438 12848 25774
rect 13004 24954 13032 25978
rect 13188 25838 13216 26318
rect 13648 25906 13676 26318
rect 13924 26246 13952 26726
rect 14292 26466 14320 26862
rect 14200 26438 14320 26466
rect 14200 26382 14228 26438
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 14568 26042 14596 26862
rect 14752 26586 14780 27474
rect 15120 27402 15148 27542
rect 15396 27470 15424 27882
rect 15384 27464 15436 27470
rect 15384 27406 15436 27412
rect 15108 27396 15160 27402
rect 15108 27338 15160 27344
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 15292 26512 15344 26518
rect 15292 26454 15344 26460
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15016 26240 15068 26246
rect 15016 26182 15068 26188
rect 14556 26036 14608 26042
rect 14556 25978 14608 25984
rect 15028 25906 15056 26182
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 15212 25838 15240 26318
rect 15304 26042 15332 26454
rect 15396 26042 15424 27406
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 13188 25498 13216 25774
rect 14188 25696 14240 25702
rect 14188 25638 14240 25644
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 15304 25650 15332 25978
rect 15752 25832 15804 25838
rect 15752 25774 15804 25780
rect 15476 25764 15528 25770
rect 15476 25706 15528 25712
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 14200 25430 14228 25638
rect 14188 25424 14240 25430
rect 14188 25366 14240 25372
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 12992 24948 13044 24954
rect 12992 24890 13044 24896
rect 13096 24410 13124 25298
rect 14004 25220 14056 25226
rect 14004 25162 14056 25168
rect 14016 24750 14044 25162
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13740 24274 13768 24550
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23594 13032 24074
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 12992 23588 13044 23594
rect 12992 23530 13044 23536
rect 13004 22506 13032 23530
rect 13648 23322 13676 23734
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 4322 22332 4630 22341
rect 4322 22330 4328 22332
rect 4384 22330 4408 22332
rect 4464 22330 4488 22332
rect 4544 22330 4568 22332
rect 4624 22330 4630 22332
rect 4384 22278 4386 22330
rect 4566 22278 4568 22330
rect 4322 22276 4328 22278
rect 4384 22276 4408 22278
rect 4464 22276 4488 22278
rect 4544 22276 4568 22278
rect 4624 22276 4630 22278
rect 4322 22267 4630 22276
rect 12096 22332 12404 22341
rect 12096 22330 12102 22332
rect 12158 22330 12182 22332
rect 12238 22330 12262 22332
rect 12318 22330 12342 22332
rect 12398 22330 12404 22332
rect 12158 22278 12160 22330
rect 12340 22278 12342 22330
rect 12096 22276 12102 22278
rect 12158 22276 12182 22278
rect 12238 22276 12262 22278
rect 12318 22276 12342 22278
rect 12398 22276 12404 22278
rect 12096 22267 12404 22276
rect 12728 22166 12756 22374
rect 12820 22234 12848 22374
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 11436 21788 11744 21797
rect 11436 21786 11442 21788
rect 11498 21786 11522 21788
rect 11578 21786 11602 21788
rect 11658 21786 11682 21788
rect 11738 21786 11744 21788
rect 11498 21734 11500 21786
rect 11680 21734 11682 21786
rect 11436 21732 11442 21734
rect 11498 21732 11522 21734
rect 11578 21732 11602 21734
rect 11658 21732 11682 21734
rect 11738 21732 11744 21734
rect 11436 21723 11744 21732
rect 13648 21690 13676 22034
rect 13832 21978 13860 24686
rect 13924 24206 13952 24686
rect 14292 24274 14320 25638
rect 15304 25622 15424 25650
rect 15200 25424 15252 25430
rect 15200 25366 15252 25372
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14280 24268 14332 24274
rect 14280 24210 14332 24216
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13924 23254 13952 24142
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 14016 22574 14044 24006
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14200 23186 14228 23666
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13924 22234 13952 22442
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 14016 22098 14044 22374
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 13832 21950 13952 21978
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 12096 21244 12404 21253
rect 12096 21242 12102 21244
rect 12158 21242 12182 21244
rect 12238 21242 12262 21244
rect 12318 21242 12342 21244
rect 12398 21242 12404 21244
rect 12158 21190 12160 21242
rect 12340 21190 12342 21242
rect 12096 21188 12102 21190
rect 12158 21188 12182 21190
rect 12238 21188 12262 21190
rect 12318 21188 12342 21190
rect 12398 21188 12404 21190
rect 12096 21179 12404 21188
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 11436 20700 11744 20709
rect 11436 20698 11442 20700
rect 11498 20698 11522 20700
rect 11578 20698 11602 20700
rect 11658 20698 11682 20700
rect 11738 20698 11744 20700
rect 11498 20646 11500 20698
rect 11680 20646 11682 20698
rect 11436 20644 11442 20646
rect 11498 20644 11522 20646
rect 11578 20644 11602 20646
rect 11658 20644 11682 20646
rect 11738 20644 11744 20646
rect 11436 20635 11744 20644
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 12096 20156 12404 20165
rect 12096 20154 12102 20156
rect 12158 20154 12182 20156
rect 12238 20154 12262 20156
rect 12318 20154 12342 20156
rect 12398 20154 12404 20156
rect 12158 20102 12160 20154
rect 12340 20102 12342 20154
rect 12096 20100 12102 20102
rect 12158 20100 12182 20102
rect 12238 20100 12262 20102
rect 12318 20100 12342 20102
rect 12398 20100 12404 20102
rect 12096 20091 12404 20100
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 11436 19612 11744 19621
rect 11436 19610 11442 19612
rect 11498 19610 11522 19612
rect 11578 19610 11602 19612
rect 11658 19610 11682 19612
rect 11738 19610 11744 19612
rect 11498 19558 11500 19610
rect 11680 19558 11682 19610
rect 11436 19556 11442 19558
rect 11498 19556 11522 19558
rect 11578 19556 11602 19558
rect 11658 19556 11682 19558
rect 11738 19556 11744 19558
rect 11436 19547 11744 19556
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 12096 19068 12404 19077
rect 12096 19066 12102 19068
rect 12158 19066 12182 19068
rect 12238 19066 12262 19068
rect 12318 19066 12342 19068
rect 12398 19066 12404 19068
rect 12158 19014 12160 19066
rect 12340 19014 12342 19066
rect 12096 19012 12102 19014
rect 12158 19012 12182 19014
rect 12238 19012 12262 19014
rect 12318 19012 12342 19014
rect 12398 19012 12404 19014
rect 12096 19003 12404 19012
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 11436 18524 11744 18533
rect 11436 18522 11442 18524
rect 11498 18522 11522 18524
rect 11578 18522 11602 18524
rect 11658 18522 11682 18524
rect 11738 18522 11744 18524
rect 11498 18470 11500 18522
rect 11680 18470 11682 18522
rect 11436 18468 11442 18470
rect 11498 18468 11522 18470
rect 11578 18468 11602 18470
rect 11658 18468 11682 18470
rect 11738 18468 11744 18470
rect 11436 18459 11744 18468
rect 13832 18222 13860 19246
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 12096 17980 12404 17989
rect 12096 17978 12102 17980
rect 12158 17978 12182 17980
rect 12238 17978 12262 17980
rect 12318 17978 12342 17980
rect 12398 17978 12404 17980
rect 12158 17926 12160 17978
rect 12340 17926 12342 17978
rect 12096 17924 12102 17926
rect 12158 17924 12182 17926
rect 12238 17924 12262 17926
rect 12318 17924 12342 17926
rect 12398 17924 12404 17926
rect 12096 17915 12404 17924
rect 13832 17898 13860 18158
rect 13648 17870 13860 17898
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 11436 17436 11744 17445
rect 11436 17434 11442 17436
rect 11498 17434 11522 17436
rect 11578 17434 11602 17436
rect 11658 17434 11682 17436
rect 11738 17434 11744 17436
rect 11498 17382 11500 17434
rect 11680 17382 11682 17434
rect 11436 17380 11442 17382
rect 11498 17380 11522 17382
rect 11578 17380 11602 17382
rect 11658 17380 11682 17382
rect 11738 17380 11744 17382
rect 11436 17371 11744 17380
rect 13648 17134 13676 17870
rect 13924 17746 13952 21950
rect 14108 21486 14136 22646
rect 14292 21894 14320 24210
rect 14384 23662 14412 24686
rect 14660 24342 14688 25094
rect 15016 24676 15068 24682
rect 15016 24618 15068 24624
rect 14648 24336 14700 24342
rect 14648 24278 14700 24284
rect 15028 24070 15056 24618
rect 15212 24138 15240 25366
rect 15396 25294 15424 25622
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15200 24132 15252 24138
rect 15200 24074 15252 24080
rect 15016 24064 15068 24070
rect 15016 24006 15068 24012
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14648 23588 14700 23594
rect 14648 23530 14700 23536
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14384 22506 14412 23258
rect 14660 23186 14688 23530
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 14648 23180 14700 23186
rect 14648 23122 14700 23128
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14384 21554 14412 22442
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14476 22166 14504 22374
rect 14464 22160 14516 22166
rect 14464 22102 14516 22108
rect 14568 21690 14596 22510
rect 14660 22234 14688 23122
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14660 21486 14688 22170
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14844 20058 14872 23054
rect 15212 22574 15240 23462
rect 15304 23254 15332 24550
rect 15292 23248 15344 23254
rect 15292 23190 15344 23196
rect 15304 22574 15332 23190
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15304 22094 15332 22510
rect 15488 22438 15516 25706
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15580 24274 15608 25094
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15764 23322 15792 25774
rect 16224 25362 16252 28426
rect 16316 28014 16344 28562
rect 16408 28218 16436 30126
rect 16500 29714 16528 30262
rect 16592 30190 16620 30806
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 16684 30394 16712 30534
rect 16672 30388 16724 30394
rect 16672 30330 16724 30336
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 16488 29708 16540 29714
rect 16488 29650 16540 29656
rect 16592 29510 16620 30126
rect 16684 29782 16712 30126
rect 16776 29850 16804 31962
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 16868 31414 16896 31758
rect 16960 31686 16988 32234
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17408 32224 17460 32230
rect 17408 32166 17460 32172
rect 17328 32026 17356 32166
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 17420 31754 17448 32166
rect 18052 31884 18104 31890
rect 18052 31826 18104 31832
rect 17132 31748 17184 31754
rect 17132 31690 17184 31696
rect 17328 31726 17448 31754
rect 16948 31680 17000 31686
rect 16948 31622 17000 31628
rect 16856 31408 16908 31414
rect 16856 31350 16908 31356
rect 16868 31278 16896 31350
rect 16856 31272 16908 31278
rect 16856 31214 16908 31220
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16868 30802 16896 31078
rect 16856 30796 16908 30802
rect 16856 30738 16908 30744
rect 16868 30122 16896 30738
rect 16856 30116 16908 30122
rect 16856 30058 16908 30064
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 16672 29776 16724 29782
rect 16672 29718 16724 29724
rect 16488 29504 16540 29510
rect 16488 29446 16540 29452
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 16304 28008 16356 28014
rect 16304 27950 16356 27956
rect 16316 27878 16344 27950
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16316 27674 16344 27814
rect 16304 27668 16356 27674
rect 16304 27610 16356 27616
rect 16500 27470 16528 29446
rect 16592 29016 16620 29446
rect 16684 29306 16712 29718
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16672 29028 16724 29034
rect 16592 28988 16672 29016
rect 16672 28970 16724 28976
rect 16684 28422 16712 28970
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16684 27946 16712 28358
rect 16868 28082 16896 28562
rect 16960 28506 16988 31622
rect 17040 31204 17092 31210
rect 17040 31146 17092 31152
rect 17052 30326 17080 31146
rect 17144 30734 17172 31690
rect 17132 30728 17184 30734
rect 17184 30688 17264 30716
rect 17132 30670 17184 30676
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 17052 29646 17080 30262
rect 17236 30190 17264 30688
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17236 29646 17264 30126
rect 17328 29714 17356 31726
rect 17776 31680 17828 31686
rect 17776 31622 17828 31628
rect 17788 31278 17816 31622
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17776 31272 17828 31278
rect 17960 31272 18012 31278
rect 17776 31214 17828 31220
rect 17880 31232 17960 31260
rect 17408 29776 17460 29782
rect 17408 29718 17460 29724
rect 17316 29708 17368 29714
rect 17316 29650 17368 29656
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 17224 29640 17276 29646
rect 17224 29582 17276 29588
rect 17420 28762 17448 29718
rect 17408 28756 17460 28762
rect 17408 28698 17460 28704
rect 16960 28478 17172 28506
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16672 27940 16724 27946
rect 16672 27882 16724 27888
rect 16776 27606 16804 28018
rect 16764 27600 16816 27606
rect 16764 27542 16816 27548
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16580 26240 16632 26246
rect 16580 26182 16632 26188
rect 16592 25838 16620 26182
rect 16776 26042 16804 26386
rect 16764 26036 16816 26042
rect 16764 25978 16816 25984
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16488 25696 16540 25702
rect 16488 25638 16540 25644
rect 16500 25362 16528 25638
rect 16960 25430 16988 26726
rect 17052 26586 17080 26862
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 17144 26466 17172 28478
rect 17316 27940 17368 27946
rect 17316 27882 17368 27888
rect 17328 27470 17356 27882
rect 17420 27538 17448 28698
rect 17512 28218 17540 31214
rect 17880 30938 17908 31232
rect 17960 31214 18012 31220
rect 18064 31210 18092 31826
rect 18052 31204 18104 31210
rect 18052 31146 18104 31152
rect 18156 30938 18184 33254
rect 18432 32978 18460 36178
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18524 34490 18552 36110
rect 18616 35630 18644 37062
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 18708 36038 18736 36722
rect 18788 36644 18840 36650
rect 18788 36586 18840 36592
rect 18800 36242 18828 36586
rect 18892 36310 18920 37334
rect 18972 37188 19024 37194
rect 18972 37130 19024 37136
rect 18984 36922 19012 37130
rect 18972 36916 19024 36922
rect 18972 36858 19024 36864
rect 19076 36786 19104 38354
rect 19444 38321 19472 39034
rect 19524 39024 19576 39030
rect 19524 38966 19576 38972
rect 19430 38312 19486 38321
rect 19536 38298 19564 38966
rect 19628 38457 19656 39442
rect 19812 39284 19840 39918
rect 19870 39740 20178 39749
rect 19870 39738 19876 39740
rect 19932 39738 19956 39740
rect 20012 39738 20036 39740
rect 20092 39738 20116 39740
rect 20172 39738 20178 39740
rect 19932 39686 19934 39738
rect 20114 39686 20116 39738
rect 19870 39684 19876 39686
rect 19932 39684 19956 39686
rect 20012 39684 20036 39686
rect 20092 39684 20116 39686
rect 20172 39684 20178 39686
rect 19870 39675 20178 39684
rect 20168 39500 20220 39506
rect 20168 39442 20220 39448
rect 20180 39370 20208 39442
rect 20168 39364 20220 39370
rect 20168 39306 20220 39312
rect 19892 39296 19944 39302
rect 19812 39256 19892 39284
rect 19892 39238 19944 39244
rect 19904 39030 19932 39238
rect 19892 39024 19944 39030
rect 19892 38966 19944 38972
rect 20180 38978 20208 39306
rect 20272 39098 20300 41006
rect 20352 40928 20404 40934
rect 20352 40870 20404 40876
rect 20364 40730 20392 40870
rect 20352 40724 20404 40730
rect 20352 40666 20404 40672
rect 20352 39908 20404 39914
rect 20352 39850 20404 39856
rect 20364 39506 20392 39850
rect 20456 39658 20484 41006
rect 20548 39846 20576 41414
rect 20720 40588 20772 40594
rect 20720 40530 20772 40536
rect 20536 39840 20588 39846
rect 20536 39782 20588 39788
rect 20628 39840 20680 39846
rect 20628 39782 20680 39788
rect 20640 39658 20668 39782
rect 20456 39630 20668 39658
rect 20352 39500 20404 39506
rect 20352 39442 20404 39448
rect 20444 39500 20496 39506
rect 20444 39442 20496 39448
rect 20364 39409 20392 39442
rect 20350 39400 20406 39409
rect 20350 39335 20406 39344
rect 20456 39302 20484 39442
rect 20640 39370 20668 39630
rect 20628 39364 20680 39370
rect 20628 39306 20680 39312
rect 20444 39296 20496 39302
rect 20444 39238 20496 39244
rect 20260 39092 20312 39098
rect 20260 39034 20312 39040
rect 20180 38950 20300 38978
rect 19800 38888 19852 38894
rect 19800 38830 19852 38836
rect 20166 38856 20222 38865
rect 19708 38752 19760 38758
rect 19708 38694 19760 38700
rect 19614 38448 19670 38457
rect 19720 38418 19748 38694
rect 19614 38383 19670 38392
rect 19708 38412 19760 38418
rect 19708 38354 19760 38360
rect 19812 38332 19840 38830
rect 20166 38791 20222 38800
rect 20180 38758 20208 38791
rect 20168 38752 20220 38758
rect 20168 38694 20220 38700
rect 19870 38652 20178 38661
rect 19870 38650 19876 38652
rect 19932 38650 19956 38652
rect 20012 38650 20036 38652
rect 20092 38650 20116 38652
rect 20172 38650 20178 38652
rect 19932 38598 19934 38650
rect 20114 38598 20116 38650
rect 19870 38596 19876 38598
rect 19932 38596 19956 38598
rect 20012 38596 20036 38598
rect 20092 38596 20116 38598
rect 20172 38596 20178 38598
rect 19870 38587 20178 38596
rect 20166 38448 20222 38457
rect 19984 38412 20036 38418
rect 20166 38383 20222 38392
rect 19984 38354 20036 38360
rect 19812 38304 19932 38332
rect 19536 38270 19748 38298
rect 19430 38247 19486 38256
rect 19210 38108 19518 38117
rect 19210 38106 19216 38108
rect 19272 38106 19296 38108
rect 19352 38106 19376 38108
rect 19432 38106 19456 38108
rect 19512 38106 19518 38108
rect 19272 38054 19274 38106
rect 19454 38054 19456 38106
rect 19210 38052 19216 38054
rect 19272 38052 19296 38054
rect 19352 38052 19376 38054
rect 19432 38052 19456 38054
rect 19512 38052 19518 38054
rect 19210 38043 19518 38052
rect 19338 37904 19394 37913
rect 19338 37839 19340 37848
rect 19392 37839 19394 37848
rect 19340 37810 19392 37816
rect 19616 37732 19668 37738
rect 19616 37674 19668 37680
rect 19524 37664 19576 37670
rect 19524 37606 19576 37612
rect 19338 37360 19394 37369
rect 19338 37295 19394 37304
rect 19352 37262 19380 37295
rect 19340 37256 19392 37262
rect 19536 37233 19564 37606
rect 19340 37198 19392 37204
rect 19522 37224 19578 37233
rect 19522 37159 19578 37168
rect 19210 37020 19518 37029
rect 19210 37018 19216 37020
rect 19272 37018 19296 37020
rect 19352 37018 19376 37020
rect 19432 37018 19456 37020
rect 19512 37018 19518 37020
rect 19272 36966 19274 37018
rect 19454 36966 19456 37018
rect 19210 36964 19216 36966
rect 19272 36964 19296 36966
rect 19352 36964 19376 36966
rect 19432 36964 19456 36966
rect 19512 36964 19518 36966
rect 19210 36955 19518 36964
rect 19522 36816 19578 36825
rect 19064 36780 19116 36786
rect 19522 36751 19578 36760
rect 19064 36722 19116 36728
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 18972 36644 19024 36650
rect 18972 36586 19024 36592
rect 18984 36378 19012 36586
rect 18972 36372 19024 36378
rect 18972 36314 19024 36320
rect 18880 36304 18932 36310
rect 18880 36246 18932 36252
rect 18788 36236 18840 36242
rect 18788 36178 18840 36184
rect 18696 36032 18748 36038
rect 18696 35974 18748 35980
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 18708 35222 18736 35974
rect 18788 35488 18840 35494
rect 18788 35430 18840 35436
rect 18696 35216 18748 35222
rect 18696 35158 18748 35164
rect 18800 35154 18828 35430
rect 18788 35148 18840 35154
rect 18788 35090 18840 35096
rect 18892 35018 18920 36246
rect 18984 36038 19012 36314
rect 19062 36272 19118 36281
rect 19062 36207 19118 36216
rect 18972 36032 19024 36038
rect 18972 35974 19024 35980
rect 18880 35012 18932 35018
rect 18880 34954 18932 34960
rect 18984 34898 19012 35974
rect 18892 34870 19012 34898
rect 18524 34462 18644 34490
rect 18510 34096 18566 34105
rect 18510 34031 18512 34040
rect 18564 34031 18566 34040
rect 18512 34002 18564 34008
rect 18524 33522 18552 34002
rect 18616 33969 18644 34462
rect 18892 34082 18920 34870
rect 19076 34746 19104 36207
rect 19260 36174 19288 36654
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19536 36106 19564 36751
rect 19628 36310 19656 37674
rect 19616 36304 19668 36310
rect 19616 36246 19668 36252
rect 19524 36100 19576 36106
rect 19524 36042 19576 36048
rect 19210 35932 19518 35941
rect 19210 35930 19216 35932
rect 19272 35930 19296 35932
rect 19352 35930 19376 35932
rect 19432 35930 19456 35932
rect 19512 35930 19518 35932
rect 19272 35878 19274 35930
rect 19454 35878 19456 35930
rect 19210 35876 19216 35878
rect 19272 35876 19296 35878
rect 19352 35876 19376 35878
rect 19432 35876 19456 35878
rect 19512 35876 19518 35878
rect 19210 35867 19518 35876
rect 19720 35494 19748 38270
rect 19904 38185 19932 38304
rect 19890 38176 19946 38185
rect 19890 38111 19946 38120
rect 19798 38040 19854 38049
rect 19996 38010 20024 38354
rect 20180 38049 20208 38383
rect 20166 38040 20222 38049
rect 19798 37975 19854 37984
rect 19984 38004 20036 38010
rect 19812 37874 19840 37975
rect 20166 37975 20222 37984
rect 19984 37946 20036 37952
rect 19800 37868 19852 37874
rect 19800 37810 19852 37816
rect 19812 35630 19840 37810
rect 20076 37800 20128 37806
rect 20074 37768 20076 37777
rect 20168 37800 20220 37806
rect 20128 37768 20130 37777
rect 20272 37788 20300 38950
rect 20352 38820 20404 38826
rect 20352 38762 20404 38768
rect 20364 38654 20392 38762
rect 20364 38626 20668 38654
rect 20536 38412 20588 38418
rect 20536 38354 20588 38360
rect 20548 38321 20576 38354
rect 20534 38312 20590 38321
rect 20534 38247 20590 38256
rect 20444 38004 20496 38010
rect 20444 37946 20496 37952
rect 20220 37760 20300 37788
rect 20168 37742 20220 37748
rect 20074 37703 20130 37712
rect 19870 37564 20178 37573
rect 19870 37562 19876 37564
rect 19932 37562 19956 37564
rect 20012 37562 20036 37564
rect 20092 37562 20116 37564
rect 20172 37562 20178 37564
rect 19932 37510 19934 37562
rect 20114 37510 20116 37562
rect 19870 37508 19876 37510
rect 19932 37508 19956 37510
rect 20012 37508 20036 37510
rect 20092 37508 20116 37510
rect 20172 37508 20178 37510
rect 19870 37499 20178 37508
rect 20166 37360 20222 37369
rect 20166 37295 20168 37304
rect 20220 37295 20222 37304
rect 20168 37266 20220 37272
rect 20272 36582 20300 37760
rect 20352 37800 20404 37806
rect 20352 37742 20404 37748
rect 20364 37466 20392 37742
rect 20352 37460 20404 37466
rect 20352 37402 20404 37408
rect 20456 37262 20484 37946
rect 20548 37806 20576 38247
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 20640 37670 20668 38626
rect 20732 38010 20760 40530
rect 20824 38486 20852 42094
rect 21008 42022 21036 42094
rect 20996 42016 21048 42022
rect 20996 41958 21048 41964
rect 21008 41546 21036 41958
rect 20996 41540 21048 41546
rect 20996 41482 21048 41488
rect 21100 39982 21128 42162
rect 21272 42016 21324 42022
rect 21272 41958 21324 41964
rect 21284 41682 21312 41958
rect 21272 41676 21324 41682
rect 21272 41618 21324 41624
rect 21364 41676 21416 41682
rect 21364 41618 21416 41624
rect 21376 41274 21404 41618
rect 21364 41268 21416 41274
rect 21364 41210 21416 41216
rect 21468 40662 21496 43590
rect 22020 43178 22048 44134
rect 22928 43852 22980 43858
rect 22928 43794 22980 43800
rect 23388 43852 23440 43858
rect 23440 43812 23520 43840
rect 23388 43794 23440 43800
rect 22376 43648 22428 43654
rect 22376 43590 22428 43596
rect 22388 43246 22416 43590
rect 22376 43240 22428 43246
rect 22376 43182 22428 43188
rect 21640 43172 21692 43178
rect 21640 43114 21692 43120
rect 22008 43172 22060 43178
rect 22008 43114 22060 43120
rect 21652 42158 21680 43114
rect 22284 42560 22336 42566
rect 22284 42502 22336 42508
rect 21640 42152 21692 42158
rect 21640 42094 21692 42100
rect 22008 42152 22060 42158
rect 22008 42094 22060 42100
rect 21916 40928 21968 40934
rect 21916 40870 21968 40876
rect 21456 40656 21508 40662
rect 21456 40598 21508 40604
rect 21928 40594 21956 40870
rect 21916 40588 21968 40594
rect 21916 40530 21968 40536
rect 21456 40384 21508 40390
rect 21456 40326 21508 40332
rect 21468 39982 21496 40326
rect 21088 39976 21140 39982
rect 21088 39918 21140 39924
rect 21456 39976 21508 39982
rect 21456 39918 21508 39924
rect 21100 39302 21128 39918
rect 21088 39296 21140 39302
rect 21088 39238 21140 39244
rect 20812 38480 20864 38486
rect 20812 38422 20864 38428
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 20628 37664 20680 37670
rect 20628 37606 20680 37612
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20352 36644 20404 36650
rect 20352 36586 20404 36592
rect 20260 36576 20312 36582
rect 20260 36518 20312 36524
rect 19870 36476 20178 36485
rect 19870 36474 19876 36476
rect 19932 36474 19956 36476
rect 20012 36474 20036 36476
rect 20092 36474 20116 36476
rect 20172 36474 20178 36476
rect 19932 36422 19934 36474
rect 20114 36422 20116 36474
rect 19870 36420 19876 36422
rect 19932 36420 19956 36422
rect 20012 36420 20036 36422
rect 20092 36420 20116 36422
rect 20172 36420 20178 36422
rect 19870 36411 20178 36420
rect 20272 36242 20300 36518
rect 20260 36236 20312 36242
rect 20260 36178 20312 36184
rect 19800 35624 19852 35630
rect 19800 35566 19852 35572
rect 19708 35488 19760 35494
rect 19708 35430 19760 35436
rect 20260 35488 20312 35494
rect 20260 35430 20312 35436
rect 19870 35388 20178 35397
rect 19870 35386 19876 35388
rect 19932 35386 19956 35388
rect 20012 35386 20036 35388
rect 20092 35386 20116 35388
rect 20172 35386 20178 35388
rect 19932 35334 19934 35386
rect 20114 35334 20116 35386
rect 19870 35332 19876 35334
rect 19932 35332 19956 35334
rect 20012 35332 20036 35334
rect 20092 35332 20116 35334
rect 20172 35332 20178 35334
rect 19870 35323 20178 35332
rect 19800 35284 19852 35290
rect 19800 35226 19852 35232
rect 19708 35012 19760 35018
rect 19708 34954 19760 34960
rect 19210 34844 19518 34853
rect 19210 34842 19216 34844
rect 19272 34842 19296 34844
rect 19352 34842 19376 34844
rect 19432 34842 19456 34844
rect 19512 34842 19518 34844
rect 19272 34790 19274 34842
rect 19454 34790 19456 34842
rect 19210 34788 19216 34790
rect 19272 34788 19296 34790
rect 19352 34788 19376 34790
rect 19432 34788 19456 34790
rect 19512 34788 19518 34790
rect 19210 34779 19518 34788
rect 19064 34740 19116 34746
rect 19064 34682 19116 34688
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 18984 34202 19012 34546
rect 18972 34196 19024 34202
rect 18972 34138 19024 34144
rect 18892 34066 19012 34082
rect 18880 34060 19012 34066
rect 18932 34054 19012 34060
rect 18880 34002 18932 34008
rect 18602 33960 18658 33969
rect 18602 33895 18658 33904
rect 18880 33924 18932 33930
rect 18616 33862 18644 33895
rect 18880 33866 18932 33872
rect 18604 33856 18656 33862
rect 18604 33798 18656 33804
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 18420 32972 18472 32978
rect 18420 32914 18472 32920
rect 18524 31414 18552 33254
rect 18512 31408 18564 31414
rect 18512 31350 18564 31356
rect 18420 31136 18472 31142
rect 18420 31078 18472 31084
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 18144 30932 18196 30938
rect 18196 30892 18276 30920
rect 18144 30874 18196 30880
rect 17880 30190 17908 30874
rect 17592 30184 17644 30190
rect 17592 30126 17644 30132
rect 17868 30184 17920 30190
rect 17868 30126 17920 30132
rect 17604 29850 17632 30126
rect 17592 29844 17644 29850
rect 17592 29786 17644 29792
rect 17880 28626 17908 30126
rect 18144 29776 18196 29782
rect 18144 29718 18196 29724
rect 17960 29708 18012 29714
rect 17960 29650 18012 29656
rect 17972 29306 18000 29650
rect 18052 29504 18104 29510
rect 18156 29492 18184 29718
rect 18104 29464 18184 29492
rect 18052 29446 18104 29452
rect 18156 29306 18184 29464
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 17868 28620 17920 28626
rect 17868 28562 17920 28568
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17972 27470 18000 28358
rect 18144 28212 18196 28218
rect 18144 28154 18196 28160
rect 18156 27674 18184 28154
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17328 26586 17356 27406
rect 17776 27056 17828 27062
rect 17776 26998 17828 27004
rect 17972 27010 18000 27406
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17512 26586 17540 26726
rect 17316 26580 17368 26586
rect 17316 26522 17368 26528
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17144 26438 17540 26466
rect 17132 26036 17184 26042
rect 17132 25978 17184 25984
rect 16948 25424 17000 25430
rect 16948 25366 17000 25372
rect 16212 25356 16264 25362
rect 16132 25316 16212 25344
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 16040 24954 16068 25230
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15856 23662 15884 24278
rect 16132 23798 16160 25316
rect 16212 25298 16264 25304
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24614 16252 25094
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 16224 24274 16252 24550
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 16132 23662 16160 23734
rect 15844 23656 15896 23662
rect 15844 23598 15896 23604
rect 15936 23656 15988 23662
rect 15936 23598 15988 23604
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15304 22066 15424 22094
rect 15396 21554 15424 22066
rect 15948 22030 15976 23598
rect 16132 22778 16160 23598
rect 16224 23322 16252 23598
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 16316 22574 16344 24006
rect 16408 23866 16436 24210
rect 16500 24138 16528 24210
rect 16488 24132 16540 24138
rect 16488 24074 16540 24080
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16500 23746 16528 24074
rect 16408 23718 16528 23746
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16304 22432 16356 22438
rect 16408 22386 16436 23718
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23254 16528 23530
rect 17052 23526 17080 23734
rect 17144 23662 17172 25978
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 16488 23248 16540 23254
rect 16488 23190 16540 23196
rect 16500 22574 16528 23190
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16592 22574 16620 22918
rect 16868 22778 16896 23122
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16356 22380 16436 22386
rect 16304 22374 16436 22380
rect 16224 22098 16252 22374
rect 16316 22358 16436 22374
rect 16316 22166 16344 22358
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 16212 22092 16264 22098
rect 16592 22094 16620 22510
rect 17052 22094 17080 23462
rect 17144 23254 17172 23598
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17316 22094 17368 22098
rect 16592 22066 16804 22094
rect 17052 22092 17368 22094
rect 17052 22066 17316 22092
rect 16212 22034 16264 22040
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15396 21010 15424 21490
rect 15580 21010 15608 21898
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 15672 21010 15700 21354
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16132 21010 16160 21286
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14844 19922 14872 19994
rect 15396 19922 15424 20946
rect 15488 20602 15516 20946
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 16500 19990 16528 21898
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19310 14688 19654
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15212 18834 15240 19178
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15212 18154 15240 18770
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 14844 17746 14872 18022
rect 15304 17882 15332 18022
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15396 17746 15424 19858
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15856 19310 15884 19790
rect 16500 19310 16528 19926
rect 16592 19446 16620 20266
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 15844 19304 15896 19310
rect 16488 19304 16540 19310
rect 15844 19246 15896 19252
rect 16408 19264 16488 19292
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14200 17134 14228 17478
rect 15304 17338 15332 17614
rect 15488 17338 15516 18090
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 12096 16892 12404 16901
rect 12096 16890 12102 16892
rect 12158 16890 12182 16892
rect 12238 16890 12262 16892
rect 12318 16890 12342 16892
rect 12398 16890 12404 16892
rect 12158 16838 12160 16890
rect 12340 16838 12342 16890
rect 12096 16836 12102 16838
rect 12158 16836 12182 16838
rect 12238 16836 12262 16838
rect 12318 16836 12342 16838
rect 12398 16836 12404 16838
rect 12096 16827 12404 16836
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 11436 16348 11744 16357
rect 11436 16346 11442 16348
rect 11498 16346 11522 16348
rect 11578 16346 11602 16348
rect 11658 16346 11682 16348
rect 11738 16346 11744 16348
rect 11498 16294 11500 16346
rect 11680 16294 11682 16346
rect 11436 16292 11442 16294
rect 11498 16292 11522 16294
rect 11578 16292 11602 16294
rect 11658 16292 11682 16294
rect 11738 16292 11744 16294
rect 11436 16283 11744 16292
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 12096 15804 12404 15813
rect 12096 15802 12102 15804
rect 12158 15802 12182 15804
rect 12238 15802 12262 15804
rect 12318 15802 12342 15804
rect 12398 15802 12404 15804
rect 12158 15750 12160 15802
rect 12340 15750 12342 15802
rect 12096 15748 12102 15750
rect 12158 15748 12182 15750
rect 12238 15748 12262 15750
rect 12318 15748 12342 15750
rect 12398 15748 12404 15750
rect 12096 15739 12404 15748
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 11436 15260 11744 15269
rect 11436 15258 11442 15260
rect 11498 15258 11522 15260
rect 11578 15258 11602 15260
rect 11658 15258 11682 15260
rect 11738 15258 11744 15260
rect 11498 15206 11500 15258
rect 11680 15206 11682 15258
rect 11436 15204 11442 15206
rect 11498 15204 11522 15206
rect 11578 15204 11602 15206
rect 11658 15204 11682 15206
rect 11738 15204 11744 15206
rect 11436 15195 11744 15204
rect 13648 14958 13676 17070
rect 15304 16658 15332 17274
rect 15672 16658 15700 19110
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15764 17134 15792 17750
rect 15856 17134 15884 18566
rect 16316 18426 16344 18770
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16040 17134 16068 17682
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15304 15434 15332 16594
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 16046 15424 16390
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 12096 14716 12404 14725
rect 12096 14714 12102 14716
rect 12158 14714 12182 14716
rect 12238 14714 12262 14716
rect 12318 14714 12342 14716
rect 12398 14714 12404 14716
rect 12158 14662 12160 14714
rect 12340 14662 12342 14714
rect 12096 14660 12102 14662
rect 12158 14660 12182 14662
rect 12238 14660 12262 14662
rect 12318 14660 12342 14662
rect 12398 14660 12404 14662
rect 12096 14651 12404 14660
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 11436 14172 11744 14181
rect 11436 14170 11442 14172
rect 11498 14170 11522 14172
rect 11578 14170 11602 14172
rect 11658 14170 11682 14172
rect 11738 14170 11744 14172
rect 11498 14118 11500 14170
rect 11680 14118 11682 14170
rect 11436 14116 11442 14118
rect 11498 14116 11522 14118
rect 11578 14116 11602 14118
rect 11658 14116 11682 14118
rect 11738 14116 11744 14118
rect 11436 14107 11744 14116
rect 13648 13870 13676 14894
rect 15396 14822 15424 15982
rect 15488 15638 15516 16594
rect 15672 16046 15700 16594
rect 16316 16574 16344 18362
rect 16408 18086 16436 19264
rect 16488 19246 16540 19252
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16500 18970 16528 19110
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16592 18834 16620 19110
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16408 17814 16436 18022
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16592 17746 16620 18090
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16224 16546 16344 16574
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16132 16046 16160 16458
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15856 15706 15884 15982
rect 16224 15978 16252 16546
rect 16500 16046 16528 16594
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 13870 14044 14214
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 12096 13628 12404 13637
rect 12096 13626 12102 13628
rect 12158 13626 12182 13628
rect 12238 13626 12262 13628
rect 12318 13626 12342 13628
rect 12398 13626 12404 13628
rect 12158 13574 12160 13626
rect 12340 13574 12342 13626
rect 12096 13572 12102 13574
rect 12158 13572 12182 13574
rect 12238 13572 12262 13574
rect 12318 13572 12342 13574
rect 12398 13572 12404 13574
rect 12096 13563 12404 13572
rect 14200 13394 14228 14758
rect 15396 14482 15424 14758
rect 15488 14550 15516 15574
rect 16224 14958 16252 15914
rect 16408 15586 16436 15982
rect 16500 15706 16528 15982
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16408 15558 16528 15586
rect 16500 15026 16528 15558
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16132 14618 16160 14894
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 11436 13084 11744 13093
rect 11436 13082 11442 13084
rect 11498 13082 11522 13084
rect 11578 13082 11602 13084
rect 11658 13082 11682 13084
rect 11738 13082 11744 13084
rect 11498 13030 11500 13082
rect 11680 13030 11682 13082
rect 11436 13028 11442 13030
rect 11498 13028 11522 13030
rect 11578 13028 11602 13030
rect 11658 13028 11682 13030
rect 11738 13028 11744 13030
rect 11436 13019 11744 13028
rect 14936 12986 14964 13330
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 15028 12782 15056 14214
rect 15304 14074 15332 14282
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15304 13530 15332 14010
rect 15488 13938 15516 14486
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15488 13258 15516 13874
rect 15580 13394 15608 14554
rect 16500 14482 16528 14962
rect 16592 14890 16620 17682
rect 16684 16726 16712 20334
rect 16776 19310 16804 22066
rect 17316 22034 17368 22040
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17144 21486 17172 21830
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17420 19446 17448 22442
rect 17512 22250 17540 26438
rect 17788 25974 17816 26998
rect 17972 26982 18092 27010
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 17868 26240 17920 26246
rect 17868 26182 17920 26188
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 17788 25786 17816 25910
rect 17880 25838 17908 26182
rect 17972 25906 18000 26862
rect 18064 26382 18092 26982
rect 18156 26586 18184 27610
rect 18248 27606 18276 30892
rect 18432 29034 18460 31078
rect 18524 30802 18552 31350
rect 18512 30796 18564 30802
rect 18512 30738 18564 30744
rect 18524 30122 18552 30738
rect 18512 30116 18564 30122
rect 18512 30058 18564 30064
rect 18524 29170 18552 30058
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18420 29028 18472 29034
rect 18420 28970 18472 28976
rect 18432 28558 18460 28970
rect 18524 28694 18552 29106
rect 18512 28688 18564 28694
rect 18512 28630 18564 28636
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18432 28150 18460 28494
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 18236 27600 18288 27606
rect 18236 27542 18288 27548
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 18340 26586 18368 26726
rect 18432 26586 18460 28086
rect 18512 26920 18564 26926
rect 18512 26862 18564 26868
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17696 25758 17816 25786
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17696 24818 17724 25758
rect 17972 25498 18000 25842
rect 18156 25702 18184 26250
rect 18524 26042 18552 26862
rect 18512 26036 18564 26042
rect 18512 25978 18564 25984
rect 18524 25770 18552 25978
rect 18512 25764 18564 25770
rect 18512 25706 18564 25712
rect 18144 25696 18196 25702
rect 18144 25638 18196 25644
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17972 24886 18000 25434
rect 18340 25362 18368 25638
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 18524 24818 18552 25706
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17604 23186 17632 23462
rect 17880 23322 17908 23666
rect 17972 23594 18000 24686
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 18144 23588 18196 23594
rect 18144 23530 18196 23536
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17684 23248 17736 23254
rect 17684 23190 17736 23196
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 17696 22642 17724 23190
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17696 22386 17724 22578
rect 17776 22568 17828 22574
rect 17880 22556 17908 23258
rect 17972 22642 18000 23530
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 18156 22574 18184 23530
rect 17828 22528 17908 22556
rect 17776 22510 17828 22516
rect 17696 22358 17816 22386
rect 17512 22222 17724 22250
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 17604 21146 17632 22034
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17512 20398 17540 20742
rect 17604 20398 17632 20946
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 16776 18952 16804 19246
rect 16856 18964 16908 18970
rect 16776 18924 16856 18952
rect 16856 18906 16908 18912
rect 16960 17882 16988 19246
rect 17236 18154 17264 19246
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17512 17814 17540 18566
rect 17500 17808 17552 17814
rect 17500 17750 17552 17756
rect 17604 17746 17632 20334
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17604 17134 17632 17682
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 17222 16688 17278 16697
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16684 16114 16712 16390
rect 16960 16182 16988 16390
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 17052 16046 17080 16662
rect 17132 16652 17184 16658
rect 17222 16623 17278 16632
rect 17408 16652 17460 16658
rect 17132 16594 17184 16600
rect 17144 16250 17172 16594
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 13802 16436 14214
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13462 16068 13670
rect 16500 13530 16528 14418
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15580 12646 15608 13330
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12782 16160 13126
rect 16592 12782 16620 14826
rect 16684 14618 16712 14894
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16868 14482 16896 15506
rect 16946 15192 17002 15201
rect 16946 15127 16948 15136
rect 17000 15127 17002 15136
rect 16948 15098 17000 15104
rect 17236 15094 17264 16623
rect 17408 16594 17460 16600
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17328 16046 17356 16390
rect 17420 16250 17448 16594
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17592 15904 17644 15910
rect 17696 15892 17724 22222
rect 17788 21690 17816 22358
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17788 18698 17816 19178
rect 17880 18902 17908 22528
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18432 22098 18460 22510
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 17972 21010 18000 21898
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17972 19174 18000 19858
rect 18064 19310 18092 20198
rect 18248 20058 18276 20470
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18340 19990 18368 20198
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17880 18222 17908 18838
rect 18248 18222 18276 19110
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17788 17338 17816 17614
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17880 16454 17908 17750
rect 18064 17746 18092 18022
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 18340 17270 18368 18158
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18236 16720 18288 16726
rect 18236 16662 18288 16668
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17788 16114 17816 16186
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17644 15864 17724 15892
rect 17592 15846 17644 15852
rect 17788 15706 17816 16050
rect 17880 16028 17908 16390
rect 17960 16040 18012 16046
rect 17880 16000 17960 16028
rect 17960 15982 18012 15988
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17788 14618 17816 14894
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 18064 14482 18092 15506
rect 18156 14890 18184 15982
rect 18248 14958 18276 16662
rect 18340 16250 18368 16730
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18432 15978 18460 21286
rect 18616 20942 18644 33798
rect 18800 32552 18828 33798
rect 18892 33658 18920 33866
rect 18880 33652 18932 33658
rect 18880 33594 18932 33600
rect 18984 33454 19012 34054
rect 19076 33590 19104 34682
rect 19616 34536 19668 34542
rect 19616 34478 19668 34484
rect 19524 34468 19576 34474
rect 19524 34410 19576 34416
rect 19156 34060 19208 34066
rect 19156 34002 19208 34008
rect 19168 33969 19196 34002
rect 19154 33960 19210 33969
rect 19154 33895 19210 33904
rect 19536 33862 19564 34410
rect 19628 34066 19656 34478
rect 19720 34066 19748 34954
rect 19812 34406 19840 35226
rect 19892 34944 19944 34950
rect 19892 34886 19944 34892
rect 19904 34542 19932 34886
rect 19892 34536 19944 34542
rect 19892 34478 19944 34484
rect 19800 34400 19852 34406
rect 19800 34342 19852 34348
rect 19812 34066 19840 34342
rect 19870 34300 20178 34309
rect 19870 34298 19876 34300
rect 19932 34298 19956 34300
rect 20012 34298 20036 34300
rect 20092 34298 20116 34300
rect 20172 34298 20178 34300
rect 19932 34246 19934 34298
rect 20114 34246 20116 34298
rect 19870 34244 19876 34246
rect 19932 34244 19956 34246
rect 20012 34244 20036 34246
rect 20092 34244 20116 34246
rect 20172 34244 20178 34246
rect 19870 34235 20178 34244
rect 19616 34060 19668 34066
rect 19616 34002 19668 34008
rect 19708 34060 19760 34066
rect 19708 34002 19760 34008
rect 19800 34060 19852 34066
rect 19800 34002 19852 34008
rect 19524 33856 19576 33862
rect 19524 33798 19576 33804
rect 19616 33856 19668 33862
rect 19668 33816 19748 33844
rect 19616 33798 19668 33804
rect 19210 33756 19518 33765
rect 19210 33754 19216 33756
rect 19272 33754 19296 33756
rect 19352 33754 19376 33756
rect 19432 33754 19456 33756
rect 19512 33754 19518 33756
rect 19272 33702 19274 33754
rect 19454 33702 19456 33754
rect 19210 33700 19216 33702
rect 19272 33700 19296 33702
rect 19352 33700 19376 33702
rect 19432 33700 19456 33702
rect 19512 33700 19518 33702
rect 19210 33691 19518 33700
rect 19064 33584 19116 33590
rect 19064 33526 19116 33532
rect 19616 33516 19668 33522
rect 19616 33458 19668 33464
rect 18972 33448 19024 33454
rect 18972 33390 19024 33396
rect 19064 33380 19116 33386
rect 19064 33322 19116 33328
rect 18972 33312 19024 33318
rect 18972 33254 19024 33260
rect 18880 32564 18932 32570
rect 18800 32524 18880 32552
rect 18880 32506 18932 32512
rect 18892 31890 18920 32506
rect 18984 32434 19012 33254
rect 19076 33114 19104 33322
rect 19064 33108 19116 33114
rect 19064 33050 19116 33056
rect 19210 32668 19518 32677
rect 19210 32666 19216 32668
rect 19272 32666 19296 32668
rect 19352 32666 19376 32668
rect 19432 32666 19456 32668
rect 19512 32666 19518 32668
rect 19272 32614 19274 32666
rect 19454 32614 19456 32666
rect 19210 32612 19216 32614
rect 19272 32612 19296 32614
rect 19352 32612 19376 32614
rect 19432 32612 19456 32614
rect 19512 32612 19518 32614
rect 19210 32603 19518 32612
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 19064 32360 19116 32366
rect 19064 32302 19116 32308
rect 18880 31884 18932 31890
rect 18880 31826 18932 31832
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30938 18736 31214
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 19076 30802 19104 32302
rect 19156 32292 19208 32298
rect 19156 32234 19208 32240
rect 19168 31890 19196 32234
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19444 31822 19472 32438
rect 19524 32224 19576 32230
rect 19524 32166 19576 32172
rect 19536 31890 19564 32166
rect 19524 31884 19576 31890
rect 19524 31826 19576 31832
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19210 31580 19518 31589
rect 19210 31578 19216 31580
rect 19272 31578 19296 31580
rect 19352 31578 19376 31580
rect 19432 31578 19456 31580
rect 19512 31578 19518 31580
rect 19272 31526 19274 31578
rect 19454 31526 19456 31578
rect 19210 31524 19216 31526
rect 19272 31524 19296 31526
rect 19352 31524 19376 31526
rect 19432 31524 19456 31526
rect 19512 31524 19518 31526
rect 19210 31515 19518 31524
rect 19064 30796 19116 30802
rect 19064 30738 19116 30744
rect 19076 30190 19104 30738
rect 19210 30492 19518 30501
rect 19210 30490 19216 30492
rect 19272 30490 19296 30492
rect 19352 30490 19376 30492
rect 19432 30490 19456 30492
rect 19512 30490 19518 30492
rect 19272 30438 19274 30490
rect 19454 30438 19456 30490
rect 19210 30436 19216 30438
rect 19272 30436 19296 30438
rect 19352 30436 19376 30438
rect 19432 30436 19456 30438
rect 19512 30436 19518 30438
rect 19210 30427 19518 30436
rect 19064 30184 19116 30190
rect 19064 30126 19116 30132
rect 18972 30048 19024 30054
rect 18972 29990 19024 29996
rect 18984 29714 19012 29990
rect 18972 29708 19024 29714
rect 18972 29650 19024 29656
rect 19076 28014 19104 30126
rect 19628 29850 19656 33458
rect 19720 32910 19748 33816
rect 19870 33212 20178 33221
rect 19870 33210 19876 33212
rect 19932 33210 19956 33212
rect 20012 33210 20036 33212
rect 20092 33210 20116 33212
rect 20172 33210 20178 33212
rect 19932 33158 19934 33210
rect 20114 33158 20116 33210
rect 19870 33156 19876 33158
rect 19932 33156 19956 33158
rect 20012 33156 20036 33158
rect 20092 33156 20116 33158
rect 20172 33156 20178 33158
rect 19870 33147 20178 33156
rect 19708 32904 19760 32910
rect 19708 32846 19760 32852
rect 19616 29844 19668 29850
rect 19616 29786 19668 29792
rect 19616 29708 19668 29714
rect 19616 29650 19668 29656
rect 19210 29404 19518 29413
rect 19210 29402 19216 29404
rect 19272 29402 19296 29404
rect 19352 29402 19376 29404
rect 19432 29402 19456 29404
rect 19512 29402 19518 29404
rect 19272 29350 19274 29402
rect 19454 29350 19456 29402
rect 19210 29348 19216 29350
rect 19272 29348 19296 29350
rect 19352 29348 19376 29350
rect 19432 29348 19456 29350
rect 19512 29348 19518 29350
rect 19210 29339 19518 29348
rect 19628 29306 19656 29650
rect 19616 29300 19668 29306
rect 19616 29242 19668 29248
rect 19522 29200 19578 29209
rect 19522 29135 19578 29144
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19444 28994 19472 29038
rect 19536 28994 19564 29135
rect 19444 28966 19564 28994
rect 19340 28960 19392 28966
rect 19340 28902 19392 28908
rect 19352 28626 19380 28902
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 19536 28506 19564 28966
rect 19536 28478 19656 28506
rect 19210 28316 19518 28325
rect 19210 28314 19216 28316
rect 19272 28314 19296 28316
rect 19352 28314 19376 28316
rect 19432 28314 19456 28316
rect 19512 28314 19518 28316
rect 19272 28262 19274 28314
rect 19454 28262 19456 28314
rect 19210 28260 19216 28262
rect 19272 28260 19296 28262
rect 19352 28260 19376 28262
rect 19432 28260 19456 28262
rect 19512 28260 19518 28262
rect 19210 28251 19518 28260
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 18696 27872 18748 27878
rect 18696 27814 18748 27820
rect 18708 27538 18736 27814
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 19210 27228 19518 27237
rect 19210 27226 19216 27228
rect 19272 27226 19296 27228
rect 19352 27226 19376 27228
rect 19432 27226 19456 27228
rect 19512 27226 19518 27228
rect 19272 27174 19274 27226
rect 19454 27174 19456 27226
rect 19210 27172 19216 27174
rect 19272 27172 19296 27174
rect 19352 27172 19376 27174
rect 19432 27172 19456 27174
rect 19512 27172 19518 27174
rect 19210 27163 19518 27172
rect 19628 27010 19656 28478
rect 19536 26982 19656 27010
rect 19536 26330 19564 26982
rect 19616 26920 19668 26926
rect 19616 26862 19668 26868
rect 19628 26518 19656 26862
rect 19720 26586 19748 32846
rect 19800 32768 19852 32774
rect 19800 32710 19852 32716
rect 19812 29034 19840 32710
rect 20272 32586 20300 35430
rect 20180 32558 20300 32586
rect 20180 32502 20208 32558
rect 20168 32496 20220 32502
rect 20074 32464 20130 32473
rect 20168 32438 20220 32444
rect 20074 32399 20130 32408
rect 20088 32298 20116 32399
rect 20168 32360 20220 32366
rect 20166 32328 20168 32337
rect 20260 32360 20312 32366
rect 20220 32328 20222 32337
rect 20076 32292 20128 32298
rect 20260 32302 20312 32308
rect 20166 32263 20222 32272
rect 20076 32234 20128 32240
rect 19870 32124 20178 32133
rect 19870 32122 19876 32124
rect 19932 32122 19956 32124
rect 20012 32122 20036 32124
rect 20092 32122 20116 32124
rect 20172 32122 20178 32124
rect 19932 32070 19934 32122
rect 20114 32070 20116 32122
rect 19870 32068 19876 32070
rect 19932 32068 19956 32070
rect 20012 32068 20036 32070
rect 20092 32068 20116 32070
rect 20172 32068 20178 32070
rect 19870 32059 20178 32068
rect 20272 31482 20300 32302
rect 20364 31929 20392 36586
rect 20456 36378 20484 37198
rect 20548 36650 20576 37198
rect 20640 37194 20668 37606
rect 20720 37324 20772 37330
rect 20720 37266 20772 37272
rect 20628 37188 20680 37194
rect 20628 37130 20680 37136
rect 20640 36768 20668 37130
rect 20732 36922 20760 37266
rect 20824 37233 20852 38422
rect 20904 38208 20956 38214
rect 20904 38150 20956 38156
rect 20916 37806 20944 38150
rect 20904 37800 20956 37806
rect 20904 37742 20956 37748
rect 21100 37330 21128 39238
rect 21272 37868 21324 37874
rect 21272 37810 21324 37816
rect 21284 37330 21312 37810
rect 21640 37732 21692 37738
rect 21640 37674 21692 37680
rect 21652 37466 21680 37674
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21640 37460 21692 37466
rect 21640 37402 21692 37408
rect 21836 37369 21864 37606
rect 21822 37360 21878 37369
rect 20904 37324 20956 37330
rect 20904 37266 20956 37272
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 21272 37324 21324 37330
rect 21822 37295 21878 37304
rect 21272 37266 21324 37272
rect 20810 37224 20866 37233
rect 20810 37159 20866 37168
rect 20916 36922 20944 37266
rect 21100 36922 21128 37266
rect 21836 37244 21864 37295
rect 21836 37216 21956 37244
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20904 36916 20956 36922
rect 20904 36858 20956 36864
rect 21088 36916 21140 36922
rect 21088 36858 21140 36864
rect 20640 36740 20760 36768
rect 20536 36644 20588 36650
rect 20536 36586 20588 36592
rect 20628 36644 20680 36650
rect 20628 36586 20680 36592
rect 20444 36372 20496 36378
rect 20444 36314 20496 36320
rect 20350 31920 20406 31929
rect 20350 31855 20406 31864
rect 20350 31648 20406 31657
rect 20350 31583 20406 31592
rect 20260 31476 20312 31482
rect 20260 31418 20312 31424
rect 19870 31036 20178 31045
rect 19870 31034 19876 31036
rect 19932 31034 19956 31036
rect 20012 31034 20036 31036
rect 20092 31034 20116 31036
rect 20172 31034 20178 31036
rect 19932 30982 19934 31034
rect 20114 30982 20116 31034
rect 19870 30980 19876 30982
rect 19932 30980 19956 30982
rect 20012 30980 20036 30982
rect 20092 30980 20116 30982
rect 20172 30980 20178 30982
rect 19870 30971 20178 30980
rect 19870 29948 20178 29957
rect 19870 29946 19876 29948
rect 19932 29946 19956 29948
rect 20012 29946 20036 29948
rect 20092 29946 20116 29948
rect 20172 29946 20178 29948
rect 19932 29894 19934 29946
rect 20114 29894 20116 29946
rect 19870 29892 19876 29894
rect 19932 29892 19956 29894
rect 20012 29892 20036 29894
rect 20092 29892 20116 29894
rect 20172 29892 20178 29894
rect 19870 29883 20178 29892
rect 19892 29776 19944 29782
rect 19892 29718 19944 29724
rect 20260 29776 20312 29782
rect 20260 29718 20312 29724
rect 19904 29238 19932 29718
rect 19892 29232 19944 29238
rect 19892 29174 19944 29180
rect 19800 29028 19852 29034
rect 19800 28970 19852 28976
rect 19870 28860 20178 28869
rect 19870 28858 19876 28860
rect 19932 28858 19956 28860
rect 20012 28858 20036 28860
rect 20092 28858 20116 28860
rect 20172 28858 20178 28860
rect 19932 28806 19934 28858
rect 20114 28806 20116 28858
rect 19870 28804 19876 28806
rect 19932 28804 19956 28806
rect 20012 28804 20036 28806
rect 20092 28804 20116 28806
rect 20172 28804 20178 28806
rect 19870 28795 20178 28804
rect 20272 28626 20300 29718
rect 20364 29510 20392 31583
rect 20456 29714 20484 36314
rect 20444 29708 20496 29714
rect 20444 29650 20496 29656
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20456 29170 20484 29446
rect 20548 29186 20576 36586
rect 20640 36378 20668 36586
rect 20628 36372 20680 36378
rect 20628 36314 20680 36320
rect 20628 36032 20680 36038
rect 20628 35974 20680 35980
rect 20640 35630 20668 35974
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20732 35476 20760 36740
rect 21928 36718 21956 37216
rect 21456 36712 21508 36718
rect 21916 36712 21968 36718
rect 21456 36654 21508 36660
rect 21914 36680 21916 36689
rect 21968 36680 21970 36689
rect 20812 36644 20864 36650
rect 20812 36586 20864 36592
rect 20824 36242 20852 36586
rect 20812 36236 20864 36242
rect 20812 36178 20864 36184
rect 21468 36038 21496 36654
rect 21914 36615 21970 36624
rect 21548 36236 21600 36242
rect 21548 36178 21600 36184
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 20812 35556 20864 35562
rect 20812 35498 20864 35504
rect 20640 35448 20760 35476
rect 20640 31668 20668 35448
rect 20720 35148 20772 35154
rect 20720 35090 20772 35096
rect 20732 34746 20760 35090
rect 20824 35086 20852 35498
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20732 33862 20760 34682
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20824 33674 20852 35022
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21100 34406 21128 34478
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 20732 33646 20852 33674
rect 20732 31754 20760 33646
rect 20812 33312 20864 33318
rect 20812 33254 20864 33260
rect 20824 32314 20852 33254
rect 20904 32496 20956 32502
rect 20902 32464 20904 32473
rect 20956 32464 20958 32473
rect 20902 32399 20958 32408
rect 21100 32366 21128 34342
rect 21272 33856 21324 33862
rect 21272 33798 21324 33804
rect 21284 33386 21312 33798
rect 21272 33380 21324 33386
rect 21272 33322 21324 33328
rect 21468 32978 21496 35974
rect 21560 35834 21588 36178
rect 21824 36032 21876 36038
rect 21824 35974 21876 35980
rect 21548 35828 21600 35834
rect 21548 35770 21600 35776
rect 21836 35698 21864 35974
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21916 35216 21968 35222
rect 22020 35204 22048 42094
rect 22100 41064 22152 41070
rect 22100 41006 22152 41012
rect 22112 39930 22140 41006
rect 22192 40588 22244 40594
rect 22192 40530 22244 40536
rect 22204 40118 22232 40530
rect 22192 40112 22244 40118
rect 22192 40054 22244 40060
rect 22112 39902 22232 39930
rect 22100 39840 22152 39846
rect 22100 39782 22152 39788
rect 22112 39574 22140 39782
rect 22100 39568 22152 39574
rect 22100 39510 22152 39516
rect 22204 39386 22232 39902
rect 22112 39358 22232 39386
rect 22112 36281 22140 39358
rect 22296 38554 22324 42502
rect 22388 42158 22416 43182
rect 22940 42770 22968 43794
rect 23204 43648 23256 43654
rect 23204 43590 23256 43596
rect 23020 43104 23072 43110
rect 23020 43046 23072 43052
rect 23032 42770 23060 43046
rect 22928 42764 22980 42770
rect 22928 42706 22980 42712
rect 23020 42764 23072 42770
rect 23020 42706 23072 42712
rect 22652 42628 22704 42634
rect 22652 42570 22704 42576
rect 22376 42152 22428 42158
rect 22376 42094 22428 42100
rect 22388 41070 22416 42094
rect 22664 41750 22692 42570
rect 23216 42158 23244 43590
rect 23492 43450 23520 43812
rect 24400 43648 24452 43654
rect 24400 43590 24452 43596
rect 23480 43444 23532 43450
rect 23480 43386 23532 43392
rect 23296 43172 23348 43178
rect 23296 43114 23348 43120
rect 23308 42906 23336 43114
rect 23296 42900 23348 42906
rect 23296 42842 23348 42848
rect 23492 42770 23520 43386
rect 23572 43104 23624 43110
rect 23572 43046 23624 43052
rect 24124 43104 24176 43110
rect 24124 43046 24176 43052
rect 23296 42764 23348 42770
rect 23296 42706 23348 42712
rect 23480 42764 23532 42770
rect 23480 42706 23532 42712
rect 23584 42752 23612 43046
rect 23756 42764 23808 42770
rect 23584 42724 23756 42752
rect 23308 42362 23336 42706
rect 23388 42560 23440 42566
rect 23388 42502 23440 42508
rect 23296 42356 23348 42362
rect 23296 42298 23348 42304
rect 23400 42158 23428 42502
rect 22928 42152 22980 42158
rect 22928 42094 22980 42100
rect 23204 42152 23256 42158
rect 23204 42094 23256 42100
rect 23388 42152 23440 42158
rect 23388 42094 23440 42100
rect 22940 42022 22968 42094
rect 22836 42016 22888 42022
rect 22836 41958 22888 41964
rect 22928 42016 22980 42022
rect 22928 41958 22980 41964
rect 22652 41744 22704 41750
rect 22652 41686 22704 41692
rect 22664 41274 22692 41686
rect 22652 41268 22704 41274
rect 22652 41210 22704 41216
rect 22376 41064 22428 41070
rect 22376 41006 22428 41012
rect 22388 39982 22416 41006
rect 22376 39976 22428 39982
rect 22376 39918 22428 39924
rect 22284 38548 22336 38554
rect 22284 38490 22336 38496
rect 22388 38418 22416 39918
rect 22744 39840 22796 39846
rect 22744 39782 22796 39788
rect 22756 39506 22784 39782
rect 22744 39500 22796 39506
rect 22744 39442 22796 39448
rect 22376 38412 22428 38418
rect 22376 38354 22428 38360
rect 22192 38208 22244 38214
rect 22192 38150 22244 38156
rect 22204 37874 22232 38150
rect 22192 37868 22244 37874
rect 22192 37810 22244 37816
rect 22284 37800 22336 37806
rect 22388 37788 22416 38354
rect 22848 38282 22876 41958
rect 22940 39846 22968 41958
rect 23492 41834 23520 42706
rect 23584 42090 23612 42724
rect 23756 42706 23808 42712
rect 23940 42764 23992 42770
rect 23940 42706 23992 42712
rect 24032 42764 24084 42770
rect 24032 42706 24084 42712
rect 23952 42634 23980 42706
rect 23940 42628 23992 42634
rect 23940 42570 23992 42576
rect 23664 42288 23716 42294
rect 23662 42256 23664 42265
rect 23716 42256 23718 42265
rect 23662 42191 23718 42200
rect 24044 42158 24072 42706
rect 24136 42158 24164 43046
rect 24216 42628 24268 42634
rect 24216 42570 24268 42576
rect 24228 42294 24256 42570
rect 24216 42288 24268 42294
rect 24216 42230 24268 42236
rect 24412 42158 24440 43590
rect 24596 43246 24624 44134
rect 25148 43926 25176 44134
rect 25136 43920 25188 43926
rect 25136 43862 25188 43868
rect 24584 43240 24636 43246
rect 24584 43182 24636 43188
rect 24492 42900 24544 42906
rect 24492 42842 24544 42848
rect 24504 42770 24532 42842
rect 25240 42838 25268 44406
rect 25516 44334 25544 44639
rect 26068 44334 26096 44639
rect 26528 44402 26556 44639
rect 26984 44636 27292 44645
rect 26984 44634 26990 44636
rect 27046 44634 27070 44636
rect 27126 44634 27150 44636
rect 27206 44634 27230 44636
rect 27286 44634 27292 44636
rect 27046 44582 27048 44634
rect 27228 44582 27230 44634
rect 26984 44580 26990 44582
rect 27046 44580 27070 44582
rect 27126 44580 27150 44582
rect 27206 44580 27230 44582
rect 27286 44580 27292 44582
rect 26984 44571 27292 44580
rect 27448 44538 27476 44775
rect 27436 44532 27488 44538
rect 27436 44474 27488 44480
rect 26516 44396 26568 44402
rect 26516 44338 26568 44344
rect 28184 44334 28212 44775
rect 28998 44704 29054 44713
rect 28998 44639 29054 44648
rect 29012 44402 29040 44639
rect 29000 44396 29052 44402
rect 29000 44338 29052 44344
rect 25504 44328 25556 44334
rect 25504 44270 25556 44276
rect 26056 44328 26108 44334
rect 26056 44270 26108 44276
rect 28172 44328 28224 44334
rect 28172 44270 28224 44276
rect 29276 44328 29328 44334
rect 29276 44270 29328 44276
rect 27436 44260 27488 44266
rect 27436 44202 27488 44208
rect 25688 44192 25740 44198
rect 25688 44134 25740 44140
rect 26240 44192 26292 44198
rect 26240 44134 26292 44140
rect 27448 44146 27476 44202
rect 28080 44192 28132 44198
rect 25412 43784 25464 43790
rect 25412 43726 25464 43732
rect 25424 43246 25452 43726
rect 25412 43240 25464 43246
rect 25412 43182 25464 43188
rect 25700 43178 25728 44134
rect 26252 43926 26280 44134
rect 27448 44118 27568 44146
rect 28080 44134 28132 44140
rect 29000 44192 29052 44198
rect 29000 44134 29052 44140
rect 26240 43920 26292 43926
rect 26240 43862 26292 43868
rect 27540 43654 27568 44118
rect 27644 44092 27952 44101
rect 27644 44090 27650 44092
rect 27706 44090 27730 44092
rect 27786 44090 27810 44092
rect 27866 44090 27890 44092
rect 27946 44090 27952 44092
rect 27706 44038 27708 44090
rect 27888 44038 27890 44090
rect 27644 44036 27650 44038
rect 27706 44036 27730 44038
rect 27786 44036 27810 44038
rect 27866 44036 27890 44038
rect 27946 44036 27952 44038
rect 27644 44027 27952 44036
rect 27528 43648 27580 43654
rect 27528 43590 27580 43596
rect 26984 43548 27292 43557
rect 26984 43546 26990 43548
rect 27046 43546 27070 43548
rect 27126 43546 27150 43548
rect 27206 43546 27230 43548
rect 27286 43546 27292 43548
rect 27046 43494 27048 43546
rect 27228 43494 27230 43546
rect 26984 43492 26990 43494
rect 27046 43492 27070 43494
rect 27126 43492 27150 43494
rect 27206 43492 27230 43494
rect 27286 43492 27292 43494
rect 26984 43483 27292 43492
rect 27540 43246 27568 43590
rect 27528 43240 27580 43246
rect 27528 43182 27580 43188
rect 25688 43172 25740 43178
rect 25688 43114 25740 43120
rect 25320 43104 25372 43110
rect 25320 43046 25372 43052
rect 26792 43104 26844 43110
rect 26792 43046 26844 43052
rect 25228 42832 25280 42838
rect 25228 42774 25280 42780
rect 24492 42764 24544 42770
rect 24492 42706 24544 42712
rect 24584 42764 24636 42770
rect 24584 42706 24636 42712
rect 24032 42152 24084 42158
rect 24032 42094 24084 42100
rect 24124 42152 24176 42158
rect 24124 42094 24176 42100
rect 24400 42152 24452 42158
rect 24400 42094 24452 42100
rect 23572 42084 23624 42090
rect 23572 42026 23624 42032
rect 23492 41806 23704 41834
rect 24044 41818 24072 42094
rect 23204 41676 23256 41682
rect 23204 41618 23256 41624
rect 23216 40730 23244 41618
rect 23480 41472 23532 41478
rect 23480 41414 23532 41420
rect 23492 41138 23520 41414
rect 23480 41132 23532 41138
rect 23480 41074 23532 41080
rect 23492 41002 23520 41074
rect 23480 40996 23532 41002
rect 23480 40938 23532 40944
rect 23296 40928 23348 40934
rect 23348 40888 23428 40916
rect 23296 40870 23348 40876
rect 23204 40724 23256 40730
rect 23204 40666 23256 40672
rect 23400 40118 23428 40888
rect 23572 40588 23624 40594
rect 23572 40530 23624 40536
rect 23480 40384 23532 40390
rect 23480 40326 23532 40332
rect 23020 40112 23072 40118
rect 23020 40054 23072 40060
rect 23388 40112 23440 40118
rect 23388 40054 23440 40060
rect 22928 39840 22980 39846
rect 22928 39782 22980 39788
rect 22940 38962 22968 39782
rect 22928 38956 22980 38962
rect 22928 38898 22980 38904
rect 22836 38276 22888 38282
rect 22836 38218 22888 38224
rect 22336 37760 22416 37788
rect 22284 37742 22336 37748
rect 22388 37330 22416 37760
rect 22376 37324 22428 37330
rect 22376 37266 22428 37272
rect 22928 37256 22980 37262
rect 22928 37198 22980 37204
rect 22940 36922 22968 37198
rect 22928 36916 22980 36922
rect 22928 36858 22980 36864
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 22098 36272 22154 36281
rect 22098 36207 22154 36216
rect 22376 36236 22428 36242
rect 21968 35176 22048 35204
rect 21916 35158 21968 35164
rect 22020 34542 22048 35176
rect 22112 35170 22140 36207
rect 22376 36178 22428 36184
rect 22560 36236 22612 36242
rect 22560 36178 22612 36184
rect 22282 36136 22338 36145
rect 22282 36071 22284 36080
rect 22336 36071 22338 36080
rect 22284 36042 22336 36048
rect 22192 35556 22244 35562
rect 22192 35498 22244 35504
rect 22204 35290 22232 35498
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 22112 35142 22232 35170
rect 22100 34944 22152 34950
rect 22100 34886 22152 34892
rect 22112 34746 22140 34886
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21744 33658 21772 33934
rect 21732 33652 21784 33658
rect 21732 33594 21784 33600
rect 21732 33448 21784 33454
rect 21732 33390 21784 33396
rect 21456 32972 21508 32978
rect 21456 32914 21508 32920
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 21192 32366 21220 32846
rect 21088 32360 21140 32366
rect 20824 32286 20944 32314
rect 21088 32302 21140 32308
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 20732 31726 20852 31754
rect 20640 31640 20760 31668
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20444 29164 20496 29170
rect 20548 29158 20668 29186
rect 20444 29106 20496 29112
rect 20260 28620 20312 28626
rect 20260 28562 20312 28568
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19996 28082 20024 28358
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 19870 27772 20178 27781
rect 19870 27770 19876 27772
rect 19932 27770 19956 27772
rect 20012 27770 20036 27772
rect 20092 27770 20116 27772
rect 20172 27770 20178 27772
rect 19932 27718 19934 27770
rect 20114 27718 20116 27770
rect 19870 27716 19876 27718
rect 19932 27716 19956 27718
rect 20012 27716 20036 27718
rect 20092 27716 20116 27718
rect 20172 27716 20178 27718
rect 19870 27707 20178 27716
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 20260 27328 20312 27334
rect 20260 27270 20312 27276
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19616 26512 19668 26518
rect 19616 26454 19668 26460
rect 19064 26308 19116 26314
rect 19536 26302 19656 26330
rect 19064 26250 19116 26256
rect 18696 26240 18748 26246
rect 18696 26182 18748 26188
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18708 25430 18736 26182
rect 18696 25424 18748 25430
rect 18696 25366 18748 25372
rect 18788 23656 18840 23662
rect 18786 23624 18788 23633
rect 18840 23624 18842 23633
rect 18786 23559 18842 23568
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18708 22574 18736 23122
rect 18800 22574 18828 23462
rect 18892 23186 18920 26182
rect 19076 25838 19104 26250
rect 19210 26140 19518 26149
rect 19210 26138 19216 26140
rect 19272 26138 19296 26140
rect 19352 26138 19376 26140
rect 19432 26138 19456 26140
rect 19512 26138 19518 26140
rect 19272 26086 19274 26138
rect 19454 26086 19456 26138
rect 19210 26084 19216 26086
rect 19272 26084 19296 26086
rect 19352 26084 19376 26086
rect 19432 26084 19456 26086
rect 19512 26084 19518 26086
rect 19210 26075 19518 26084
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 18984 24818 19012 25706
rect 19076 25158 19104 25774
rect 19064 25152 19116 25158
rect 19064 25094 19116 25100
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 19076 24750 19104 25094
rect 19210 25052 19518 25061
rect 19210 25050 19216 25052
rect 19272 25050 19296 25052
rect 19352 25050 19376 25052
rect 19432 25050 19456 25052
rect 19512 25050 19518 25052
rect 19272 24998 19274 25050
rect 19454 24998 19456 25050
rect 19210 24996 19216 24998
rect 19272 24996 19296 24998
rect 19352 24996 19376 24998
rect 19432 24996 19456 24998
rect 19512 24996 19518 24998
rect 19210 24987 19518 24996
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18800 22234 18828 22510
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18892 22098 18920 22918
rect 18984 22166 19012 24142
rect 19076 23662 19104 24686
rect 19210 23964 19518 23973
rect 19210 23962 19216 23964
rect 19272 23962 19296 23964
rect 19352 23962 19376 23964
rect 19432 23962 19456 23964
rect 19512 23962 19518 23964
rect 19272 23910 19274 23962
rect 19454 23910 19456 23962
rect 19210 23908 19216 23910
rect 19272 23908 19296 23910
rect 19352 23908 19376 23910
rect 19432 23908 19456 23910
rect 19512 23908 19518 23910
rect 19210 23899 19518 23908
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 19246 23624 19302 23633
rect 19246 23559 19248 23568
rect 19300 23559 19302 23568
rect 19248 23530 19300 23536
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19168 23186 19196 23462
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 19628 23050 19656 26302
rect 19812 26246 19840 27270
rect 20272 26926 20300 27270
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 19870 26684 20178 26693
rect 19870 26682 19876 26684
rect 19932 26682 19956 26684
rect 20012 26682 20036 26684
rect 20092 26682 20116 26684
rect 20172 26682 20178 26684
rect 19932 26630 19934 26682
rect 20114 26630 20116 26682
rect 19870 26628 19876 26630
rect 19932 26628 19956 26630
rect 20012 26628 20036 26630
rect 20092 26628 20116 26630
rect 20172 26628 20178 26630
rect 19870 26619 20178 26628
rect 20364 26602 20392 29106
rect 20444 29028 20496 29034
rect 20444 28970 20496 28976
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20456 28082 20484 28970
rect 20548 28762 20576 28970
rect 20536 28756 20588 28762
rect 20536 28698 20588 28704
rect 20536 28552 20588 28558
rect 20536 28494 20588 28500
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20548 27538 20576 28494
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20536 27532 20588 27538
rect 20536 27474 20588 27480
rect 20272 26574 20392 26602
rect 20456 26586 20484 27474
rect 20548 27441 20576 27474
rect 20534 27432 20590 27441
rect 20534 27367 20590 27376
rect 20536 26852 20588 26858
rect 20536 26794 20588 26800
rect 20444 26580 20496 26586
rect 19800 26240 19852 26246
rect 19800 26182 19852 26188
rect 19812 25838 19840 26182
rect 19800 25832 19852 25838
rect 19800 25774 19852 25780
rect 19812 24750 19840 25774
rect 19870 25596 20178 25605
rect 19870 25594 19876 25596
rect 19932 25594 19956 25596
rect 20012 25594 20036 25596
rect 20092 25594 20116 25596
rect 20172 25594 20178 25596
rect 19932 25542 19934 25594
rect 20114 25542 20116 25594
rect 19870 25540 19876 25542
rect 19932 25540 19956 25542
rect 20012 25540 20036 25542
rect 20092 25540 20116 25542
rect 20172 25540 20178 25542
rect 19870 25531 20178 25540
rect 20272 25242 20300 26574
rect 20444 26522 20496 26528
rect 20352 26512 20404 26518
rect 20548 26466 20576 26794
rect 20352 26454 20404 26460
rect 20364 25362 20392 26454
rect 20456 26450 20576 26466
rect 20444 26444 20576 26450
rect 20496 26438 20576 26444
rect 20444 26386 20496 26392
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20272 25214 20576 25242
rect 20260 25152 20312 25158
rect 20260 25094 20312 25100
rect 20272 24818 20300 25094
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19720 23186 19748 23802
rect 19812 23594 19840 24686
rect 20260 24676 20312 24682
rect 20260 24618 20312 24624
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 19870 24508 20178 24517
rect 19870 24506 19876 24508
rect 19932 24506 19956 24508
rect 20012 24506 20036 24508
rect 20092 24506 20116 24508
rect 20172 24506 20178 24508
rect 19932 24454 19934 24506
rect 20114 24454 20116 24506
rect 19870 24452 19876 24454
rect 19932 24452 19956 24454
rect 20012 24452 20036 24454
rect 20092 24452 20116 24454
rect 20172 24452 20178 24454
rect 19870 24443 20178 24452
rect 20272 24449 20300 24618
rect 20258 24440 20314 24449
rect 20364 24410 20392 24618
rect 20258 24375 20314 24384
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20350 23896 20406 23905
rect 20350 23831 20352 23840
rect 20404 23831 20406 23840
rect 20352 23802 20404 23808
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19870 23420 20178 23429
rect 19870 23418 19876 23420
rect 19932 23418 19956 23420
rect 20012 23418 20036 23420
rect 20092 23418 20116 23420
rect 20172 23418 20178 23420
rect 19932 23366 19934 23418
rect 20114 23366 20116 23418
rect 19870 23364 19876 23366
rect 19932 23364 19956 23366
rect 20012 23364 20036 23366
rect 20092 23364 20116 23366
rect 20172 23364 20178 23366
rect 19870 23355 20178 23364
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19616 23044 19668 23050
rect 19616 22986 19668 22992
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19210 22876 19518 22885
rect 19210 22874 19216 22876
rect 19272 22874 19296 22876
rect 19352 22874 19376 22876
rect 19432 22874 19456 22876
rect 19512 22874 19518 22876
rect 19272 22822 19274 22874
rect 19454 22822 19456 22874
rect 19210 22820 19216 22822
rect 19272 22820 19296 22822
rect 19352 22820 19376 22822
rect 19432 22820 19456 22822
rect 19512 22820 19518 22822
rect 19210 22811 19518 22820
rect 19720 22778 19748 22918
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19996 22574 20024 22918
rect 20364 22642 20392 22986
rect 20352 22636 20404 22642
rect 20352 22578 20404 22584
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19870 22332 20178 22341
rect 19870 22330 19876 22332
rect 19932 22330 19956 22332
rect 20012 22330 20036 22332
rect 20092 22330 20116 22332
rect 20172 22330 20178 22332
rect 19932 22278 19934 22330
rect 20114 22278 20116 22330
rect 19870 22276 19876 22278
rect 19932 22276 19956 22278
rect 20012 22276 20036 22278
rect 20092 22276 20116 22278
rect 20172 22276 20178 22278
rect 19870 22267 20178 22276
rect 18972 22160 19024 22166
rect 18972 22102 19024 22108
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18708 21078 18736 21286
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18524 16658 18552 19994
rect 18892 18766 18920 20334
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 18222 18920 18702
rect 18984 18290 19012 22102
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 20168 22092 20220 22098
rect 20364 22094 20392 22578
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20456 22234 20484 22374
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20444 22094 20496 22098
rect 20364 22092 20496 22094
rect 20364 22066 20444 22092
rect 20168 22034 20220 22040
rect 20444 22034 20496 22040
rect 19076 21690 19104 22034
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19210 21788 19518 21797
rect 19210 21786 19216 21788
rect 19272 21786 19296 21788
rect 19352 21786 19376 21788
rect 19432 21786 19456 21788
rect 19512 21786 19518 21788
rect 19272 21734 19274 21786
rect 19454 21734 19456 21786
rect 19210 21732 19216 21734
rect 19272 21732 19296 21734
rect 19352 21732 19376 21734
rect 19432 21732 19456 21734
rect 19512 21732 19518 21734
rect 19210 21723 19518 21732
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 19996 21418 20024 21830
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19800 21344 19852 21350
rect 20088 21332 20116 21626
rect 20180 21468 20208 22034
rect 20444 21956 20496 21962
rect 20444 21898 20496 21904
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20272 21622 20300 21830
rect 20456 21690 20484 21898
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20548 21536 20576 25214
rect 20364 21508 20576 21536
rect 20180 21440 20300 21468
rect 20168 21344 20220 21350
rect 20088 21304 20168 21332
rect 19800 21286 19852 21292
rect 20168 21286 20220 21292
rect 19210 20700 19518 20709
rect 19210 20698 19216 20700
rect 19272 20698 19296 20700
rect 19352 20698 19376 20700
rect 19432 20698 19456 20700
rect 19512 20698 19518 20700
rect 19272 20646 19274 20698
rect 19454 20646 19456 20698
rect 19210 20644 19216 20646
rect 19272 20644 19296 20646
rect 19352 20644 19376 20646
rect 19432 20644 19456 20646
rect 19512 20644 19518 20646
rect 19210 20635 19518 20644
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19168 19922 19196 20198
rect 19260 20058 19288 20334
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19616 19984 19668 19990
rect 19616 19926 19668 19932
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19210 19612 19518 19621
rect 19210 19610 19216 19612
rect 19272 19610 19296 19612
rect 19352 19610 19376 19612
rect 19432 19610 19456 19612
rect 19512 19610 19518 19612
rect 19272 19558 19274 19610
rect 19454 19558 19456 19610
rect 19210 19556 19216 19558
rect 19272 19556 19296 19558
rect 19352 19556 19376 19558
rect 19432 19556 19456 19558
rect 19512 19556 19518 19558
rect 19210 19547 19518 19556
rect 19628 19514 19656 19926
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19720 19378 19748 20198
rect 19812 19718 19840 21286
rect 19870 21244 20178 21253
rect 19870 21242 19876 21244
rect 19932 21242 19956 21244
rect 20012 21242 20036 21244
rect 20092 21242 20116 21244
rect 20172 21242 20178 21244
rect 19932 21190 19934 21242
rect 20114 21190 20116 21242
rect 19870 21188 19876 21190
rect 19932 21188 19956 21190
rect 20012 21188 20036 21190
rect 20092 21188 20116 21190
rect 20172 21188 20178 21190
rect 19870 21179 20178 21188
rect 20272 20466 20300 21440
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 19870 20156 20178 20165
rect 19870 20154 19876 20156
rect 19932 20154 19956 20156
rect 20012 20154 20036 20156
rect 20092 20154 20116 20156
rect 20172 20154 20178 20156
rect 19932 20102 19934 20154
rect 20114 20102 20116 20154
rect 19870 20100 19876 20102
rect 19932 20100 19956 20102
rect 20012 20100 20036 20102
rect 20092 20100 20116 20102
rect 20172 20100 20178 20102
rect 19870 20091 20178 20100
rect 20272 19990 20300 20402
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19812 19310 19840 19654
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19812 18698 19840 19246
rect 19870 19068 20178 19077
rect 19870 19066 19876 19068
rect 19932 19066 19956 19068
rect 20012 19066 20036 19068
rect 20092 19066 20116 19068
rect 20172 19066 20178 19068
rect 19932 19014 19934 19066
rect 20114 19014 20116 19066
rect 19870 19012 19876 19014
rect 19932 19012 19956 19014
rect 20012 19012 20036 19014
rect 20092 19012 20116 19014
rect 20172 19012 20178 19014
rect 19870 19003 20178 19012
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19210 18524 19518 18533
rect 19210 18522 19216 18524
rect 19272 18522 19296 18524
rect 19352 18522 19376 18524
rect 19432 18522 19456 18524
rect 19512 18522 19518 18524
rect 19272 18470 19274 18522
rect 19454 18470 19456 18522
rect 19210 18468 19216 18470
rect 19272 18468 19296 18470
rect 19352 18468 19376 18470
rect 19432 18468 19456 18470
rect 19512 18468 19518 18470
rect 19210 18459 19518 18468
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18892 17134 18920 18158
rect 19628 17882 19656 18566
rect 19812 18154 19840 18634
rect 20272 18290 20300 19926
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18892 16658 18920 17070
rect 19076 17066 19104 17478
rect 19210 17436 19518 17445
rect 19210 17434 19216 17436
rect 19272 17434 19296 17436
rect 19352 17434 19376 17436
rect 19432 17434 19456 17436
rect 19512 17434 19518 17436
rect 19272 17382 19274 17434
rect 19454 17382 19456 17434
rect 19210 17380 19216 17382
rect 19272 17380 19296 17382
rect 19352 17380 19376 17382
rect 19432 17380 19456 17382
rect 19512 17380 19518 17382
rect 19210 17371 19518 17380
rect 19628 17338 19656 17682
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19720 17134 19748 18022
rect 19812 17134 19840 18090
rect 19870 17980 20178 17989
rect 19870 17978 19876 17980
rect 19932 17978 19956 17980
rect 20012 17978 20036 17980
rect 20092 17978 20116 17980
rect 20172 17978 20178 17980
rect 19932 17926 19934 17978
rect 20114 17926 20116 17978
rect 19870 17924 19876 17926
rect 19932 17924 19956 17926
rect 20012 17924 20036 17926
rect 20092 17924 20116 17926
rect 20172 17924 20178 17926
rect 19870 17915 20178 17924
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18156 14550 18184 14826
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 17500 14476 17552 14482
rect 18052 14476 18104 14482
rect 17500 14418 17552 14424
rect 17972 14436 18052 14464
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16684 12986 16712 13806
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16868 12850 16896 14418
rect 17512 14074 17540 14418
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17604 13394 17632 13670
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 12096 12540 12404 12549
rect 12096 12538 12102 12540
rect 12158 12538 12182 12540
rect 12238 12538 12262 12540
rect 12318 12538 12342 12540
rect 12398 12538 12404 12540
rect 12158 12486 12160 12538
rect 12340 12486 12342 12538
rect 12096 12484 12102 12486
rect 12158 12484 12182 12486
rect 12238 12484 12262 12486
rect 12318 12484 12342 12486
rect 12398 12484 12404 12486
rect 12096 12475 12404 12484
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 11436 11996 11744 12005
rect 11436 11994 11442 11996
rect 11498 11994 11522 11996
rect 11578 11994 11602 11996
rect 11658 11994 11682 11996
rect 11738 11994 11744 11996
rect 11498 11942 11500 11994
rect 11680 11942 11682 11994
rect 11436 11940 11442 11942
rect 11498 11940 11522 11942
rect 11578 11940 11602 11942
rect 11658 11940 11682 11942
rect 11738 11940 11744 11942
rect 11436 11931 11744 11940
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 12096 11452 12404 11461
rect 12096 11450 12102 11452
rect 12158 11450 12182 11452
rect 12238 11450 12262 11452
rect 12318 11450 12342 11452
rect 12398 11450 12404 11452
rect 12158 11398 12160 11450
rect 12340 11398 12342 11450
rect 12096 11396 12102 11398
rect 12158 11396 12182 11398
rect 12238 11396 12262 11398
rect 12318 11396 12342 11398
rect 12398 11396 12404 11398
rect 12096 11387 12404 11396
rect 15580 11218 15608 12582
rect 16500 12442 16528 12650
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15672 11354 15700 11562
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15764 11218 15792 12038
rect 16592 11898 16620 12718
rect 16868 12306 16896 12786
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16868 11778 16896 12242
rect 16776 11750 16896 11778
rect 16776 11558 16804 11750
rect 17144 11694 17172 12582
rect 17512 12442 17540 12718
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17972 12306 18000 14436
rect 18052 14418 18104 14424
rect 18248 14414 18276 14894
rect 18340 14822 18368 14894
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18064 12442 18092 12650
rect 18248 12646 18276 14214
rect 18432 13938 18460 14758
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18432 13326 18460 13874
rect 18524 13530 18552 16118
rect 18616 16046 18644 16390
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18432 12782 18460 13262
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 11898 18000 12242
rect 18248 12102 18276 12582
rect 18340 12306 18368 12582
rect 18524 12374 18552 13194
rect 18892 12782 18920 16594
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18984 16046 19012 16458
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 19076 15978 19104 17002
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19628 16697 19656 16934
rect 19870 16892 20178 16901
rect 19870 16890 19876 16892
rect 19932 16890 19956 16892
rect 20012 16890 20036 16892
rect 20092 16890 20116 16892
rect 20172 16890 20178 16892
rect 19932 16838 19934 16890
rect 20114 16838 20116 16890
rect 19870 16836 19876 16838
rect 19932 16836 19956 16838
rect 20012 16836 20036 16838
rect 20092 16836 20116 16838
rect 20172 16836 20178 16838
rect 19870 16827 20178 16836
rect 19614 16688 19670 16697
rect 19614 16623 19670 16632
rect 19708 16652 19760 16658
rect 19628 16590 19656 16623
rect 19708 16594 19760 16600
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19210 16348 19518 16357
rect 19210 16346 19216 16348
rect 19272 16346 19296 16348
rect 19352 16346 19376 16348
rect 19432 16346 19456 16348
rect 19512 16346 19518 16348
rect 19272 16294 19274 16346
rect 19454 16294 19456 16346
rect 19210 16292 19216 16294
rect 19272 16292 19296 16294
rect 19352 16292 19376 16294
rect 19432 16292 19456 16294
rect 19512 16292 19518 16294
rect 19210 16283 19518 16292
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 19352 15348 19380 15982
rect 19536 15502 19564 16186
rect 19628 16046 19656 16526
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19720 15570 19748 16594
rect 20364 16250 20392 21508
rect 20640 21434 20668 29158
rect 20732 27554 20760 31640
rect 20824 31278 20852 31726
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20824 29646 20852 31214
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20916 28762 20944 32286
rect 20996 32292 21048 32298
rect 20996 32234 21048 32240
rect 21008 31414 21036 32234
rect 20996 31408 21048 31414
rect 20996 31350 21048 31356
rect 21008 31278 21036 31350
rect 20996 31272 21048 31278
rect 20996 31214 21048 31220
rect 20904 28756 20956 28762
rect 20904 28698 20956 28704
rect 20902 28520 20958 28529
rect 20902 28455 20958 28464
rect 20916 28014 20944 28455
rect 20904 28008 20956 28014
rect 20904 27950 20956 27956
rect 20732 27526 20944 27554
rect 21100 27538 21128 32302
rect 21284 31346 21312 32302
rect 21364 32020 21416 32026
rect 21364 31962 21416 31968
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 21376 31278 21404 31962
rect 21364 31272 21416 31278
rect 21364 31214 21416 31220
rect 21180 29572 21232 29578
rect 21180 29514 21232 29520
rect 21192 28558 21220 29514
rect 21468 28744 21496 32914
rect 21744 32366 21772 33390
rect 21836 33114 21864 33934
rect 21824 33108 21876 33114
rect 21824 33050 21876 33056
rect 22020 32978 22048 34478
rect 22100 34128 22152 34134
rect 22100 34070 22152 34076
rect 22112 33386 22140 34070
rect 22204 33674 22232 35142
rect 22388 34542 22416 36178
rect 22572 35834 22600 36178
rect 22848 36106 22876 36722
rect 23032 36718 23060 40054
rect 23400 39982 23428 40054
rect 23204 39976 23256 39982
rect 23204 39918 23256 39924
rect 23388 39976 23440 39982
rect 23388 39918 23440 39924
rect 23216 39794 23244 39918
rect 23492 39794 23520 40326
rect 23584 39914 23612 40530
rect 23676 39982 23704 41806
rect 24032 41812 24084 41818
rect 24032 41754 24084 41760
rect 23940 41676 23992 41682
rect 23940 41618 23992 41624
rect 23952 41585 23980 41618
rect 23938 41576 23994 41585
rect 23938 41511 23940 41520
rect 23992 41511 23994 41520
rect 23940 41482 23992 41488
rect 24596 41478 24624 42706
rect 25332 42702 25360 43046
rect 25320 42696 25372 42702
rect 25320 42638 25372 42644
rect 26804 42226 26832 43046
rect 27540 42770 27568 43182
rect 28092 43178 28120 44134
rect 29012 43858 29040 44134
rect 29000 43852 29052 43858
rect 29000 43794 29052 43800
rect 28080 43172 28132 43178
rect 28080 43114 28132 43120
rect 27644 43004 27952 43013
rect 27644 43002 27650 43004
rect 27706 43002 27730 43004
rect 27786 43002 27810 43004
rect 27866 43002 27890 43004
rect 27946 43002 27952 43004
rect 27706 42950 27708 43002
rect 27888 42950 27890 43002
rect 27644 42948 27650 42950
rect 27706 42948 27730 42950
rect 27786 42948 27810 42950
rect 27866 42948 27890 42950
rect 27946 42948 27952 42950
rect 27644 42939 27952 42948
rect 27528 42764 27580 42770
rect 27528 42706 27580 42712
rect 26984 42460 27292 42469
rect 26984 42458 26990 42460
rect 27046 42458 27070 42460
rect 27126 42458 27150 42460
rect 27206 42458 27230 42460
rect 27286 42458 27292 42460
rect 27046 42406 27048 42458
rect 27228 42406 27230 42458
rect 26984 42404 26990 42406
rect 27046 42404 27070 42406
rect 27126 42404 27150 42406
rect 27206 42404 27230 42406
rect 27286 42404 27292 42406
rect 26984 42395 27292 42404
rect 26792 42220 26844 42226
rect 26792 42162 26844 42168
rect 27540 42158 27568 42706
rect 29288 42634 29316 44270
rect 29276 42628 29328 42634
rect 29276 42570 29328 42576
rect 29368 42560 29420 42566
rect 29368 42502 29420 42508
rect 26240 42152 26292 42158
rect 26240 42094 26292 42100
rect 27528 42152 27580 42158
rect 27528 42094 27580 42100
rect 23756 41472 23808 41478
rect 23756 41414 23808 41420
rect 24584 41472 24636 41478
rect 24584 41414 24636 41420
rect 23768 41070 23796 41414
rect 23756 41064 23808 41070
rect 23756 41006 23808 41012
rect 23940 41064 23992 41070
rect 23940 41006 23992 41012
rect 25320 41064 25372 41070
rect 25320 41006 25372 41012
rect 26148 41064 26200 41070
rect 26148 41006 26200 41012
rect 23952 40730 23980 41006
rect 24676 40996 24728 41002
rect 24676 40938 24728 40944
rect 24860 40996 24912 41002
rect 24860 40938 24912 40944
rect 23940 40724 23992 40730
rect 23940 40666 23992 40672
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23572 39908 23624 39914
rect 23572 39850 23624 39856
rect 23216 39766 23520 39794
rect 23216 39574 23244 39766
rect 23584 39658 23612 39850
rect 24216 39840 24268 39846
rect 24216 39782 24268 39788
rect 23492 39642 23612 39658
rect 23492 39636 23624 39642
rect 23492 39630 23572 39636
rect 23204 39568 23256 39574
rect 23204 39510 23256 39516
rect 23020 36712 23072 36718
rect 23072 36672 23152 36700
rect 23020 36654 23072 36660
rect 22836 36100 22888 36106
rect 22836 36042 22888 36048
rect 22560 35828 22612 35834
rect 22560 35770 22612 35776
rect 22572 35290 22600 35770
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 22376 34536 22428 34542
rect 22376 34478 22428 34484
rect 22572 34474 22600 35226
rect 22744 35012 22796 35018
rect 22744 34954 22796 34960
rect 22560 34468 22612 34474
rect 22560 34410 22612 34416
rect 22376 34400 22428 34406
rect 22376 34342 22428 34348
rect 22284 34196 22336 34202
rect 22284 34138 22336 34144
rect 22296 33862 22324 34138
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22204 33646 22324 33674
rect 22100 33380 22152 33386
rect 22100 33322 22152 33328
rect 22008 32972 22060 32978
rect 22008 32914 22060 32920
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21548 32224 21600 32230
rect 21548 32166 21600 32172
rect 21640 32224 21692 32230
rect 21640 32166 21692 32172
rect 21560 31890 21588 32166
rect 21652 31958 21680 32166
rect 21640 31952 21692 31958
rect 21640 31894 21692 31900
rect 21548 31884 21600 31890
rect 21548 31826 21600 31832
rect 21836 31414 21864 32438
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 21824 31408 21876 31414
rect 21824 31350 21876 31356
rect 21836 31210 21864 31350
rect 21916 31340 21968 31346
rect 21916 31282 21968 31288
rect 21928 31210 21956 31282
rect 21824 31204 21876 31210
rect 21376 28716 21496 28744
rect 21652 31164 21824 31192
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 20732 26314 20760 27066
rect 20824 26314 20852 27270
rect 20916 26382 20944 27526
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 21008 26450 21036 26726
rect 20996 26444 21048 26450
rect 20996 26386 21048 26392
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20812 26308 20864 26314
rect 20812 26250 20864 26256
rect 20916 25786 20944 26318
rect 21008 26042 21036 26386
rect 20996 26036 21048 26042
rect 20996 25978 21048 25984
rect 20916 25758 21036 25786
rect 21008 24342 21036 25758
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20732 22506 20760 23122
rect 20824 22574 20852 23802
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21008 22710 21036 23122
rect 20996 22704 21048 22710
rect 20996 22646 21048 22652
rect 21100 22574 21128 27474
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21192 26586 21220 26862
rect 21180 26580 21232 26586
rect 21180 26522 21232 26528
rect 21376 25702 21404 28716
rect 21652 28694 21680 31164
rect 21824 31146 21876 31152
rect 21916 31204 21968 31210
rect 21916 31146 21968 31152
rect 21732 29844 21784 29850
rect 21732 29786 21784 29792
rect 21744 29714 21772 29786
rect 21732 29708 21784 29714
rect 21732 29650 21784 29656
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 21732 28960 21784 28966
rect 21732 28902 21784 28908
rect 21640 28688 21692 28694
rect 21640 28630 21692 28636
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 21468 28150 21496 28562
rect 21652 28490 21680 28630
rect 21640 28484 21692 28490
rect 21640 28426 21692 28432
rect 21744 28422 21772 28902
rect 21732 28416 21784 28422
rect 21732 28358 21784 28364
rect 21456 28144 21508 28150
rect 21456 28086 21508 28092
rect 21732 28076 21784 28082
rect 21732 28018 21784 28024
rect 21640 27600 21692 27606
rect 21560 27560 21640 27588
rect 21456 27328 21508 27334
rect 21456 27270 21508 27276
rect 21468 26926 21496 27270
rect 21456 26920 21508 26926
rect 21456 26862 21508 26868
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21456 25288 21508 25294
rect 21560 25276 21588 27560
rect 21640 27542 21692 27548
rect 21744 27470 21772 28018
rect 21732 27464 21784 27470
rect 21732 27406 21784 27412
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21652 25430 21680 26250
rect 21640 25424 21692 25430
rect 21640 25366 21692 25372
rect 21508 25248 21588 25276
rect 21456 25230 21508 25236
rect 21468 24274 21496 25230
rect 21652 25140 21680 25366
rect 21560 25112 21680 25140
rect 21456 24268 21508 24274
rect 21560 24256 21588 25112
rect 21732 24948 21784 24954
rect 21732 24890 21784 24896
rect 21744 24682 21772 24890
rect 21732 24676 21784 24682
rect 21732 24618 21784 24624
rect 21640 24608 21692 24614
rect 21638 24576 21640 24585
rect 21692 24576 21694 24585
rect 21638 24511 21694 24520
rect 21652 24410 21680 24511
rect 21640 24404 21692 24410
rect 21640 24346 21692 24352
rect 21744 24342 21772 24618
rect 21732 24336 21784 24342
rect 21732 24278 21784 24284
rect 21640 24268 21692 24274
rect 21560 24228 21640 24256
rect 21456 24210 21508 24216
rect 21640 24210 21692 24216
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21376 23186 21404 24074
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21192 22574 21220 22918
rect 21284 22778 21312 23122
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21376 22658 21404 23122
rect 21652 23118 21680 24210
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21468 22778 21496 23054
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21284 22630 21404 22658
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 20732 22098 20760 22442
rect 20720 22092 20772 22098
rect 21284 22094 21312 22630
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21560 22166 21588 22374
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 20720 22034 20772 22040
rect 21192 22066 21312 22094
rect 20456 21406 20668 21434
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20456 16114 20484 21406
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20640 20466 20668 21286
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 19786 20576 20198
rect 20640 19802 20668 20402
rect 20732 20330 20760 22034
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20824 20398 20852 21422
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20720 20324 20772 20330
rect 20720 20266 20772 20272
rect 21088 19848 21140 19854
rect 20536 19780 20588 19786
rect 20640 19774 20760 19802
rect 21088 19790 21140 19796
rect 20536 19722 20588 19728
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19242 20668 19654
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20732 18408 20760 19774
rect 21100 19514 21128 19790
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 20640 18380 20760 18408
rect 20640 18290 20668 18380
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20548 17746 20576 18226
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20732 17338 20760 18226
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20824 17921 20852 18022
rect 20810 17912 20866 17921
rect 20810 17847 20812 17856
rect 20864 17847 20866 17856
rect 20812 17818 20864 17824
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20548 16794 20576 17002
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20916 16046 20944 16390
rect 21192 16114 21220 22066
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21284 21690 21312 21966
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21652 21418 21680 23054
rect 21744 22094 21772 24142
rect 21836 22778 21864 29650
rect 21928 29050 21956 31146
rect 22020 30802 22048 32370
rect 22008 30796 22060 30802
rect 22008 30738 22060 30744
rect 22008 30184 22060 30190
rect 22008 30126 22060 30132
rect 22020 29714 22048 30126
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 21928 29022 22048 29050
rect 21916 28960 21968 28966
rect 21916 28902 21968 28908
rect 21928 28762 21956 28902
rect 21916 28756 21968 28762
rect 21916 28698 21968 28704
rect 21914 28656 21970 28665
rect 21914 28591 21916 28600
rect 21968 28591 21970 28600
rect 21916 28562 21968 28568
rect 21928 24449 21956 28562
rect 22020 28558 22048 29022
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 22020 26790 22048 28494
rect 22112 28218 22140 33322
rect 22192 32360 22244 32366
rect 22192 32302 22244 32308
rect 22204 31482 22232 32302
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22296 31346 22324 33646
rect 22388 33590 22416 34342
rect 22560 34060 22612 34066
rect 22560 34002 22612 34008
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 22388 33454 22416 33526
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22572 33114 22600 34002
rect 22560 33108 22612 33114
rect 22560 33050 22612 33056
rect 22468 32972 22520 32978
rect 22468 32914 22520 32920
rect 22480 32570 22508 32914
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22560 32360 22612 32366
rect 22558 32328 22560 32337
rect 22612 32328 22614 32337
rect 22558 32263 22614 32272
rect 22376 32224 22428 32230
rect 22376 32166 22428 32172
rect 22388 31822 22416 32166
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22388 31278 22416 31622
rect 22572 31278 22600 32263
rect 22652 31476 22704 31482
rect 22652 31418 22704 31424
rect 22376 31272 22428 31278
rect 22376 31214 22428 31220
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22468 31136 22520 31142
rect 22572 31124 22600 31214
rect 22664 31210 22692 31418
rect 22756 31226 22784 34954
rect 22848 34678 22876 36042
rect 22928 35080 22980 35086
rect 22928 35022 22980 35028
rect 22940 34746 22968 35022
rect 22928 34740 22980 34746
rect 22928 34682 22980 34688
rect 22836 34672 22888 34678
rect 22836 34614 22888 34620
rect 22848 32366 22876 34614
rect 23124 33862 23152 36672
rect 23216 36174 23244 39510
rect 23492 39030 23520 39630
rect 23572 39578 23624 39584
rect 24228 39506 24256 39782
rect 23572 39500 23624 39506
rect 23572 39442 23624 39448
rect 24216 39500 24268 39506
rect 24216 39442 24268 39448
rect 24492 39500 24544 39506
rect 24492 39442 24544 39448
rect 23480 39024 23532 39030
rect 23480 38966 23532 38972
rect 23584 38554 23612 39442
rect 23848 39296 23900 39302
rect 23848 39238 23900 39244
rect 23860 38758 23888 39238
rect 24504 39098 24532 39442
rect 24492 39092 24544 39098
rect 24492 39034 24544 39040
rect 23848 38752 23900 38758
rect 23848 38694 23900 38700
rect 23572 38548 23624 38554
rect 23572 38490 23624 38496
rect 23756 38412 23808 38418
rect 23756 38354 23808 38360
rect 23296 38004 23348 38010
rect 23296 37946 23348 37952
rect 23308 37194 23336 37946
rect 23388 37732 23440 37738
rect 23388 37674 23440 37680
rect 23400 37466 23428 37674
rect 23388 37460 23440 37466
rect 23388 37402 23440 37408
rect 23480 37392 23532 37398
rect 23480 37334 23532 37340
rect 23296 37188 23348 37194
rect 23296 37130 23348 37136
rect 23492 37126 23520 37334
rect 23572 37324 23624 37330
rect 23572 37266 23624 37272
rect 23664 37324 23716 37330
rect 23664 37266 23716 37272
rect 23480 37120 23532 37126
rect 23480 37062 23532 37068
rect 23492 36582 23520 37062
rect 23584 36922 23612 37266
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23676 36802 23704 37266
rect 23584 36774 23704 36802
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23492 36378 23520 36518
rect 23480 36372 23532 36378
rect 23480 36314 23532 36320
rect 23480 36236 23532 36242
rect 23584 36224 23612 36774
rect 23664 36712 23716 36718
rect 23664 36654 23716 36660
rect 23676 36242 23704 36654
rect 23768 36378 23796 38354
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23532 36196 23612 36224
rect 23480 36178 23532 36184
rect 23204 36168 23256 36174
rect 23204 36110 23256 36116
rect 23112 33856 23164 33862
rect 23112 33798 23164 33804
rect 23124 32366 23152 33798
rect 22836 32360 22888 32366
rect 22836 32302 22888 32308
rect 23020 32360 23072 32366
rect 23020 32302 23072 32308
rect 23112 32360 23164 32366
rect 23112 32302 23164 32308
rect 23032 32212 23060 32302
rect 23032 32184 23152 32212
rect 23020 31272 23072 31278
rect 22756 31220 23020 31226
rect 22756 31214 23072 31220
rect 22652 31204 22704 31210
rect 22756 31198 23060 31214
rect 22652 31146 22704 31152
rect 22520 31096 22600 31124
rect 22468 31078 22520 31084
rect 22376 30796 22428 30802
rect 22376 30738 22428 30744
rect 22388 29714 22416 30738
rect 22284 29708 22336 29714
rect 22284 29650 22336 29656
rect 22376 29708 22428 29714
rect 22376 29650 22428 29656
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22204 29034 22232 29446
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 22296 28762 22324 29650
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22284 28756 22336 28762
rect 22284 28698 22336 28704
rect 22480 28626 22508 28902
rect 22572 28626 22600 31096
rect 23032 30394 23060 31198
rect 23124 31142 23152 32184
rect 23112 31136 23164 31142
rect 23112 31078 23164 31084
rect 23020 30388 23072 30394
rect 23020 30330 23072 30336
rect 23216 30258 23244 36110
rect 23480 34536 23532 34542
rect 23480 34478 23532 34484
rect 23584 34490 23612 36196
rect 23664 36236 23716 36242
rect 23664 36178 23716 36184
rect 23676 35834 23704 36178
rect 23860 36174 23888 38694
rect 23940 38344 23992 38350
rect 23940 38286 23992 38292
rect 23952 36786 23980 38286
rect 24032 38004 24084 38010
rect 24032 37946 24084 37952
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 24044 36650 24072 37946
rect 24584 37324 24636 37330
rect 24584 37266 24636 37272
rect 24124 36712 24176 36718
rect 24124 36654 24176 36660
rect 24400 36712 24452 36718
rect 24400 36654 24452 36660
rect 24032 36644 24084 36650
rect 24032 36586 24084 36592
rect 24136 36378 24164 36654
rect 24412 36378 24440 36654
rect 24124 36372 24176 36378
rect 24124 36314 24176 36320
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 24596 36242 24624 37266
rect 24124 36236 24176 36242
rect 24124 36178 24176 36184
rect 24584 36236 24636 36242
rect 24584 36178 24636 36184
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 24032 36168 24084 36174
rect 24032 36110 24084 36116
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 23940 35624 23992 35630
rect 23940 35566 23992 35572
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 23492 33454 23520 34478
rect 23584 34462 23704 34490
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 23584 34134 23612 34342
rect 23572 34128 23624 34134
rect 23572 34070 23624 34076
rect 23480 33448 23532 33454
rect 23480 33390 23532 33396
rect 23492 32570 23520 33390
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23492 32366 23520 32506
rect 23480 32360 23532 32366
rect 23480 32302 23532 32308
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23308 31958 23336 32166
rect 23296 31952 23348 31958
rect 23296 31894 23348 31900
rect 23492 31278 23520 32302
rect 23676 31414 23704 34462
rect 23860 33658 23888 35022
rect 23952 34746 23980 35566
rect 24044 35018 24072 36110
rect 24136 35630 24164 36178
rect 24596 35834 24624 36178
rect 24584 35828 24636 35834
rect 24584 35770 24636 35776
rect 24124 35624 24176 35630
rect 24124 35566 24176 35572
rect 24032 35012 24084 35018
rect 24032 34954 24084 34960
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 24124 34468 24176 34474
rect 24124 34410 24176 34416
rect 24492 34468 24544 34474
rect 24492 34410 24544 34416
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 24136 32978 24164 34410
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 24412 33454 24440 33798
rect 24504 33454 24532 34410
rect 24584 34400 24636 34406
rect 24584 34342 24636 34348
rect 24596 34066 24624 34342
rect 24584 34060 24636 34066
rect 24584 34002 24636 34008
rect 24216 33448 24268 33454
rect 24216 33390 24268 33396
rect 24308 33448 24360 33454
rect 24308 33390 24360 33396
rect 24400 33448 24452 33454
rect 24400 33390 24452 33396
rect 24492 33448 24544 33454
rect 24492 33390 24544 33396
rect 24228 33114 24256 33390
rect 24216 33108 24268 33114
rect 24216 33050 24268 33056
rect 24124 32972 24176 32978
rect 24124 32914 24176 32920
rect 24320 32026 24348 33390
rect 24412 32502 24440 33390
rect 24400 32496 24452 32502
rect 24400 32438 24452 32444
rect 24308 32020 24360 32026
rect 24308 31962 24360 31968
rect 24492 31952 24544 31958
rect 24492 31894 24544 31900
rect 24504 31754 24532 31894
rect 24032 31748 24084 31754
rect 24032 31690 24084 31696
rect 24412 31726 24532 31754
rect 24688 31754 24716 40938
rect 24872 40730 24900 40938
rect 25228 40928 25280 40934
rect 25332 40916 25360 41006
rect 25280 40888 25360 40916
rect 25504 40928 25556 40934
rect 25228 40870 25280 40876
rect 25504 40870 25556 40876
rect 24860 40724 24912 40730
rect 24860 40666 24912 40672
rect 24952 40588 25004 40594
rect 24952 40530 25004 40536
rect 24860 39840 24912 39846
rect 24860 39782 24912 39788
rect 24872 39506 24900 39782
rect 24860 39500 24912 39506
rect 24860 39442 24912 39448
rect 24872 39098 24900 39442
rect 24860 39092 24912 39098
rect 24860 39034 24912 39040
rect 24964 37806 24992 40530
rect 25044 40520 25096 40526
rect 25044 40462 25096 40468
rect 25056 39914 25084 40462
rect 25136 40452 25188 40458
rect 25136 40394 25188 40400
rect 25044 39908 25096 39914
rect 25044 39850 25096 39856
rect 25148 39302 25176 40394
rect 25240 39914 25268 40870
rect 25516 40594 25544 40870
rect 25504 40588 25556 40594
rect 25504 40530 25556 40536
rect 26160 40526 26188 41006
rect 26252 40662 26280 42094
rect 28724 42084 28776 42090
rect 28724 42026 28776 42032
rect 26424 42016 26476 42022
rect 26424 41958 26476 41964
rect 27988 42016 28040 42022
rect 27988 41958 28040 41964
rect 26436 41682 26464 41958
rect 27644 41916 27952 41925
rect 27644 41914 27650 41916
rect 27706 41914 27730 41916
rect 27786 41914 27810 41916
rect 27866 41914 27890 41916
rect 27946 41914 27952 41916
rect 27706 41862 27708 41914
rect 27888 41862 27890 41914
rect 27644 41860 27650 41862
rect 27706 41860 27730 41862
rect 27786 41860 27810 41862
rect 27866 41860 27890 41862
rect 27946 41860 27952 41862
rect 27644 41851 27952 41860
rect 28000 41682 28028 41958
rect 26424 41676 26476 41682
rect 26424 41618 26476 41624
rect 26700 41676 26752 41682
rect 26700 41618 26752 41624
rect 27988 41676 28040 41682
rect 27988 41618 28040 41624
rect 28172 41676 28224 41682
rect 28172 41618 28224 41624
rect 26608 41268 26660 41274
rect 26608 41210 26660 41216
rect 26332 41200 26384 41206
rect 26332 41142 26384 41148
rect 26240 40656 26292 40662
rect 26240 40598 26292 40604
rect 26148 40520 26200 40526
rect 26148 40462 26200 40468
rect 26056 40112 26108 40118
rect 26056 40054 26108 40060
rect 25596 39976 25648 39982
rect 25596 39918 25648 39924
rect 25228 39908 25280 39914
rect 25228 39850 25280 39856
rect 25240 39370 25268 39850
rect 25412 39840 25464 39846
rect 25412 39782 25464 39788
rect 25228 39364 25280 39370
rect 25228 39306 25280 39312
rect 25136 39296 25188 39302
rect 25136 39238 25188 39244
rect 25148 38978 25176 39238
rect 25056 38950 25176 38978
rect 25056 38894 25084 38950
rect 25240 38894 25268 39306
rect 25424 39030 25452 39782
rect 25608 39642 25636 39918
rect 25596 39636 25648 39642
rect 25596 39578 25648 39584
rect 25608 39030 25636 39578
rect 26068 39302 26096 40054
rect 26344 39982 26372 41142
rect 26516 40928 26568 40934
rect 26516 40870 26568 40876
rect 26528 40594 26556 40870
rect 26620 40594 26648 41210
rect 26712 40730 26740 41618
rect 27804 41472 27856 41478
rect 27804 41414 27856 41420
rect 26984 41372 27292 41381
rect 26984 41370 26990 41372
rect 27046 41370 27070 41372
rect 27126 41370 27150 41372
rect 27206 41370 27230 41372
rect 27286 41370 27292 41372
rect 27046 41318 27048 41370
rect 27228 41318 27230 41370
rect 26984 41316 26990 41318
rect 27046 41316 27070 41318
rect 27126 41316 27150 41318
rect 27206 41316 27230 41318
rect 27286 41316 27292 41318
rect 26984 41307 27292 41316
rect 27816 41138 27844 41414
rect 28184 41274 28212 41618
rect 28172 41268 28224 41274
rect 28172 41210 28224 41216
rect 26792 41132 26844 41138
rect 26792 41074 26844 41080
rect 27804 41132 27856 41138
rect 27804 41074 27856 41080
rect 26700 40724 26752 40730
rect 26700 40666 26752 40672
rect 26516 40588 26568 40594
rect 26516 40530 26568 40536
rect 26608 40588 26660 40594
rect 26608 40530 26660 40536
rect 26620 40202 26648 40530
rect 26804 40526 26832 41074
rect 28632 41064 28684 41070
rect 28632 41006 28684 41012
rect 27436 40996 27488 41002
rect 27436 40938 27488 40944
rect 27344 40656 27396 40662
rect 27344 40598 27396 40604
rect 26792 40520 26844 40526
rect 26792 40462 26844 40468
rect 26528 40174 26648 40202
rect 26528 39982 26556 40174
rect 26332 39976 26384 39982
rect 26332 39918 26384 39924
rect 26516 39976 26568 39982
rect 26516 39918 26568 39924
rect 26344 39658 26372 39918
rect 26344 39630 26464 39658
rect 26332 39568 26384 39574
rect 26332 39510 26384 39516
rect 26056 39296 26108 39302
rect 26056 39238 26108 39244
rect 26344 39098 26372 39510
rect 26332 39092 26384 39098
rect 26332 39034 26384 39040
rect 25412 39024 25464 39030
rect 25412 38966 25464 38972
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 25870 38992 25926 39001
rect 26436 38978 26464 39630
rect 26528 39438 26556 39918
rect 26804 39574 26832 40462
rect 26984 40284 27292 40293
rect 26984 40282 26990 40284
rect 27046 40282 27070 40284
rect 27126 40282 27150 40284
rect 27206 40282 27230 40284
rect 27286 40282 27292 40284
rect 27046 40230 27048 40282
rect 27228 40230 27230 40282
rect 26984 40228 26990 40230
rect 27046 40228 27070 40230
rect 27126 40228 27150 40230
rect 27206 40228 27230 40230
rect 27286 40228 27292 40230
rect 26984 40219 27292 40228
rect 26884 40180 26936 40186
rect 26884 40122 26936 40128
rect 26792 39568 26844 39574
rect 26792 39510 26844 39516
rect 26896 39438 26924 40122
rect 27356 39506 27384 40598
rect 27448 40526 27476 40938
rect 28540 40928 28592 40934
rect 28540 40870 28592 40876
rect 27644 40828 27952 40837
rect 27644 40826 27650 40828
rect 27706 40826 27730 40828
rect 27786 40826 27810 40828
rect 27866 40826 27890 40828
rect 27946 40826 27952 40828
rect 27706 40774 27708 40826
rect 27888 40774 27890 40826
rect 27644 40772 27650 40774
rect 27706 40772 27730 40774
rect 27786 40772 27810 40774
rect 27866 40772 27890 40774
rect 27946 40772 27952 40774
rect 27644 40763 27952 40772
rect 28552 40594 28580 40870
rect 28356 40588 28408 40594
rect 28540 40588 28592 40594
rect 28356 40530 28408 40536
rect 28460 40548 28540 40576
rect 27436 40520 27488 40526
rect 27436 40462 27488 40468
rect 27448 40186 27476 40462
rect 27436 40180 27488 40186
rect 27436 40122 27488 40128
rect 28368 40050 28396 40530
rect 28460 40118 28488 40548
rect 28540 40530 28592 40536
rect 28644 40390 28672 41006
rect 28632 40384 28684 40390
rect 28632 40326 28684 40332
rect 28540 40180 28592 40186
rect 28540 40122 28592 40128
rect 28448 40112 28500 40118
rect 28448 40054 28500 40060
rect 28356 40044 28408 40050
rect 28356 39986 28408 39992
rect 28552 39982 28580 40122
rect 28540 39976 28592 39982
rect 27724 39902 28028 39930
rect 28540 39918 28592 39924
rect 27724 39846 27752 39902
rect 27712 39840 27764 39846
rect 27712 39782 27764 39788
rect 27644 39740 27952 39749
rect 27644 39738 27650 39740
rect 27706 39738 27730 39740
rect 27786 39738 27810 39740
rect 27866 39738 27890 39740
rect 27946 39738 27952 39740
rect 27706 39686 27708 39738
rect 27888 39686 27890 39738
rect 27644 39684 27650 39686
rect 27706 39684 27730 39686
rect 27786 39684 27810 39686
rect 27866 39684 27890 39686
rect 27946 39684 27952 39686
rect 27644 39675 27952 39684
rect 27344 39500 27396 39506
rect 27344 39442 27396 39448
rect 26516 39432 26568 39438
rect 26884 39432 26936 39438
rect 26516 39374 26568 39380
rect 26620 39380 26884 39386
rect 26620 39374 26936 39380
rect 26620 39358 26924 39374
rect 26620 39098 26648 39358
rect 26792 39296 26844 39302
rect 26792 39238 26844 39244
rect 26884 39296 26936 39302
rect 26884 39238 26936 39244
rect 26608 39092 26660 39098
rect 26608 39034 26660 39040
rect 26436 38950 26556 38978
rect 26620 38962 26648 39034
rect 26804 38962 26832 39238
rect 25870 38927 25872 38936
rect 25924 38927 25926 38936
rect 25872 38898 25924 38904
rect 25044 38888 25096 38894
rect 25044 38830 25096 38836
rect 25228 38888 25280 38894
rect 25228 38830 25280 38836
rect 25136 38480 25188 38486
rect 25136 38422 25188 38428
rect 24952 37800 25004 37806
rect 24952 37742 25004 37748
rect 24964 37398 24992 37742
rect 24952 37392 25004 37398
rect 24952 37334 25004 37340
rect 25148 37330 25176 38422
rect 25884 38010 25912 38898
rect 26424 38888 26476 38894
rect 26424 38830 26476 38836
rect 26436 38758 26464 38830
rect 26424 38752 26476 38758
rect 26424 38694 26476 38700
rect 25872 38004 25924 38010
rect 25872 37946 25924 37952
rect 25136 37324 25188 37330
rect 25136 37266 25188 37272
rect 24952 37120 25004 37126
rect 24952 37062 25004 37068
rect 24768 36644 24820 36650
rect 24768 36586 24820 36592
rect 24780 36242 24808 36586
rect 24964 36242 24992 37062
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 24952 36236 25004 36242
rect 24952 36178 25004 36184
rect 24860 35148 24912 35154
rect 24860 35090 24912 35096
rect 24768 34536 24820 34542
rect 24872 34524 24900 35090
rect 25044 35080 25096 35086
rect 25044 35022 25096 35028
rect 24952 34672 25004 34678
rect 24952 34614 25004 34620
rect 24820 34496 24900 34524
rect 24768 34478 24820 34484
rect 24780 33522 24808 34478
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 24872 33114 24900 34002
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24964 32978 24992 34614
rect 25056 34542 25084 35022
rect 25044 34536 25096 34542
rect 25044 34478 25096 34484
rect 25148 34474 25176 37266
rect 25872 37120 25924 37126
rect 25872 37062 25924 37068
rect 25884 36786 25912 37062
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25228 36644 25280 36650
rect 25228 36586 25280 36592
rect 25240 36310 25268 36586
rect 25780 36576 25832 36582
rect 25780 36518 25832 36524
rect 25792 36310 25820 36518
rect 25228 36304 25280 36310
rect 25228 36246 25280 36252
rect 25780 36304 25832 36310
rect 25780 36246 25832 36252
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 26424 36236 26476 36242
rect 26424 36178 26476 36184
rect 25320 35556 25372 35562
rect 25320 35498 25372 35504
rect 25332 35290 25360 35498
rect 25320 35284 25372 35290
rect 25320 35226 25372 35232
rect 25424 34610 25452 36178
rect 25688 36032 25740 36038
rect 25688 35974 25740 35980
rect 25700 35154 25728 35974
rect 25688 35148 25740 35154
rect 25688 35090 25740 35096
rect 25700 34746 25728 35090
rect 25688 34740 25740 34746
rect 25688 34682 25740 34688
rect 25412 34604 25464 34610
rect 25412 34546 25464 34552
rect 25136 34468 25188 34474
rect 25136 34410 25188 34416
rect 25148 34202 25176 34410
rect 25596 34400 25648 34406
rect 25596 34342 25648 34348
rect 25136 34196 25188 34202
rect 25136 34138 25188 34144
rect 25608 33930 25636 34342
rect 25700 33998 25728 34682
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 26252 34066 26280 34546
rect 26436 34134 26464 36178
rect 26528 35834 26556 38950
rect 26608 38956 26660 38962
rect 26608 38898 26660 38904
rect 26792 38956 26844 38962
rect 26792 38898 26844 38904
rect 26896 38418 26924 39238
rect 26984 39196 27292 39205
rect 26984 39194 26990 39196
rect 27046 39194 27070 39196
rect 27126 39194 27150 39196
rect 27206 39194 27230 39196
rect 27286 39194 27292 39196
rect 27046 39142 27048 39194
rect 27228 39142 27230 39194
rect 26984 39140 26990 39142
rect 27046 39140 27070 39142
rect 27126 39140 27150 39142
rect 27206 39140 27230 39142
rect 27286 39140 27292 39142
rect 26984 39131 27292 39140
rect 27356 39098 27384 39442
rect 27436 39296 27488 39302
rect 27436 39238 27488 39244
rect 27712 39296 27764 39302
rect 27712 39238 27764 39244
rect 27344 39092 27396 39098
rect 27344 39034 27396 39040
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 26884 38412 26936 38418
rect 26884 38354 26936 38360
rect 26988 38298 27016 38694
rect 26896 38270 27016 38298
rect 26896 37330 26924 38270
rect 26984 38108 27292 38117
rect 26984 38106 26990 38108
rect 27046 38106 27070 38108
rect 27126 38106 27150 38108
rect 27206 38106 27230 38108
rect 27286 38106 27292 38108
rect 27046 38054 27048 38106
rect 27228 38054 27230 38106
rect 26984 38052 26990 38054
rect 27046 38052 27070 38054
rect 27126 38052 27150 38054
rect 27206 38052 27230 38054
rect 27286 38052 27292 38054
rect 26984 38043 27292 38052
rect 27344 37392 27396 37398
rect 27344 37334 27396 37340
rect 26884 37324 26936 37330
rect 26884 37266 26936 37272
rect 26700 37256 26752 37262
rect 26700 37198 26752 37204
rect 26608 36644 26660 36650
rect 26608 36586 26660 36592
rect 26620 36242 26648 36586
rect 26712 36378 26740 37198
rect 26884 37188 26936 37194
rect 26884 37130 26936 37136
rect 26792 37120 26844 37126
rect 26792 37062 26844 37068
rect 26700 36372 26752 36378
rect 26700 36314 26752 36320
rect 26712 36242 26740 36314
rect 26804 36242 26832 37062
rect 26896 36242 26924 37130
rect 26984 37020 27292 37029
rect 26984 37018 26990 37020
rect 27046 37018 27070 37020
rect 27126 37018 27150 37020
rect 27206 37018 27230 37020
rect 27286 37018 27292 37020
rect 27046 36966 27048 37018
rect 27228 36966 27230 37018
rect 26984 36964 26990 36966
rect 27046 36964 27070 36966
rect 27126 36964 27150 36966
rect 27206 36964 27230 36966
rect 27286 36964 27292 36966
rect 26984 36955 27292 36964
rect 27356 36922 27384 37334
rect 27448 37194 27476 39238
rect 27724 39001 27752 39238
rect 27710 38992 27766 39001
rect 27710 38927 27766 38936
rect 27644 38652 27952 38661
rect 27644 38650 27650 38652
rect 27706 38650 27730 38652
rect 27786 38650 27810 38652
rect 27866 38650 27890 38652
rect 27946 38650 27952 38652
rect 27706 38598 27708 38650
rect 27888 38598 27890 38650
rect 27644 38596 27650 38598
rect 27706 38596 27730 38598
rect 27786 38596 27810 38598
rect 27866 38596 27890 38598
rect 27946 38596 27952 38598
rect 27644 38587 27952 38596
rect 28000 38486 28028 39902
rect 28356 39908 28408 39914
rect 28356 39850 28408 39856
rect 28368 39506 28396 39850
rect 28356 39500 28408 39506
rect 28356 39442 28408 39448
rect 28552 39438 28580 39918
rect 28644 39846 28672 40326
rect 28736 40050 28764 42026
rect 29000 42016 29052 42022
rect 29000 41958 29052 41964
rect 29276 42016 29328 42022
rect 29276 41958 29328 41964
rect 28816 41812 28868 41818
rect 28816 41754 28868 41760
rect 28724 40044 28776 40050
rect 28724 39986 28776 39992
rect 28632 39840 28684 39846
rect 28632 39782 28684 39788
rect 28736 39438 28764 39986
rect 28828 39914 28856 41754
rect 29012 41154 29040 41958
rect 28920 41138 29040 41154
rect 28908 41132 29040 41138
rect 28960 41126 29040 41132
rect 28908 41074 28960 41080
rect 29288 41070 29316 41958
rect 29380 41682 29408 42502
rect 29552 42152 29604 42158
rect 29552 42094 29604 42100
rect 30748 42152 30800 42158
rect 30748 42094 30800 42100
rect 29564 41818 29592 42094
rect 30760 41818 30788 42094
rect 29552 41812 29604 41818
rect 29552 41754 29604 41760
rect 30748 41812 30800 41818
rect 30748 41754 30800 41760
rect 29368 41676 29420 41682
rect 29368 41618 29420 41624
rect 29460 41676 29512 41682
rect 29460 41618 29512 41624
rect 29472 41274 29500 41618
rect 29460 41268 29512 41274
rect 29460 41210 29512 41216
rect 29552 41132 29604 41138
rect 29552 41074 29604 41080
rect 29276 41064 29328 41070
rect 29276 41006 29328 41012
rect 29460 40928 29512 40934
rect 29460 40870 29512 40876
rect 29472 40594 29500 40870
rect 29460 40588 29512 40594
rect 29460 40530 29512 40536
rect 28908 40112 28960 40118
rect 28908 40054 28960 40060
rect 28816 39908 28868 39914
rect 28816 39850 28868 39856
rect 28080 39432 28132 39438
rect 28080 39374 28132 39380
rect 28540 39432 28592 39438
rect 28540 39374 28592 39380
rect 28724 39432 28776 39438
rect 28724 39374 28776 39380
rect 28092 38826 28120 39374
rect 28080 38820 28132 38826
rect 28080 38762 28132 38768
rect 28552 38554 28580 39374
rect 28724 39296 28776 39302
rect 28724 39238 28776 39244
rect 28540 38548 28592 38554
rect 28540 38490 28592 38496
rect 27988 38480 28040 38486
rect 27988 38422 28040 38428
rect 27644 37564 27952 37573
rect 27644 37562 27650 37564
rect 27706 37562 27730 37564
rect 27786 37562 27810 37564
rect 27866 37562 27890 37564
rect 27946 37562 27952 37564
rect 27706 37510 27708 37562
rect 27888 37510 27890 37562
rect 27644 37508 27650 37510
rect 27706 37508 27730 37510
rect 27786 37508 27810 37510
rect 27866 37508 27890 37510
rect 27946 37508 27952 37510
rect 27644 37499 27952 37508
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 27436 37188 27488 37194
rect 27436 37130 27488 37136
rect 27804 37120 27856 37126
rect 27804 37062 27856 37068
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27816 36786 27844 37062
rect 27804 36780 27856 36786
rect 27804 36722 27856 36728
rect 28080 36576 28132 36582
rect 28080 36518 28132 36524
rect 27644 36476 27952 36485
rect 27644 36474 27650 36476
rect 27706 36474 27730 36476
rect 27786 36474 27810 36476
rect 27866 36474 27890 36476
rect 27946 36474 27952 36476
rect 27706 36422 27708 36474
rect 27888 36422 27890 36474
rect 27644 36420 27650 36422
rect 27706 36420 27730 36422
rect 27786 36420 27810 36422
rect 27866 36420 27890 36422
rect 27946 36420 27952 36422
rect 27644 36411 27952 36420
rect 26608 36236 26660 36242
rect 26608 36178 26660 36184
rect 26700 36236 26752 36242
rect 26700 36178 26752 36184
rect 26792 36236 26844 36242
rect 26792 36178 26844 36184
rect 26884 36236 26936 36242
rect 26884 36178 26936 36184
rect 26792 36032 26844 36038
rect 26792 35974 26844 35980
rect 26516 35828 26568 35834
rect 26516 35770 26568 35776
rect 26700 35624 26752 35630
rect 26700 35566 26752 35572
rect 26712 35222 26740 35566
rect 26700 35216 26752 35222
rect 26700 35158 26752 35164
rect 26712 34746 26740 35158
rect 26700 34740 26752 34746
rect 26700 34682 26752 34688
rect 26804 34218 26832 35974
rect 26984 35932 27292 35941
rect 26984 35930 26990 35932
rect 27046 35930 27070 35932
rect 27126 35930 27150 35932
rect 27206 35930 27230 35932
rect 27286 35930 27292 35932
rect 27046 35878 27048 35930
rect 27228 35878 27230 35930
rect 26984 35876 26990 35878
rect 27046 35876 27070 35878
rect 27126 35876 27150 35878
rect 27206 35876 27230 35878
rect 27286 35876 27292 35878
rect 26984 35867 27292 35876
rect 27160 35828 27212 35834
rect 27160 35770 27212 35776
rect 26884 35692 26936 35698
rect 26884 35634 26936 35640
rect 26896 35222 26924 35634
rect 26884 35216 26936 35222
rect 26884 35158 26936 35164
rect 27172 34950 27200 35770
rect 27988 35692 28040 35698
rect 27988 35634 28040 35640
rect 28000 35494 28028 35634
rect 27252 35488 27304 35494
rect 27252 35430 27304 35436
rect 27988 35488 28040 35494
rect 27988 35430 28040 35436
rect 27264 35290 27292 35430
rect 27644 35388 27952 35397
rect 27644 35386 27650 35388
rect 27706 35386 27730 35388
rect 27786 35386 27810 35388
rect 27866 35386 27890 35388
rect 27946 35386 27952 35388
rect 27706 35334 27708 35386
rect 27888 35334 27890 35386
rect 27644 35332 27650 35334
rect 27706 35332 27730 35334
rect 27786 35332 27810 35334
rect 27866 35332 27890 35334
rect 27946 35332 27952 35334
rect 27644 35323 27952 35332
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 28000 35086 28028 35430
rect 28092 35290 28120 36518
rect 28080 35284 28132 35290
rect 28080 35226 28132 35232
rect 28172 35148 28224 35154
rect 28276 35136 28304 37198
rect 28736 37126 28764 39238
rect 28920 39030 28948 40054
rect 29276 39908 29328 39914
rect 29276 39850 29328 39856
rect 29184 39364 29236 39370
rect 29184 39306 29236 39312
rect 28908 39024 28960 39030
rect 28908 38966 28960 38972
rect 29196 38826 29224 39306
rect 29288 38894 29316 39850
rect 29472 39574 29500 40530
rect 29564 40526 29592 41074
rect 31116 41064 31168 41070
rect 31116 41006 31168 41012
rect 30748 40996 30800 41002
rect 30748 40938 30800 40944
rect 30760 40730 30788 40938
rect 30932 40928 30984 40934
rect 30932 40870 30984 40876
rect 30748 40724 30800 40730
rect 30748 40666 30800 40672
rect 30944 40594 30972 40870
rect 31128 40730 31156 41006
rect 31116 40724 31168 40730
rect 31116 40666 31168 40672
rect 30932 40588 30984 40594
rect 30932 40530 30984 40536
rect 31024 40588 31076 40594
rect 31024 40530 31076 40536
rect 29552 40520 29604 40526
rect 29552 40462 29604 40468
rect 29460 39568 29512 39574
rect 29460 39510 29512 39516
rect 29472 39098 29500 39510
rect 29564 39438 29592 40462
rect 30380 40384 30432 40390
rect 30380 40326 30432 40332
rect 29920 39976 29972 39982
rect 29920 39918 29972 39924
rect 29828 39840 29880 39846
rect 29828 39782 29880 39788
rect 29840 39506 29868 39782
rect 29828 39500 29880 39506
rect 29828 39442 29880 39448
rect 29552 39432 29604 39438
rect 29552 39374 29604 39380
rect 29460 39092 29512 39098
rect 29460 39034 29512 39040
rect 29276 38888 29328 38894
rect 29276 38830 29328 38836
rect 29184 38820 29236 38826
rect 29184 38762 29236 38768
rect 28816 38752 28868 38758
rect 28816 38694 28868 38700
rect 28828 37262 28856 38694
rect 29092 38208 29144 38214
rect 29092 38150 29144 38156
rect 29104 37874 29132 38150
rect 29092 37868 29144 37874
rect 29092 37810 29144 37816
rect 29196 37754 29224 38762
rect 29288 38418 29316 38830
rect 29276 38412 29328 38418
rect 29276 38354 29328 38360
rect 29104 37726 29224 37754
rect 29000 37460 29052 37466
rect 29000 37402 29052 37408
rect 29012 37330 29040 37402
rect 29104 37330 29132 37726
rect 29000 37324 29052 37330
rect 29000 37266 29052 37272
rect 29092 37324 29144 37330
rect 29092 37266 29144 37272
rect 28816 37256 28868 37262
rect 28816 37198 28868 37204
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28448 35828 28500 35834
rect 28448 35770 28500 35776
rect 28460 35494 28488 35770
rect 28448 35488 28500 35494
rect 28448 35430 28500 35436
rect 28224 35108 28304 35136
rect 28356 35148 28408 35154
rect 28172 35090 28224 35096
rect 28356 35090 28408 35096
rect 27988 35080 28040 35086
rect 27988 35022 28040 35028
rect 27160 34944 27212 34950
rect 27160 34886 27212 34892
rect 27344 34944 27396 34950
rect 27344 34886 27396 34892
rect 27988 34944 28040 34950
rect 27988 34886 28040 34892
rect 26984 34844 27292 34853
rect 26984 34842 26990 34844
rect 27046 34842 27070 34844
rect 27126 34842 27150 34844
rect 27206 34842 27230 34844
rect 27286 34842 27292 34844
rect 27046 34790 27048 34842
rect 27228 34790 27230 34842
rect 26984 34788 26990 34790
rect 27046 34788 27070 34790
rect 27126 34788 27150 34790
rect 27206 34788 27230 34790
rect 27286 34788 27292 34790
rect 26984 34779 27292 34788
rect 27356 34474 27384 34886
rect 27344 34468 27396 34474
rect 27344 34410 27396 34416
rect 27644 34300 27952 34309
rect 27644 34298 27650 34300
rect 27706 34298 27730 34300
rect 27786 34298 27810 34300
rect 27866 34298 27890 34300
rect 27946 34298 27952 34300
rect 27706 34246 27708 34298
rect 27888 34246 27890 34298
rect 27644 34244 27650 34246
rect 27706 34244 27730 34246
rect 27786 34244 27810 34246
rect 27866 34244 27890 34246
rect 27946 34244 27952 34246
rect 27644 34235 27952 34244
rect 26804 34190 26924 34218
rect 26424 34128 26476 34134
rect 26424 34070 26476 34076
rect 26792 34128 26844 34134
rect 26792 34070 26844 34076
rect 26240 34060 26292 34066
rect 26240 34002 26292 34008
rect 25688 33992 25740 33998
rect 25688 33934 25740 33940
rect 25596 33924 25648 33930
rect 25596 33866 25648 33872
rect 25136 33516 25188 33522
rect 25136 33458 25188 33464
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 25148 32910 25176 33458
rect 25700 32978 25728 33934
rect 26148 33856 26200 33862
rect 26148 33798 26200 33804
rect 26160 33658 26188 33798
rect 26148 33652 26200 33658
rect 26148 33594 26200 33600
rect 26056 33448 26108 33454
rect 26252 33402 26280 34002
rect 26516 33924 26568 33930
rect 26516 33866 26568 33872
rect 26332 33856 26384 33862
rect 26332 33798 26384 33804
rect 26108 33396 26280 33402
rect 26056 33390 26280 33396
rect 26068 33374 26280 33390
rect 25688 32972 25740 32978
rect 25688 32914 25740 32920
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 25136 32904 25188 32910
rect 25136 32846 25188 32852
rect 24688 31726 24808 31754
rect 24044 31482 24072 31690
rect 24032 31476 24084 31482
rect 24032 31418 24084 31424
rect 23664 31408 23716 31414
rect 23664 31350 23716 31356
rect 24124 31408 24176 31414
rect 24124 31350 24176 31356
rect 23480 31272 23532 31278
rect 23480 31214 23532 31220
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23492 29782 23520 31214
rect 23664 31204 23716 31210
rect 23664 31146 23716 31152
rect 23676 30938 23704 31146
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23940 30796 23992 30802
rect 23940 30738 23992 30744
rect 23952 30394 23980 30738
rect 24136 30394 24164 31350
rect 24216 31136 24268 31142
rect 24216 31078 24268 31084
rect 24228 30802 24256 31078
rect 24216 30796 24268 30802
rect 24216 30738 24268 30744
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 24124 30388 24176 30394
rect 24124 30330 24176 30336
rect 23570 30288 23626 30297
rect 23570 30223 23626 30232
rect 23848 30252 23900 30258
rect 23480 29776 23532 29782
rect 23480 29718 23532 29724
rect 23584 29714 23612 30223
rect 23848 30194 23900 30200
rect 23572 29708 23624 29714
rect 23572 29650 23624 29656
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 22652 29504 22704 29510
rect 22652 29446 22704 29452
rect 22664 29102 22692 29446
rect 22652 29096 22704 29102
rect 22652 29038 22704 29044
rect 23124 28626 23152 29514
rect 23204 29504 23256 29510
rect 23204 29446 23256 29452
rect 23216 29034 23244 29446
rect 23664 29164 23716 29170
rect 23664 29106 23716 29112
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23216 28694 23244 28970
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23204 28688 23256 28694
rect 23204 28630 23256 28636
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 22112 25242 22140 28154
rect 22572 28150 22600 28562
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22284 28008 22336 28014
rect 22284 27950 22336 27956
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22204 26518 22232 27814
rect 22296 26586 22324 27950
rect 22388 27334 22416 28086
rect 22836 27940 22888 27946
rect 22836 27882 22888 27888
rect 22744 27464 22796 27470
rect 22848 27452 22876 27882
rect 23308 27674 23336 28902
rect 23400 28694 23428 29038
rect 23388 28688 23440 28694
rect 23388 28630 23440 28636
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23676 27606 23704 29106
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 22796 27424 22876 27452
rect 22744 27406 22796 27412
rect 22468 27396 22520 27402
rect 22468 27338 22520 27344
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22376 27328 22428 27334
rect 22376 27270 22428 27276
rect 22388 26858 22416 27270
rect 22480 26994 22508 27338
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22376 26852 22428 26858
rect 22376 26794 22428 26800
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22192 26512 22244 26518
rect 22192 26454 22244 26460
rect 22296 25362 22324 26522
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22112 25214 22232 25242
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22008 24744 22060 24750
rect 22112 24732 22140 25094
rect 22060 24704 22140 24732
rect 22008 24686 22060 24692
rect 21914 24440 21970 24449
rect 21914 24375 21970 24384
rect 22204 23322 22232 25214
rect 22376 25152 22428 25158
rect 22376 25094 22428 25100
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22296 24410 22324 24618
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22388 24342 22416 25094
rect 22480 24698 22508 26930
rect 22572 26790 22600 27338
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 26926 22784 27270
rect 22744 26920 22796 26926
rect 22744 26862 22796 26868
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22664 26518 22692 26726
rect 22652 26512 22704 26518
rect 22652 26454 22704 26460
rect 22480 24670 22600 24698
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22480 24449 22508 24550
rect 22466 24440 22522 24449
rect 22466 24375 22522 24384
rect 22376 24336 22428 24342
rect 22376 24278 22428 24284
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 22020 22574 22048 23190
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 22112 22710 22140 23122
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22204 22574 22232 22646
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 21744 22066 21864 22094
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 21640 21412 21692 21418
rect 21640 21354 21692 21360
rect 21652 20398 21680 21354
rect 21744 21146 21772 21422
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21652 19922 21680 20334
rect 21732 20324 21784 20330
rect 21732 20266 21784 20272
rect 21744 19922 21772 20266
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21284 17678 21312 18906
rect 21468 18816 21496 19246
rect 21560 18970 21588 19246
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21548 18828 21600 18834
rect 21468 18788 21548 18816
rect 21548 18770 21600 18776
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 16658 21312 17478
rect 21376 16658 21404 17682
rect 21560 17134 21588 18770
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21652 18222 21680 18634
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21652 17814 21680 18158
rect 21744 18154 21772 19858
rect 21836 18290 21864 22066
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22112 21010 22140 21626
rect 22296 21486 22324 22986
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 22020 19990 22048 20334
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22112 20058 22140 20198
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 22020 19514 22048 19926
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22112 18970 22140 19178
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22204 18834 22232 20198
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22296 18902 22324 19790
rect 22388 19174 22416 21286
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21732 18148 21784 18154
rect 21732 18090 21784 18096
rect 21640 17808 21692 17814
rect 21640 17750 21692 17756
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21560 16046 21588 17070
rect 21652 16726 21680 17750
rect 21744 17746 21772 18090
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21744 16726 21772 17682
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 19870 15804 20178 15813
rect 19870 15802 19876 15804
rect 19932 15802 19956 15804
rect 20012 15802 20036 15804
rect 20092 15802 20116 15804
rect 20172 15802 20178 15804
rect 19932 15750 19934 15802
rect 20114 15750 20116 15802
rect 19870 15748 19876 15750
rect 19932 15748 19956 15750
rect 20012 15748 20036 15750
rect 20092 15748 20116 15750
rect 20172 15748 20178 15750
rect 19870 15739 20178 15748
rect 21100 15638 21128 15846
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 21284 15570 21312 15846
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19076 15320 19380 15348
rect 18972 14952 19024 14958
rect 19076 14940 19104 15320
rect 19210 15260 19518 15269
rect 19210 15258 19216 15260
rect 19272 15258 19296 15260
rect 19352 15258 19376 15260
rect 19432 15258 19456 15260
rect 19512 15258 19518 15260
rect 19272 15206 19274 15258
rect 19454 15206 19456 15258
rect 19210 15204 19216 15206
rect 19272 15204 19296 15206
rect 19352 15204 19376 15206
rect 19432 15204 19456 15206
rect 19512 15204 19518 15206
rect 19210 15195 19518 15204
rect 19628 15026 19656 15370
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19720 14958 19748 15302
rect 20916 15162 20944 15438
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 19024 14912 19104 14940
rect 19708 14952 19760 14958
rect 18972 14894 19024 14900
rect 19708 14894 19760 14900
rect 20916 14890 20944 15098
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18984 14006 19012 14758
rect 19870 14716 20178 14725
rect 19870 14714 19876 14716
rect 19932 14714 19956 14716
rect 20012 14714 20036 14716
rect 20092 14714 20116 14716
rect 20172 14714 20178 14716
rect 19932 14662 19934 14714
rect 20114 14662 20116 14714
rect 19870 14660 19876 14662
rect 19932 14660 19956 14662
rect 20012 14660 20036 14662
rect 20092 14660 20116 14662
rect 20172 14660 20178 14662
rect 19870 14651 20178 14660
rect 21560 14482 21588 15982
rect 21836 14958 21864 17478
rect 21928 17338 21956 17818
rect 22020 17746 22048 18226
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22112 17377 22140 17614
rect 22098 17368 22154 17377
rect 21916 17332 21968 17338
rect 22098 17303 22154 17312
rect 21916 17274 21968 17280
rect 22480 16658 22508 24375
rect 22572 23186 22600 24670
rect 22560 23180 22612 23186
rect 22560 23122 22612 23128
rect 22756 22710 22784 26726
rect 22848 26518 22876 27424
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23032 26926 23060 27270
rect 23308 26926 23336 27474
rect 23480 27464 23532 27470
rect 23676 27441 23704 27542
rect 23480 27406 23532 27412
rect 23662 27432 23718 27441
rect 23020 26920 23072 26926
rect 23020 26862 23072 26868
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23400 26772 23428 26862
rect 23308 26744 23428 26772
rect 23308 26586 23336 26744
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 23296 26580 23348 26586
rect 23296 26522 23348 26528
rect 22836 26512 22888 26518
rect 22836 26454 22888 26460
rect 22848 25362 22876 26454
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22848 24954 22876 25298
rect 23020 25288 23072 25294
rect 23020 25230 23072 25236
rect 22928 25220 22980 25226
rect 22928 25162 22980 25168
rect 22940 24954 22968 25162
rect 22836 24948 22888 24954
rect 22836 24890 22888 24896
rect 22928 24948 22980 24954
rect 22928 24890 22980 24896
rect 23032 24614 23060 25230
rect 23124 24750 23152 26522
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23204 25696 23256 25702
rect 23204 25638 23256 25644
rect 23216 25226 23244 25638
rect 23400 25430 23428 26386
rect 23492 26246 23520 27406
rect 23662 27367 23718 27376
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23584 26382 23612 26726
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23572 26240 23624 26246
rect 23572 26182 23624 26188
rect 23388 25424 23440 25430
rect 23388 25366 23440 25372
rect 23584 25362 23612 26182
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 23204 25220 23256 25226
rect 23204 25162 23256 25168
rect 23112 24744 23164 24750
rect 23216 24732 23244 25162
rect 23492 24970 23520 25298
rect 23584 25158 23612 25298
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23492 24942 23612 24970
rect 23216 24704 23336 24732
rect 23112 24686 23164 24692
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 23124 23254 23152 24686
rect 23112 23248 23164 23254
rect 23032 23208 23112 23236
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 23032 22574 23060 23208
rect 23112 23190 23164 23196
rect 23112 22976 23164 22982
rect 23112 22918 23164 22924
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22848 21894 22876 22034
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22756 21146 22784 21830
rect 23032 21690 23060 22510
rect 23124 22098 23152 22918
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23216 22273 23244 22374
rect 23202 22264 23258 22273
rect 23202 22199 23258 22208
rect 23204 22160 23256 22166
rect 23204 22102 23256 22108
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 23216 21690 23244 22102
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23204 21480 23256 21486
rect 23202 21448 23204 21457
rect 23256 21448 23258 21457
rect 23202 21383 23258 21392
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 23308 20466 23336 24704
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23492 24342 23520 24550
rect 23584 24410 23612 24942
rect 23676 24682 23704 27367
rect 23768 26246 23796 27950
rect 23756 26240 23808 26246
rect 23756 26182 23808 26188
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23768 24750 23796 25094
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23664 24676 23716 24682
rect 23664 24618 23716 24624
rect 23572 24404 23624 24410
rect 23572 24346 23624 24352
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 23676 24070 23704 24618
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23768 24274 23796 24550
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22572 20262 22600 20334
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 22572 19514 22600 20198
rect 23400 19990 23428 23258
rect 23676 22438 23704 24006
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23570 22264 23626 22273
rect 23480 22228 23532 22234
rect 23570 22199 23626 22208
rect 23480 22170 23532 22176
rect 23492 20398 23520 22170
rect 23584 21554 23612 22199
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23584 21350 23612 21490
rect 23754 21448 23810 21457
rect 23754 21383 23810 21392
rect 23768 21350 23796 21383
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23388 19984 23440 19990
rect 23860 19938 23888 30194
rect 23940 30184 23992 30190
rect 23940 30126 23992 30132
rect 23952 28014 23980 30126
rect 24136 30104 24164 30330
rect 24216 30116 24268 30122
rect 24136 30076 24216 30104
rect 24216 30058 24268 30064
rect 24308 30116 24360 30122
rect 24308 30058 24360 30064
rect 24032 29096 24084 29102
rect 24032 29038 24084 29044
rect 24044 28218 24072 29038
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 24228 28014 24256 30058
rect 24320 29850 24348 30058
rect 24308 29844 24360 29850
rect 24308 29786 24360 29792
rect 23940 28008 23992 28014
rect 23940 27950 23992 27956
rect 24216 28008 24268 28014
rect 24216 27950 24268 27956
rect 24320 27946 24348 29786
rect 24308 27940 24360 27946
rect 24308 27882 24360 27888
rect 23940 27872 23992 27878
rect 23940 27814 23992 27820
rect 23952 21146 23980 27814
rect 24412 27538 24440 31726
rect 24584 28620 24636 28626
rect 24584 28562 24636 28568
rect 24490 28112 24546 28121
rect 24490 28047 24546 28056
rect 24504 28014 24532 28047
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 24032 27532 24084 27538
rect 24032 27474 24084 27480
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24492 27532 24544 27538
rect 24492 27474 24544 27480
rect 24044 26586 24072 27474
rect 24216 27464 24268 27470
rect 24216 27406 24268 27412
rect 24124 27328 24176 27334
rect 24124 27270 24176 27276
rect 24136 26926 24164 27270
rect 24228 27130 24256 27406
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24412 26926 24440 27474
rect 24124 26920 24176 26926
rect 24124 26862 24176 26868
rect 24400 26920 24452 26926
rect 24400 26862 24452 26868
rect 24032 26580 24084 26586
rect 24032 26522 24084 26528
rect 24504 26518 24532 27474
rect 24596 27334 24624 28562
rect 24676 27940 24728 27946
rect 24676 27882 24728 27888
rect 24688 27402 24716 27882
rect 24676 27396 24728 27402
rect 24676 27338 24728 27344
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24492 26512 24544 26518
rect 24492 26454 24544 26460
rect 24124 25424 24176 25430
rect 24124 25366 24176 25372
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 24044 24954 24072 25094
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 24136 24585 24164 25366
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24504 24818 24532 25162
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 24122 24576 24178 24585
rect 24122 24511 24178 24520
rect 24136 24206 24164 24511
rect 24308 24268 24360 24274
rect 24308 24210 24360 24216
rect 24124 24200 24176 24206
rect 24124 24142 24176 24148
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24216 23180 24268 23186
rect 24216 23122 24268 23128
rect 24044 22438 24072 23122
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23952 20806 23980 21082
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 24044 20482 24072 22374
rect 24228 21690 24256 23122
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 23952 20454 24072 20482
rect 23952 20330 23980 20454
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 23940 20324 23992 20330
rect 23940 20266 23992 20272
rect 23388 19926 23440 19932
rect 23676 19922 23888 19938
rect 23664 19916 23888 19922
rect 23716 19910 23888 19916
rect 23664 19858 23716 19864
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23308 19174 23336 19314
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23032 17746 23060 18770
rect 23308 18766 23336 19110
rect 23584 18970 23612 19246
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22572 16726 22600 17614
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22848 16726 22876 17274
rect 22940 17134 22968 17478
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 23032 16794 23060 17546
rect 23124 16794 23152 17682
rect 23308 17678 23336 18702
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22836 16720 22888 16726
rect 22836 16662 22888 16668
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 23032 15706 23060 16730
rect 23308 16726 23336 17614
rect 23676 17134 23704 18770
rect 23768 17814 23796 19790
rect 23860 18850 23888 19910
rect 23952 18970 23980 20266
rect 23940 18964 23992 18970
rect 23940 18906 23992 18912
rect 23860 18822 23980 18850
rect 24044 18834 24072 20334
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 23952 18698 23980 18822
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 23940 18692 23992 18698
rect 23940 18634 23992 18640
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 23756 17808 23808 17814
rect 23756 17750 23808 17756
rect 23664 17128 23716 17134
rect 23492 17076 23664 17082
rect 23492 17070 23716 17076
rect 23492 17054 23704 17070
rect 23492 16794 23520 17054
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23308 15162 23336 16662
rect 23492 16658 23520 16730
rect 23676 16658 23704 16934
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23768 15162 23796 17750
rect 24044 17270 24072 18566
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23952 16046 23980 16390
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22112 14618 22140 14894
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 24136 14498 24164 19858
rect 24228 19854 24256 20334
rect 24320 19922 24348 24210
rect 24596 23662 24624 26726
rect 24688 25226 24716 27338
rect 24780 26790 24808 31726
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24860 30388 24912 30394
rect 24860 30330 24912 30336
rect 24872 30190 24900 30330
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 24964 30122 24992 31078
rect 24952 30116 25004 30122
rect 24952 30058 25004 30064
rect 24964 30002 24992 30058
rect 24872 29974 24992 30002
rect 24872 28150 24900 29974
rect 24952 28416 25004 28422
rect 24952 28358 25004 28364
rect 24964 28218 24992 28358
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 24860 27600 24912 27606
rect 24860 27542 24912 27548
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 24872 25498 24900 27542
rect 24964 27062 24992 28154
rect 25056 27674 25084 32846
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25136 31680 25188 31686
rect 25136 31622 25188 31628
rect 25148 29646 25176 31622
rect 25228 30592 25280 30598
rect 25228 30534 25280 30540
rect 25240 30326 25268 30534
rect 25228 30320 25280 30326
rect 25228 30262 25280 30268
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 25136 29640 25188 29646
rect 25136 29582 25188 29588
rect 25148 29102 25176 29582
rect 25240 29102 25268 29650
rect 25136 29096 25188 29102
rect 25136 29038 25188 29044
rect 25228 29096 25280 29102
rect 25228 29038 25280 29044
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 25148 27538 25176 27814
rect 25136 27532 25188 27538
rect 25136 27474 25188 27480
rect 25228 27532 25280 27538
rect 25228 27474 25280 27480
rect 24952 27056 25004 27062
rect 24952 26998 25004 27004
rect 25240 26926 25268 27474
rect 25332 26926 25360 32166
rect 25516 31754 25544 32710
rect 26252 32366 26280 33374
rect 26344 33046 26372 33798
rect 26424 33380 26476 33386
rect 26424 33322 26476 33328
rect 26436 33114 26464 33322
rect 26424 33108 26476 33114
rect 26424 33050 26476 33056
rect 26332 33040 26384 33046
rect 26332 32982 26384 32988
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 26528 32212 26556 33866
rect 26608 32972 26660 32978
rect 26608 32914 26660 32920
rect 26252 32184 26556 32212
rect 25516 31726 25728 31754
rect 25596 30592 25648 30598
rect 25596 30534 25648 30540
rect 25608 30054 25636 30534
rect 25596 30048 25648 30054
rect 25596 29990 25648 29996
rect 25608 29306 25636 29990
rect 25596 29300 25648 29306
rect 25596 29242 25648 29248
rect 25608 28694 25636 29242
rect 25596 28688 25648 28694
rect 25596 28630 25648 28636
rect 25608 28098 25636 28630
rect 25516 28070 25636 28098
rect 25516 28014 25544 28070
rect 25504 28008 25556 28014
rect 25504 27950 25556 27956
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25412 26784 25464 26790
rect 25464 26744 25544 26772
rect 25412 26726 25464 26732
rect 25516 26518 25544 26744
rect 25504 26512 25556 26518
rect 25504 26454 25556 26460
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 25228 25424 25280 25430
rect 25228 25366 25280 25372
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 24688 24410 24716 24618
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24872 24206 24900 25094
rect 25240 24750 25268 25366
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25332 24750 25360 25230
rect 25516 24750 25544 26454
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25504 24744 25556 24750
rect 25504 24686 25556 24692
rect 25596 24744 25648 24750
rect 25596 24686 25648 24692
rect 25056 24410 25084 24686
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 25332 24018 25360 24686
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25424 24274 25452 24550
rect 25516 24410 25544 24686
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25608 24274 25636 24686
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25240 23990 25360 24018
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24504 22710 24532 23054
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24412 22098 24440 22510
rect 24400 22092 24452 22098
rect 24400 22034 24452 22040
rect 24596 21554 24624 23598
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24688 22574 24716 23122
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24688 22234 24716 22510
rect 25136 22500 25188 22506
rect 25136 22442 25188 22448
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24676 22228 24728 22234
rect 24676 22170 24728 22176
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24688 21418 24716 22170
rect 24780 21554 24808 22374
rect 25148 22234 25176 22442
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24872 21468 24900 21830
rect 24952 21480 25004 21486
rect 24872 21440 24952 21468
rect 24676 21412 24728 21418
rect 24676 21354 24728 21360
rect 24872 20942 24900 21440
rect 24952 21422 25004 21428
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 21146 25176 21422
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24308 19916 24360 19922
rect 24308 19858 24360 19864
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24412 18970 24440 19246
rect 24492 19236 24544 19242
rect 24492 19178 24544 19184
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24504 18834 24532 19178
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 24504 18222 24532 18770
rect 24492 18216 24544 18222
rect 24492 18158 24544 18164
rect 24504 17746 24532 18158
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 16658 24256 17478
rect 24306 17368 24362 17377
rect 24306 17303 24362 17312
rect 24320 17270 24348 17303
rect 24308 17264 24360 17270
rect 24308 17206 24360 17212
rect 24412 17134 24440 17614
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24216 16652 24268 16658
rect 24216 16594 24268 16600
rect 24044 14482 24164 14498
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 24032 14476 24164 14482
rect 24084 14470 24164 14476
rect 24216 14476 24268 14482
rect 24032 14418 24084 14424
rect 24216 14418 24268 14424
rect 19210 14172 19518 14181
rect 19210 14170 19216 14172
rect 19272 14170 19296 14172
rect 19352 14170 19376 14172
rect 19432 14170 19456 14172
rect 19512 14170 19518 14172
rect 19272 14118 19274 14170
rect 19454 14118 19456 14170
rect 19210 14116 19216 14118
rect 19272 14116 19296 14118
rect 19352 14116 19376 14118
rect 19432 14116 19456 14118
rect 19512 14116 19518 14118
rect 19210 14107 19518 14116
rect 19720 14074 19748 14418
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 23492 13802 23520 14214
rect 23584 14074 23612 14282
rect 24044 14074 24072 14418
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 19870 13628 20178 13637
rect 19870 13626 19876 13628
rect 19932 13626 19956 13628
rect 20012 13626 20036 13628
rect 20092 13626 20116 13628
rect 20172 13626 20178 13628
rect 19932 13574 19934 13626
rect 20114 13574 20116 13626
rect 19870 13572 19876 13574
rect 19932 13572 19956 13574
rect 20012 13572 20036 13574
rect 20092 13572 20116 13574
rect 20172 13572 20178 13574
rect 19870 13563 20178 13572
rect 23308 13530 23336 13738
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 24044 13462 24072 14010
rect 24228 13462 24256 14418
rect 24504 13870 24532 17682
rect 24596 17202 24624 20742
rect 24952 20528 25004 20534
rect 24952 20470 25004 20476
rect 24964 19922 24992 20470
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 25240 19530 25268 23990
rect 25412 23248 25464 23254
rect 25412 23190 25464 23196
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25332 22234 25360 22918
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25332 21418 25360 22170
rect 25424 21962 25452 23190
rect 25504 22092 25556 22098
rect 25504 22034 25556 22040
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 25516 21622 25544 22034
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25504 21616 25556 21622
rect 25504 21558 25556 21564
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25320 21412 25372 21418
rect 25320 21354 25372 21360
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 25320 19984 25372 19990
rect 25320 19926 25372 19932
rect 25148 19502 25268 19530
rect 25148 18834 25176 19502
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 25240 18902 25268 19382
rect 25332 19310 25360 19926
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25228 18896 25280 18902
rect 25228 18838 25280 18844
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 17338 24716 17682
rect 24780 17678 24808 18702
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24780 17066 24808 17614
rect 24872 17134 24900 18566
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 25148 17082 25176 18770
rect 24768 17060 24820 17066
rect 24768 17002 24820 17008
rect 25056 16794 25084 17070
rect 25148 17054 25268 17082
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25148 16250 25176 16934
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24780 14346 24808 14418
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24872 13462 24900 14214
rect 24964 14074 24992 14486
rect 25056 14414 25084 14894
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25240 14278 25268 17054
rect 25424 14550 25452 21082
rect 25516 20398 25544 21422
rect 25608 20602 25636 21830
rect 25700 21690 25728 31726
rect 26056 31272 26108 31278
rect 26056 31214 26108 31220
rect 26068 30938 26096 31214
rect 26056 30932 26108 30938
rect 26056 30874 26108 30880
rect 25780 29572 25832 29578
rect 25780 29514 25832 29520
rect 25792 29170 25820 29514
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25872 29096 25924 29102
rect 25872 29038 25924 29044
rect 25964 29096 26016 29102
rect 25964 29038 26016 29044
rect 25884 28218 25912 29038
rect 25976 28490 26004 29038
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25792 27470 25820 27950
rect 25780 27464 25832 27470
rect 25780 27406 25832 27412
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25884 26790 25912 27338
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 25780 24676 25832 24682
rect 25780 24618 25832 24624
rect 25792 24274 25820 24618
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25700 21350 25728 21490
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25700 20330 25728 21286
rect 25792 20602 25820 24210
rect 25976 23866 26004 28426
rect 26056 27940 26108 27946
rect 26056 27882 26108 27888
rect 26068 27402 26096 27882
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26056 26920 26108 26926
rect 26056 26862 26108 26868
rect 26068 26314 26096 26862
rect 26056 26308 26108 26314
rect 26056 26250 26108 26256
rect 26160 25922 26188 27066
rect 26068 25894 26188 25922
rect 26068 24750 26096 25894
rect 26148 25424 26200 25430
rect 26148 25366 26200 25372
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 26068 24274 26096 24686
rect 26160 24342 26188 25366
rect 26252 24664 26280 32184
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 26344 31142 26372 31826
rect 26516 31680 26568 31686
rect 26516 31622 26568 31628
rect 26424 31340 26476 31346
rect 26424 31282 26476 31288
rect 26332 31136 26384 31142
rect 26332 31078 26384 31084
rect 26332 30932 26384 30938
rect 26332 30874 26384 30880
rect 26344 27470 26372 30874
rect 26436 30802 26464 31282
rect 26528 30802 26556 31622
rect 26424 30796 26476 30802
rect 26424 30738 26476 30744
rect 26516 30796 26568 30802
rect 26516 30738 26568 30744
rect 26516 29844 26568 29850
rect 26516 29786 26568 29792
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 26332 27328 26384 27334
rect 26332 27270 26384 27276
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 26344 27130 26372 27270
rect 26436 27130 26464 27270
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26424 27124 26476 27130
rect 26424 27066 26476 27072
rect 26528 26976 26556 29786
rect 26620 29782 26648 32914
rect 26700 31884 26752 31890
rect 26700 31826 26752 31832
rect 26712 31210 26740 31826
rect 26700 31204 26752 31210
rect 26700 31146 26752 31152
rect 26712 30705 26740 31146
rect 26698 30696 26754 30705
rect 26698 30631 26754 30640
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26608 29776 26660 29782
rect 26608 29718 26660 29724
rect 26712 29714 26740 30534
rect 26804 29850 26832 34070
rect 26896 32978 26924 34190
rect 28000 34134 28028 34886
rect 28368 34746 28396 35090
rect 28356 34740 28408 34746
rect 28356 34682 28408 34688
rect 27344 34128 27396 34134
rect 27344 34070 27396 34076
rect 27988 34128 28040 34134
rect 27988 34070 28040 34076
rect 26984 33756 27292 33765
rect 26984 33754 26990 33756
rect 27046 33754 27070 33756
rect 27126 33754 27150 33756
rect 27206 33754 27230 33756
rect 27286 33754 27292 33756
rect 27046 33702 27048 33754
rect 27228 33702 27230 33754
rect 26984 33700 26990 33702
rect 27046 33700 27070 33702
rect 27126 33700 27150 33702
rect 27206 33700 27230 33702
rect 27286 33700 27292 33702
rect 26984 33691 27292 33700
rect 27356 33658 27384 34070
rect 27988 33924 28040 33930
rect 27988 33866 28040 33872
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27344 33652 27396 33658
rect 27344 33594 27396 33600
rect 27540 33114 27568 33798
rect 27644 33212 27952 33221
rect 27644 33210 27650 33212
rect 27706 33210 27730 33212
rect 27786 33210 27810 33212
rect 27866 33210 27890 33212
rect 27946 33210 27952 33212
rect 27706 33158 27708 33210
rect 27888 33158 27890 33210
rect 27644 33156 27650 33158
rect 27706 33156 27730 33158
rect 27786 33156 27810 33158
rect 27866 33156 27890 33158
rect 27946 33156 27952 33158
rect 27644 33147 27952 33156
rect 27528 33108 27580 33114
rect 27528 33050 27580 33056
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 27436 32972 27488 32978
rect 27436 32914 27488 32920
rect 26984 32668 27292 32677
rect 26984 32666 26990 32668
rect 27046 32666 27070 32668
rect 27126 32666 27150 32668
rect 27206 32666 27230 32668
rect 27286 32666 27292 32668
rect 27046 32614 27048 32666
rect 27228 32614 27230 32666
rect 26984 32612 26990 32614
rect 27046 32612 27070 32614
rect 27126 32612 27150 32614
rect 27206 32612 27230 32614
rect 27286 32612 27292 32614
rect 26984 32603 27292 32612
rect 27344 32292 27396 32298
rect 27344 32234 27396 32240
rect 26884 31748 26936 31754
rect 26884 31690 26936 31696
rect 26896 31278 26924 31690
rect 26984 31580 27292 31589
rect 26984 31578 26990 31580
rect 27046 31578 27070 31580
rect 27126 31578 27150 31580
rect 27206 31578 27230 31580
rect 27286 31578 27292 31580
rect 27046 31526 27048 31578
rect 27228 31526 27230 31578
rect 26984 31524 26990 31526
rect 27046 31524 27070 31526
rect 27126 31524 27150 31526
rect 27206 31524 27230 31526
rect 27286 31524 27292 31526
rect 26984 31515 27292 31524
rect 26884 31272 26936 31278
rect 26884 31214 26936 31220
rect 26884 31136 26936 31142
rect 26884 31078 26936 31084
rect 26976 31136 27028 31142
rect 26976 31078 27028 31084
rect 26896 30938 26924 31078
rect 26988 30938 27016 31078
rect 26884 30932 26936 30938
rect 26884 30874 26936 30880
rect 26976 30932 27028 30938
rect 26976 30874 27028 30880
rect 26984 30492 27292 30501
rect 26984 30490 26990 30492
rect 27046 30490 27070 30492
rect 27126 30490 27150 30492
rect 27206 30490 27230 30492
rect 27286 30490 27292 30492
rect 27046 30438 27048 30490
rect 27228 30438 27230 30490
rect 26984 30436 26990 30438
rect 27046 30436 27070 30438
rect 27126 30436 27150 30438
rect 27206 30436 27230 30438
rect 27286 30436 27292 30438
rect 26984 30427 27292 30436
rect 27356 30122 27384 32234
rect 27448 30870 27476 32914
rect 27896 32904 27948 32910
rect 28000 32892 28028 33866
rect 28460 33862 28488 35430
rect 28736 35018 28764 37062
rect 29184 36712 29236 36718
rect 29288 36700 29316 38354
rect 29460 37120 29512 37126
rect 29460 37062 29512 37068
rect 29236 36672 29316 36700
rect 29184 36654 29236 36660
rect 29472 36650 29500 37062
rect 29460 36644 29512 36650
rect 29460 36586 29512 36592
rect 29564 36038 29592 39374
rect 29932 39370 29960 39918
rect 30392 39846 30420 40326
rect 31036 39982 31064 40530
rect 30564 39976 30616 39982
rect 30564 39918 30616 39924
rect 31024 39976 31076 39982
rect 31024 39918 31076 39924
rect 30380 39840 30432 39846
rect 30380 39782 30432 39788
rect 30196 39500 30248 39506
rect 30196 39442 30248 39448
rect 29920 39364 29972 39370
rect 29920 39306 29972 39312
rect 29644 39296 29696 39302
rect 29644 39238 29696 39244
rect 29656 38894 29684 39238
rect 30208 39098 30236 39442
rect 30196 39092 30248 39098
rect 30196 39034 30248 39040
rect 30392 38894 30420 39782
rect 30576 39302 30604 39918
rect 30564 39296 30616 39302
rect 30564 39238 30616 39244
rect 29644 38888 29696 38894
rect 29644 38830 29696 38836
rect 30380 38888 30432 38894
rect 30380 38830 30432 38836
rect 30576 38826 30604 39238
rect 30564 38820 30616 38826
rect 30564 38762 30616 38768
rect 30472 37664 30524 37670
rect 30472 37606 30524 37612
rect 30484 37466 30512 37606
rect 30576 37466 30604 38762
rect 31116 37868 31168 37874
rect 31116 37810 31168 37816
rect 30472 37460 30524 37466
rect 30472 37402 30524 37408
rect 30564 37460 30616 37466
rect 30564 37402 30616 37408
rect 30196 37324 30248 37330
rect 30196 37266 30248 37272
rect 30012 36644 30064 36650
rect 30012 36586 30064 36592
rect 29644 36576 29696 36582
rect 29644 36518 29696 36524
rect 29656 36174 29684 36518
rect 30024 36378 30052 36586
rect 30012 36372 30064 36378
rect 30012 36314 30064 36320
rect 30208 36258 30236 37266
rect 30748 37256 30800 37262
rect 30748 37198 30800 37204
rect 30288 37188 30340 37194
rect 30288 37130 30340 37136
rect 30300 36922 30328 37130
rect 30564 37120 30616 37126
rect 30564 37062 30616 37068
rect 30288 36916 30340 36922
rect 30288 36858 30340 36864
rect 30300 36378 30328 36858
rect 30576 36582 30604 37062
rect 30564 36576 30616 36582
rect 30564 36518 30616 36524
rect 30288 36372 30340 36378
rect 30288 36314 30340 36320
rect 30208 36230 30328 36258
rect 30576 36242 30604 36518
rect 30300 36174 30328 36230
rect 30564 36236 30616 36242
rect 30564 36178 30616 36184
rect 29644 36168 29696 36174
rect 29644 36110 29696 36116
rect 30288 36168 30340 36174
rect 30288 36110 30340 36116
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 28908 35692 28960 35698
rect 28908 35634 28960 35640
rect 28920 35018 28948 35634
rect 29644 35624 29696 35630
rect 29644 35566 29696 35572
rect 29184 35284 29236 35290
rect 29184 35226 29236 35232
rect 28724 35012 28776 35018
rect 28724 34954 28776 34960
rect 28908 35012 28960 35018
rect 28908 34954 28960 34960
rect 28632 34944 28684 34950
rect 28632 34886 28684 34892
rect 28644 34542 28672 34886
rect 28632 34536 28684 34542
rect 28632 34478 28684 34484
rect 28920 33930 28948 34954
rect 29196 34066 29224 35226
rect 29656 35154 29684 35566
rect 30300 35290 30328 36110
rect 30760 36038 30788 37198
rect 31128 37194 31156 37810
rect 31300 37460 31352 37466
rect 31300 37402 31352 37408
rect 31312 37330 31340 37402
rect 31300 37324 31352 37330
rect 31300 37266 31352 37272
rect 31024 37188 31076 37194
rect 31024 37130 31076 37136
rect 31116 37188 31168 37194
rect 31116 37130 31168 37136
rect 31036 36378 31064 37130
rect 31024 36372 31076 36378
rect 31024 36314 31076 36320
rect 31300 36372 31352 36378
rect 31300 36314 31352 36320
rect 30748 36032 30800 36038
rect 30748 35974 30800 35980
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 30196 35216 30248 35222
rect 30196 35158 30248 35164
rect 29644 35148 29696 35154
rect 29644 35090 29696 35096
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 29656 35034 29684 35090
rect 29564 35006 29684 35034
rect 29276 34468 29328 34474
rect 29276 34410 29328 34416
rect 29288 34202 29316 34410
rect 29276 34196 29328 34202
rect 29276 34138 29328 34144
rect 29184 34060 29236 34066
rect 29184 34002 29236 34008
rect 29564 33998 29592 35006
rect 29748 34898 29776 35090
rect 29920 35012 29972 35018
rect 29920 34954 29972 34960
rect 29656 34870 29776 34898
rect 29656 34746 29684 34870
rect 29644 34740 29696 34746
rect 29644 34682 29696 34688
rect 29736 34740 29788 34746
rect 29736 34682 29788 34688
rect 29656 34134 29684 34682
rect 29644 34128 29696 34134
rect 29644 34070 29696 34076
rect 29748 34066 29776 34682
rect 29932 34066 29960 34954
rect 30208 34746 30236 35158
rect 30564 35148 30616 35154
rect 30564 35090 30616 35096
rect 30288 34944 30340 34950
rect 30288 34886 30340 34892
rect 30196 34740 30248 34746
rect 30196 34682 30248 34688
rect 30300 34134 30328 34886
rect 30576 34746 30604 35090
rect 30852 35086 30880 35430
rect 30840 35080 30892 35086
rect 30840 35022 30892 35028
rect 30564 34740 30616 34746
rect 30564 34682 30616 34688
rect 31312 34542 31340 36314
rect 31300 34536 31352 34542
rect 31300 34478 31352 34484
rect 31312 34202 31340 34478
rect 31300 34196 31352 34202
rect 31300 34138 31352 34144
rect 30288 34128 30340 34134
rect 30288 34070 30340 34076
rect 29736 34060 29788 34066
rect 29736 34002 29788 34008
rect 29920 34060 29972 34066
rect 29920 34002 29972 34008
rect 29552 33992 29604 33998
rect 29552 33934 29604 33940
rect 28908 33924 28960 33930
rect 28908 33866 28960 33872
rect 28448 33856 28500 33862
rect 28448 33798 28500 33804
rect 28356 33584 28408 33590
rect 28356 33526 28408 33532
rect 28080 33448 28132 33454
rect 28080 33390 28132 33396
rect 27948 32864 28028 32892
rect 27896 32846 27948 32852
rect 27712 32768 27764 32774
rect 27712 32710 27764 32716
rect 27724 32298 27752 32710
rect 27712 32292 27764 32298
rect 27712 32234 27764 32240
rect 27644 32124 27952 32133
rect 27644 32122 27650 32124
rect 27706 32122 27730 32124
rect 27786 32122 27810 32124
rect 27866 32122 27890 32124
rect 27946 32122 27952 32124
rect 27706 32070 27708 32122
rect 27888 32070 27890 32122
rect 27644 32068 27650 32070
rect 27706 32068 27730 32070
rect 27786 32068 27810 32070
rect 27866 32068 27890 32070
rect 27946 32068 27952 32070
rect 27644 32059 27952 32068
rect 28000 31754 28028 32864
rect 28092 32026 28120 33390
rect 28368 32978 28396 33526
rect 28460 33522 28488 33798
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28356 32972 28408 32978
rect 28356 32914 28408 32920
rect 28460 32842 28488 33458
rect 28920 33454 28948 33866
rect 29564 33522 29592 33934
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 28908 33448 28960 33454
rect 28908 33390 28960 33396
rect 28920 33046 28948 33390
rect 29092 33312 29144 33318
rect 29092 33254 29144 33260
rect 29104 33114 29132 33254
rect 29092 33108 29144 33114
rect 29092 33050 29144 33056
rect 28908 33040 28960 33046
rect 28908 32982 28960 32988
rect 28448 32836 28500 32842
rect 28448 32778 28500 32784
rect 28920 32570 28948 32982
rect 29000 32768 29052 32774
rect 29000 32710 29052 32716
rect 28908 32564 28960 32570
rect 28908 32506 28960 32512
rect 28080 32020 28132 32026
rect 28080 31962 28132 31968
rect 29012 31958 29040 32710
rect 29368 32224 29420 32230
rect 29368 32166 29420 32172
rect 29000 31952 29052 31958
rect 29000 31894 29052 31900
rect 29380 31890 29408 32166
rect 29368 31884 29420 31890
rect 29368 31826 29420 31832
rect 28000 31726 28120 31754
rect 27988 31272 28040 31278
rect 27988 31214 28040 31220
rect 27528 31136 27580 31142
rect 27528 31078 27580 31084
rect 27436 30864 27488 30870
rect 27436 30806 27488 30812
rect 27540 30802 27568 31078
rect 27644 31036 27952 31045
rect 27644 31034 27650 31036
rect 27706 31034 27730 31036
rect 27786 31034 27810 31036
rect 27866 31034 27890 31036
rect 27946 31034 27952 31036
rect 27706 30982 27708 31034
rect 27888 30982 27890 31034
rect 27644 30980 27650 30982
rect 27706 30980 27730 30982
rect 27786 30980 27810 30982
rect 27866 30980 27890 30982
rect 27946 30980 27952 30982
rect 27644 30971 27952 30980
rect 28000 30802 28028 31214
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27988 30796 28040 30802
rect 27988 30738 28040 30744
rect 27988 30592 28040 30598
rect 27988 30534 28040 30540
rect 27344 30116 27396 30122
rect 27344 30058 27396 30064
rect 27528 30116 27580 30122
rect 27528 30058 27580 30064
rect 26792 29844 26844 29850
rect 26792 29786 26844 29792
rect 26700 29708 26752 29714
rect 26700 29650 26752 29656
rect 26608 29640 26660 29646
rect 26608 29582 26660 29588
rect 26792 29640 26844 29646
rect 26792 29582 26844 29588
rect 26436 26948 26556 26976
rect 26332 26920 26384 26926
rect 26436 26908 26464 26948
rect 26384 26880 26464 26908
rect 26332 26862 26384 26868
rect 26344 26450 26372 26862
rect 26516 26852 26568 26858
rect 26516 26794 26568 26800
rect 26528 26450 26556 26794
rect 26620 26586 26648 29582
rect 26804 28762 26832 29582
rect 26984 29404 27292 29413
rect 26984 29402 26990 29404
rect 27046 29402 27070 29404
rect 27126 29402 27150 29404
rect 27206 29402 27230 29404
rect 27286 29402 27292 29404
rect 27046 29350 27048 29402
rect 27228 29350 27230 29402
rect 26984 29348 26990 29350
rect 27046 29348 27070 29350
rect 27126 29348 27150 29350
rect 27206 29348 27230 29350
rect 27286 29348 27292 29350
rect 26984 29339 27292 29348
rect 26884 29232 26936 29238
rect 26884 29174 26936 29180
rect 26792 28756 26844 28762
rect 26792 28698 26844 28704
rect 26896 28626 26924 29174
rect 27356 29102 27384 30058
rect 27540 29832 27568 30058
rect 27644 29948 27952 29957
rect 27644 29946 27650 29948
rect 27706 29946 27730 29948
rect 27786 29946 27810 29948
rect 27866 29946 27890 29948
rect 27946 29946 27952 29948
rect 27706 29894 27708 29946
rect 27888 29894 27890 29946
rect 27644 29892 27650 29894
rect 27706 29892 27730 29894
rect 27786 29892 27810 29894
rect 27866 29892 27890 29894
rect 27946 29892 27952 29894
rect 27644 29883 27952 29892
rect 27620 29844 27672 29850
rect 27540 29804 27620 29832
rect 27620 29786 27672 29792
rect 27436 29640 27488 29646
rect 27436 29582 27488 29588
rect 27344 29096 27396 29102
rect 27344 29038 27396 29044
rect 26884 28620 26936 28626
rect 26884 28562 26936 28568
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 26792 28416 26844 28422
rect 26792 28358 26844 28364
rect 26700 27464 26752 27470
rect 26700 27406 26752 27412
rect 26712 26874 26740 27406
rect 26804 27130 26832 28358
rect 26984 28316 27292 28325
rect 26984 28314 26990 28316
rect 27046 28314 27070 28316
rect 27126 28314 27150 28316
rect 27206 28314 27230 28316
rect 27286 28314 27292 28316
rect 27046 28262 27048 28314
rect 27228 28262 27230 28314
rect 26984 28260 26990 28262
rect 27046 28260 27070 28262
rect 27126 28260 27150 28262
rect 27206 28260 27230 28262
rect 27286 28260 27292 28262
rect 26984 28251 27292 28260
rect 26884 27328 26936 27334
rect 26884 27270 26936 27276
rect 26792 27124 26844 27130
rect 26792 27066 26844 27072
rect 26712 26846 26832 26874
rect 26700 26784 26752 26790
rect 26700 26726 26752 26732
rect 26608 26580 26660 26586
rect 26608 26522 26660 26528
rect 26712 26518 26740 26726
rect 26804 26518 26832 26846
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 26792 26512 26844 26518
rect 26792 26454 26844 26460
rect 26896 26450 26924 27270
rect 26984 27228 27292 27237
rect 26984 27226 26990 27228
rect 27046 27226 27070 27228
rect 27126 27226 27150 27228
rect 27206 27226 27230 27228
rect 27286 27226 27292 27228
rect 27046 27174 27048 27226
rect 27228 27174 27230 27226
rect 26984 27172 26990 27174
rect 27046 27172 27070 27174
rect 27126 27172 27150 27174
rect 27206 27172 27230 27174
rect 27286 27172 27292 27174
rect 26984 27163 27292 27172
rect 26332 26444 26384 26450
rect 26332 26386 26384 26392
rect 26424 26444 26476 26450
rect 26424 26386 26476 26392
rect 26516 26444 26568 26450
rect 26516 26386 26568 26392
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26344 24834 26372 26250
rect 26436 25498 26464 26386
rect 26424 25492 26476 25498
rect 26424 25434 26476 25440
rect 26344 24806 26464 24834
rect 26332 24676 26384 24682
rect 26252 24636 26332 24664
rect 26332 24618 26384 24624
rect 26436 24614 26464 24806
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26148 24336 26200 24342
rect 26148 24278 26200 24284
rect 26056 24268 26108 24274
rect 26056 24210 26108 24216
rect 25964 23860 26016 23866
rect 25964 23802 26016 23808
rect 26160 22794 26188 24278
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 26240 24132 26292 24138
rect 26240 24074 26292 24080
rect 25884 22766 26188 22794
rect 25884 21350 25912 22766
rect 26252 22522 26280 24074
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 26344 22642 26372 23054
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26252 22494 26372 22522
rect 25964 22160 26016 22166
rect 25964 22102 26016 22108
rect 26238 22128 26294 22137
rect 25976 21622 26004 22102
rect 26056 22092 26108 22098
rect 26344 22098 26372 22494
rect 26436 22273 26464 24210
rect 26422 22264 26478 22273
rect 26422 22199 26478 22208
rect 26422 22128 26478 22137
rect 26238 22063 26294 22072
rect 26332 22092 26384 22098
rect 26056 22034 26108 22040
rect 25964 21616 26016 21622
rect 25964 21558 26016 21564
rect 26068 21468 26096 22034
rect 25976 21440 26096 21468
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25688 20324 25740 20330
rect 25688 20266 25740 20272
rect 25792 19922 25820 20538
rect 25872 20324 25924 20330
rect 25872 20266 25924 20272
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25700 17921 25728 19790
rect 25884 19718 25912 20266
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25976 19334 26004 21440
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 26068 19718 26096 20198
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 25792 19306 26004 19334
rect 25686 17912 25742 17921
rect 25686 17847 25742 17856
rect 25700 17746 25728 17847
rect 25792 17814 25820 19306
rect 26068 18970 26096 19654
rect 26160 19242 26188 21286
rect 26252 20346 26280 22063
rect 26422 22063 26478 22072
rect 26332 22034 26384 22040
rect 26344 21146 26372 22034
rect 26436 22030 26464 22063
rect 26424 22024 26476 22030
rect 26424 21966 26476 21972
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26436 21622 26464 21830
rect 26424 21616 26476 21622
rect 26424 21558 26476 21564
rect 26528 21570 26556 26386
rect 26792 26308 26844 26314
rect 26792 26250 26844 26256
rect 26608 24880 26660 24886
rect 26608 24822 26660 24828
rect 26620 24274 26648 24822
rect 26804 24750 26832 26250
rect 26984 26140 27292 26149
rect 26984 26138 26990 26140
rect 27046 26138 27070 26140
rect 27126 26138 27150 26140
rect 27206 26138 27230 26140
rect 27286 26138 27292 26140
rect 27046 26086 27048 26138
rect 27228 26086 27230 26138
rect 26984 26084 26990 26086
rect 27046 26084 27070 26086
rect 27126 26084 27150 26086
rect 27206 26084 27230 26086
rect 27286 26084 27292 26086
rect 26984 26075 27292 26084
rect 26984 25052 27292 25061
rect 26984 25050 26990 25052
rect 27046 25050 27070 25052
rect 27126 25050 27150 25052
rect 27206 25050 27230 25052
rect 27286 25050 27292 25052
rect 27046 24998 27048 25050
rect 27228 24998 27230 25050
rect 26984 24996 26990 24998
rect 27046 24996 27070 24998
rect 27126 24996 27150 24998
rect 27206 24996 27230 24998
rect 27286 24996 27292 24998
rect 26984 24987 27292 24996
rect 26792 24744 26844 24750
rect 26844 24704 26924 24732
rect 26792 24686 26844 24692
rect 26700 24676 26752 24682
rect 26700 24618 26752 24624
rect 26608 24268 26660 24274
rect 26608 24210 26660 24216
rect 26608 22976 26660 22982
rect 26608 22918 26660 22924
rect 26620 22166 26648 22918
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 26712 21962 26740 24618
rect 26792 23316 26844 23322
rect 26792 23258 26844 23264
rect 26804 22556 26832 23258
rect 26896 23050 26924 24704
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 27080 24070 27108 24550
rect 27356 24342 27384 28494
rect 27448 24954 27476 29582
rect 28000 29510 28028 30534
rect 28092 29850 28120 31726
rect 28448 30864 28500 30870
rect 28448 30806 28500 30812
rect 28080 29844 28132 29850
rect 28080 29786 28132 29792
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 28092 29050 28120 29786
rect 28460 29714 28488 30806
rect 28908 30796 28960 30802
rect 28908 30738 28960 30744
rect 28920 30054 28948 30738
rect 28908 30048 28960 30054
rect 28908 29990 28960 29996
rect 28448 29708 28500 29714
rect 28276 29668 28448 29696
rect 28172 29572 28224 29578
rect 28172 29514 28224 29520
rect 28000 29022 28120 29050
rect 28184 29034 28212 29514
rect 28172 29028 28224 29034
rect 27644 28860 27952 28869
rect 27644 28858 27650 28860
rect 27706 28858 27730 28860
rect 27786 28858 27810 28860
rect 27866 28858 27890 28860
rect 27946 28858 27952 28860
rect 27706 28806 27708 28858
rect 27888 28806 27890 28858
rect 27644 28804 27650 28806
rect 27706 28804 27730 28806
rect 27786 28804 27810 28806
rect 27866 28804 27890 28806
rect 27946 28804 27952 28806
rect 27644 28795 27952 28804
rect 27620 28008 27672 28014
rect 27540 27956 27620 27962
rect 27540 27950 27672 27956
rect 27540 27934 27660 27950
rect 28000 27946 28028 29022
rect 28172 28970 28224 28976
rect 28080 28960 28132 28966
rect 28080 28902 28132 28908
rect 28092 28422 28120 28902
rect 28276 28744 28304 29668
rect 28448 29650 28500 29656
rect 28920 29646 28948 29990
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28184 28716 28304 28744
rect 28080 28416 28132 28422
rect 28080 28358 28132 28364
rect 27988 27940 28040 27946
rect 27540 27538 27568 27934
rect 27988 27882 28040 27888
rect 27644 27772 27952 27781
rect 27644 27770 27650 27772
rect 27706 27770 27730 27772
rect 27786 27770 27810 27772
rect 27866 27770 27890 27772
rect 27946 27770 27952 27772
rect 27706 27718 27708 27770
rect 27888 27718 27890 27770
rect 27644 27716 27650 27718
rect 27706 27716 27730 27718
rect 27786 27716 27810 27718
rect 27866 27716 27890 27718
rect 27946 27716 27952 27718
rect 27644 27707 27952 27716
rect 27528 27532 27580 27538
rect 27528 27474 27580 27480
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27540 26790 27568 27338
rect 27988 26920 28040 26926
rect 27988 26862 28040 26868
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 27540 26450 27568 26726
rect 27644 26684 27952 26693
rect 27644 26682 27650 26684
rect 27706 26682 27730 26684
rect 27786 26682 27810 26684
rect 27866 26682 27890 26684
rect 27946 26682 27952 26684
rect 27706 26630 27708 26682
rect 27888 26630 27890 26682
rect 27644 26628 27650 26630
rect 27706 26628 27730 26630
rect 27786 26628 27810 26630
rect 27866 26628 27890 26630
rect 27946 26628 27952 26630
rect 27644 26619 27952 26628
rect 27712 26512 27764 26518
rect 27712 26454 27764 26460
rect 27528 26444 27580 26450
rect 27528 26386 27580 26392
rect 27540 25702 27568 26386
rect 27724 25809 27752 26454
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 27908 25838 27936 26318
rect 27896 25832 27948 25838
rect 27710 25800 27766 25809
rect 27896 25774 27948 25780
rect 27710 25735 27766 25744
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27436 24948 27488 24954
rect 27436 24890 27488 24896
rect 27540 24834 27568 25638
rect 27644 25596 27952 25605
rect 27644 25594 27650 25596
rect 27706 25594 27730 25596
rect 27786 25594 27810 25596
rect 27866 25594 27890 25596
rect 27946 25594 27952 25596
rect 27706 25542 27708 25594
rect 27888 25542 27890 25594
rect 27644 25540 27650 25542
rect 27706 25540 27730 25542
rect 27786 25540 27810 25542
rect 27866 25540 27890 25542
rect 27946 25540 27952 25542
rect 27644 25531 27952 25540
rect 28000 25362 28028 26862
rect 28092 26314 28120 27406
rect 28184 26586 28212 28716
rect 28264 28620 28316 28626
rect 28264 28562 28316 28568
rect 28276 28218 28304 28562
rect 28264 28212 28316 28218
rect 28264 28154 28316 28160
rect 28368 28150 28396 29106
rect 28448 28416 28500 28422
rect 28500 28376 28580 28404
rect 28448 28358 28500 28364
rect 28356 28144 28408 28150
rect 28356 28086 28408 28092
rect 28264 27940 28316 27946
rect 28264 27882 28316 27888
rect 28172 26580 28224 26586
rect 28172 26522 28224 26528
rect 28184 26314 28212 26522
rect 28276 26382 28304 27882
rect 28356 27532 28408 27538
rect 28356 27474 28408 27480
rect 28368 26586 28396 27474
rect 28448 26852 28500 26858
rect 28448 26794 28500 26800
rect 28356 26580 28408 26586
rect 28356 26522 28408 26528
rect 28460 26466 28488 26794
rect 28368 26438 28488 26466
rect 28264 26376 28316 26382
rect 28264 26318 28316 26324
rect 28080 26308 28132 26314
rect 28080 26250 28132 26256
rect 28172 26308 28224 26314
rect 28172 26250 28224 26256
rect 28092 25838 28120 26250
rect 28080 25832 28132 25838
rect 28080 25774 28132 25780
rect 28172 25696 28224 25702
rect 28078 25664 28134 25673
rect 28172 25638 28224 25644
rect 28078 25599 28134 25608
rect 27988 25356 28040 25362
rect 27988 25298 28040 25304
rect 28092 25242 28120 25599
rect 28000 25214 28120 25242
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 27448 24806 27568 24834
rect 27344 24336 27396 24342
rect 27344 24278 27396 24284
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27068 24064 27120 24070
rect 27068 24006 27120 24012
rect 26984 23964 27292 23973
rect 26984 23962 26990 23964
rect 27046 23962 27070 23964
rect 27126 23962 27150 23964
rect 27206 23962 27230 23964
rect 27286 23962 27292 23964
rect 27046 23910 27048 23962
rect 27228 23910 27230 23962
rect 26984 23908 26990 23910
rect 27046 23908 27070 23910
rect 27126 23908 27150 23910
rect 27206 23908 27230 23910
rect 27286 23908 27292 23910
rect 26984 23899 27292 23908
rect 26884 23044 26936 23050
rect 26884 22986 26936 22992
rect 26896 22692 26924 22986
rect 26984 22876 27292 22885
rect 26984 22874 26990 22876
rect 27046 22874 27070 22876
rect 27126 22874 27150 22876
rect 27206 22874 27230 22876
rect 27286 22874 27292 22876
rect 27046 22822 27048 22874
rect 27228 22822 27230 22874
rect 26984 22820 26990 22822
rect 27046 22820 27070 22822
rect 27126 22820 27150 22822
rect 27206 22820 27230 22822
rect 27286 22820 27292 22822
rect 26984 22811 27292 22820
rect 26896 22664 27016 22692
rect 26804 22528 26929 22556
rect 26901 22488 26929 22528
rect 26896 22460 26929 22488
rect 26792 22432 26844 22438
rect 26792 22374 26844 22380
rect 26804 22098 26832 22374
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 26700 21956 26752 21962
rect 26700 21898 26752 21904
rect 26528 21542 26740 21570
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 26252 20318 26464 20346
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 26252 19854 26280 19994
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26148 19236 26200 19242
rect 26148 19178 26200 19184
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 26056 18420 26108 18426
rect 26056 18362 26108 18368
rect 25780 17808 25832 17814
rect 25780 17750 25832 17756
rect 26068 17746 26096 18362
rect 25688 17740 25740 17746
rect 25688 17682 25740 17688
rect 26056 17740 26108 17746
rect 26056 17682 26108 17688
rect 25504 17604 25556 17610
rect 25504 17546 25556 17552
rect 25516 17134 25544 17546
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25608 16794 25636 17138
rect 26252 17134 26280 17478
rect 26344 17338 26372 19246
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 26436 17218 26464 20318
rect 26528 19514 26556 21422
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26620 19922 26648 20402
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26712 19802 26740 21542
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26620 19774 26740 19802
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 26528 17882 26556 18702
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26620 17338 26648 19774
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26712 19378 26740 19654
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26436 17190 26556 17218
rect 25964 17128 26016 17134
rect 25964 17070 26016 17076
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 25976 16998 26004 17070
rect 26436 16998 26464 17070
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25884 16658 25912 16934
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 26436 16454 26464 16934
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25700 14618 25728 14894
rect 26148 14816 26200 14822
rect 26148 14758 26200 14764
rect 26160 14618 26188 14758
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 25412 14544 25464 14550
rect 25464 14492 25544 14498
rect 25412 14486 25544 14492
rect 25424 14470 25544 14486
rect 26252 14482 26280 15846
rect 26436 15570 26464 16390
rect 26528 16182 26556 17190
rect 26804 16726 26832 21422
rect 26896 18834 26924 22460
rect 26988 22098 27016 22664
rect 27158 22672 27214 22681
rect 27158 22607 27160 22616
rect 27212 22607 27214 22616
rect 27160 22578 27212 22584
rect 27160 22500 27212 22506
rect 27160 22442 27212 22448
rect 27172 22166 27200 22442
rect 27160 22160 27212 22166
rect 27160 22102 27212 22108
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 26984 21788 27292 21797
rect 26984 21786 26990 21788
rect 27046 21786 27070 21788
rect 27126 21786 27150 21788
rect 27206 21786 27230 21788
rect 27286 21786 27292 21788
rect 27046 21734 27048 21786
rect 27228 21734 27230 21786
rect 26984 21732 26990 21734
rect 27046 21732 27070 21734
rect 27126 21732 27150 21734
rect 27206 21732 27230 21734
rect 27286 21732 27292 21734
rect 26984 21723 27292 21732
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27264 21146 27292 21626
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27356 21010 27384 24142
rect 27448 23322 27476 24806
rect 27528 24744 27580 24750
rect 27632 24732 27660 25094
rect 27580 24704 27660 24732
rect 27528 24686 27580 24692
rect 27528 24608 27580 24614
rect 27528 24550 27580 24556
rect 27540 24410 27568 24550
rect 27644 24508 27952 24517
rect 27644 24506 27650 24508
rect 27706 24506 27730 24508
rect 27786 24506 27810 24508
rect 27866 24506 27890 24508
rect 27946 24506 27952 24508
rect 27706 24454 27708 24506
rect 27888 24454 27890 24506
rect 27644 24452 27650 24454
rect 27706 24452 27730 24454
rect 27786 24452 27810 24454
rect 27866 24452 27890 24454
rect 27946 24452 27952 24454
rect 27644 24443 27952 24452
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 27436 23044 27488 23050
rect 27436 22986 27488 22992
rect 27448 22710 27476 22986
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27436 22568 27488 22574
rect 27436 22510 27488 22516
rect 27448 22234 27476 22510
rect 27436 22228 27488 22234
rect 27540 22216 27568 24210
rect 27632 23730 27660 24278
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27644 23420 27952 23429
rect 27644 23418 27650 23420
rect 27706 23418 27730 23420
rect 27786 23418 27810 23420
rect 27866 23418 27890 23420
rect 27946 23418 27952 23420
rect 27706 23366 27708 23418
rect 27888 23366 27890 23418
rect 27644 23364 27650 23366
rect 27706 23364 27730 23366
rect 27786 23364 27810 23366
rect 27866 23364 27890 23366
rect 27946 23364 27952 23366
rect 27644 23355 27952 23364
rect 28000 23254 28028 25214
rect 28080 24132 28132 24138
rect 28080 24074 28132 24080
rect 28092 23866 28120 24074
rect 28184 24070 28212 25638
rect 28276 24410 28304 26318
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28368 24274 28396 26438
rect 28448 26308 28500 26314
rect 28448 26250 28500 26256
rect 28460 24342 28488 26250
rect 28552 25809 28580 28376
rect 28920 26246 28948 29582
rect 29092 29028 29144 29034
rect 29092 28970 29144 28976
rect 29104 28626 29132 28970
rect 29092 28620 29144 28626
rect 29092 28562 29144 28568
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 29104 26858 29132 27270
rect 29092 26852 29144 26858
rect 29092 26794 29144 26800
rect 28908 26240 28960 26246
rect 28908 26182 28960 26188
rect 28816 25900 28868 25906
rect 28816 25842 28868 25848
rect 28538 25800 28594 25809
rect 28538 25735 28594 25744
rect 28632 25356 28684 25362
rect 28632 25298 28684 25304
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 28448 24336 28500 24342
rect 28448 24278 28500 24284
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 28172 24064 28224 24070
rect 28172 24006 28224 24012
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 28368 23866 28396 24006
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28448 23792 28500 23798
rect 28448 23734 28500 23740
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 28172 23656 28224 23662
rect 28172 23598 28224 23604
rect 28080 23520 28132 23526
rect 28080 23462 28132 23468
rect 28092 23254 28120 23462
rect 27988 23248 28040 23254
rect 27988 23190 28040 23196
rect 28080 23248 28132 23254
rect 28080 23190 28132 23196
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27632 22545 27660 23122
rect 28092 22982 28120 23190
rect 28184 22982 28212 23598
rect 28276 23050 28304 23666
rect 28356 23520 28408 23526
rect 28356 23462 28408 23468
rect 28368 23050 28396 23462
rect 28264 23044 28316 23050
rect 28264 22986 28316 22992
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28080 22976 28132 22982
rect 28080 22918 28132 22924
rect 28172 22976 28224 22982
rect 28172 22918 28224 22924
rect 27618 22536 27674 22545
rect 27618 22471 27674 22480
rect 27988 22432 28040 22438
rect 27988 22374 28040 22380
rect 27644 22332 27952 22341
rect 27644 22330 27650 22332
rect 27706 22330 27730 22332
rect 27786 22330 27810 22332
rect 27866 22330 27890 22332
rect 27946 22330 27952 22332
rect 27706 22278 27708 22330
rect 27888 22278 27890 22330
rect 27644 22276 27650 22278
rect 27706 22276 27730 22278
rect 27786 22276 27810 22278
rect 27866 22276 27890 22278
rect 27946 22276 27952 22278
rect 27644 22267 27952 22276
rect 28000 22216 28028 22374
rect 27540 22188 27660 22216
rect 27436 22170 27488 22176
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 26984 20700 27292 20709
rect 26984 20698 26990 20700
rect 27046 20698 27070 20700
rect 27126 20698 27150 20700
rect 27206 20698 27230 20700
rect 27286 20698 27292 20700
rect 27046 20646 27048 20698
rect 27228 20646 27230 20698
rect 26984 20644 26990 20646
rect 27046 20644 27070 20646
rect 27126 20644 27150 20646
rect 27206 20644 27230 20646
rect 27286 20644 27292 20646
rect 26984 20635 27292 20644
rect 27448 20330 27476 21966
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27344 19712 27396 19718
rect 27344 19654 27396 19660
rect 26984 19612 27292 19621
rect 26984 19610 26990 19612
rect 27046 19610 27070 19612
rect 27126 19610 27150 19612
rect 27206 19610 27230 19612
rect 27286 19610 27292 19612
rect 27046 19558 27048 19610
rect 27228 19558 27230 19610
rect 26984 19556 26990 19558
rect 27046 19556 27070 19558
rect 27126 19556 27150 19558
rect 27206 19556 27230 19558
rect 27286 19556 27292 19558
rect 26984 19547 27292 19556
rect 27356 19310 27384 19654
rect 27448 19446 27476 19790
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 26976 19304 27028 19310
rect 26976 19246 27028 19252
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 26988 18766 27016 19246
rect 26976 18760 27028 18766
rect 27436 18760 27488 18766
rect 26976 18702 27028 18708
rect 27356 18708 27436 18714
rect 27356 18702 27488 18708
rect 27356 18686 27476 18702
rect 26984 18524 27292 18533
rect 26984 18522 26990 18524
rect 27046 18522 27070 18524
rect 27126 18522 27150 18524
rect 27206 18522 27230 18524
rect 27286 18522 27292 18524
rect 27046 18470 27048 18522
rect 27228 18470 27230 18522
rect 26984 18468 26990 18470
rect 27046 18468 27070 18470
rect 27126 18468 27150 18470
rect 27206 18468 27230 18470
rect 27286 18468 27292 18470
rect 26984 18459 27292 18468
rect 26984 17436 27292 17445
rect 26984 17434 26990 17436
rect 27046 17434 27070 17436
rect 27126 17434 27150 17436
rect 27206 17434 27230 17436
rect 27286 17434 27292 17436
rect 27046 17382 27048 17434
rect 27228 17382 27230 17434
rect 26984 17380 26990 17382
rect 27046 17380 27070 17382
rect 27126 17380 27150 17382
rect 27206 17380 27230 17382
rect 27286 17380 27292 17382
rect 26984 17371 27292 17380
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27264 16794 27292 17070
rect 27356 16810 27384 18686
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27448 18222 27476 18566
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27540 17338 27568 22034
rect 27632 21690 27660 22188
rect 27908 22188 28028 22216
rect 27804 22160 27856 22166
rect 27804 22102 27856 22108
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27816 21486 27844 22102
rect 27908 22098 27936 22188
rect 27896 22092 27948 22098
rect 27896 22034 27948 22040
rect 27988 22092 28040 22098
rect 27988 22034 28040 22040
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 28000 21418 28028 22034
rect 28092 21894 28120 22918
rect 28184 22234 28212 22918
rect 28172 22228 28224 22234
rect 28172 22170 28224 22176
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 27988 21412 28040 21418
rect 27988 21354 28040 21360
rect 27644 21244 27952 21253
rect 27644 21242 27650 21244
rect 27706 21242 27730 21244
rect 27786 21242 27810 21244
rect 27866 21242 27890 21244
rect 27946 21242 27952 21244
rect 27706 21190 27708 21242
rect 27888 21190 27890 21242
rect 27644 21188 27650 21190
rect 27706 21188 27730 21190
rect 27786 21188 27810 21190
rect 27866 21188 27890 21190
rect 27946 21188 27952 21190
rect 27644 21179 27952 21188
rect 28000 21146 28028 21354
rect 28092 21350 28120 21830
rect 28172 21616 28224 21622
rect 28172 21558 28224 21564
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 27712 21140 27764 21146
rect 27712 21082 27764 21088
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 27724 20262 27752 21082
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 27816 20534 27844 20946
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 27804 20528 27856 20534
rect 27804 20470 27856 20476
rect 28000 20398 28028 20878
rect 28092 20602 28120 20946
rect 28080 20596 28132 20602
rect 28080 20538 28132 20544
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27644 20156 27952 20165
rect 27644 20154 27650 20156
rect 27706 20154 27730 20156
rect 27786 20154 27810 20156
rect 27866 20154 27890 20156
rect 27946 20154 27952 20156
rect 27706 20102 27708 20154
rect 27888 20102 27890 20154
rect 27644 20100 27650 20102
rect 27706 20100 27730 20102
rect 27786 20100 27810 20102
rect 27866 20100 27890 20102
rect 27946 20100 27952 20102
rect 27644 20091 27952 20100
rect 28000 19310 28028 20334
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 28092 19514 28120 20198
rect 28184 19922 28212 21558
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 27644 19068 27952 19077
rect 27644 19066 27650 19068
rect 27706 19066 27730 19068
rect 27786 19066 27810 19068
rect 27866 19066 27890 19068
rect 27946 19066 27952 19068
rect 27706 19014 27708 19066
rect 27888 19014 27890 19066
rect 27644 19012 27650 19014
rect 27706 19012 27730 19014
rect 27786 19012 27810 19014
rect 27866 19012 27890 19014
rect 27946 19012 27952 19014
rect 27644 19003 27952 19012
rect 28000 18426 28028 19246
rect 28092 18766 28120 19450
rect 28276 19242 28304 22986
rect 28460 22930 28488 23734
rect 28552 23254 28580 24346
rect 28644 23662 28672 25298
rect 28828 24954 28856 25842
rect 28816 24948 28868 24954
rect 28816 24890 28868 24896
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28736 23866 28764 24210
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28632 23656 28684 23662
rect 28632 23598 28684 23604
rect 28540 23248 28592 23254
rect 28540 23190 28592 23196
rect 28368 22902 28488 22930
rect 28368 21978 28396 22902
rect 28448 22432 28500 22438
rect 28448 22374 28500 22380
rect 28460 22098 28488 22374
rect 28448 22092 28500 22098
rect 28448 22034 28500 22040
rect 28368 21950 28488 21978
rect 28460 21894 28488 21950
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 28448 21888 28500 21894
rect 28448 21830 28500 21836
rect 28368 21486 28396 21830
rect 28460 21622 28488 21830
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 28368 20398 28396 21422
rect 28552 21418 28580 23190
rect 28644 22681 28672 23598
rect 28736 23322 28764 23802
rect 28724 23316 28776 23322
rect 28724 23258 28776 23264
rect 28828 23118 28856 24890
rect 28920 23186 28948 26182
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28724 23044 28776 23050
rect 28724 22986 28776 22992
rect 28630 22672 28686 22681
rect 28630 22607 28686 22616
rect 28644 22574 28672 22607
rect 28632 22568 28684 22574
rect 28632 22510 28684 22516
rect 28736 22386 28764 22986
rect 28816 22976 28868 22982
rect 28816 22918 28868 22924
rect 28644 22358 28764 22386
rect 28540 21412 28592 21418
rect 28540 21354 28592 21360
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28264 19236 28316 19242
rect 28264 19178 28316 19184
rect 28276 18766 28304 19178
rect 28460 19174 28488 20810
rect 28644 20806 28672 22358
rect 28724 22092 28776 22098
rect 28724 22034 28776 22040
rect 28736 21690 28764 22034
rect 28724 21684 28776 21690
rect 28724 21626 28776 21632
rect 28828 21434 28856 22918
rect 28736 21406 28856 21434
rect 28632 20800 28684 20806
rect 28632 20742 28684 20748
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28460 18834 28488 19110
rect 28552 18902 28580 19246
rect 28644 19174 28672 20742
rect 28736 20534 28764 21406
rect 28816 21344 28868 21350
rect 28816 21286 28868 21292
rect 28828 21010 28856 21286
rect 28816 21004 28868 21010
rect 28816 20946 28868 20952
rect 28724 20528 28776 20534
rect 28724 20470 28776 20476
rect 28920 19990 28948 23122
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 29012 21486 29040 22510
rect 29000 21480 29052 21486
rect 29000 21422 29052 21428
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 28540 18896 28592 18902
rect 28540 18838 28592 18844
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28644 18630 28672 19110
rect 29380 18902 29408 19110
rect 29368 18896 29420 18902
rect 29368 18838 29420 18844
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 28724 18692 28776 18698
rect 28724 18634 28776 18640
rect 28632 18624 28684 18630
rect 28632 18566 28684 18572
rect 27988 18420 28040 18426
rect 27988 18362 28040 18368
rect 28736 18086 28764 18634
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18222 29592 18566
rect 30392 18426 30420 18770
rect 30380 18420 30432 18426
rect 30380 18362 30432 18368
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 29552 18216 29604 18222
rect 29552 18158 29604 18164
rect 27988 18080 28040 18086
rect 27988 18022 28040 18028
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 27644 17980 27952 17989
rect 27644 17978 27650 17980
rect 27706 17978 27730 17980
rect 27786 17978 27810 17980
rect 27866 17978 27890 17980
rect 27946 17978 27952 17980
rect 27706 17926 27708 17978
rect 27888 17926 27890 17978
rect 27644 17924 27650 17926
rect 27706 17924 27730 17926
rect 27786 17924 27810 17926
rect 27866 17924 27890 17926
rect 27946 17924 27952 17926
rect 27644 17915 27952 17924
rect 28000 17746 28028 18022
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27644 16892 27952 16901
rect 27644 16890 27650 16892
rect 27706 16890 27730 16892
rect 27786 16890 27810 16892
rect 27866 16890 27890 16892
rect 27946 16890 27952 16892
rect 27706 16838 27708 16890
rect 27888 16838 27890 16890
rect 27644 16836 27650 16838
rect 27706 16836 27730 16838
rect 27786 16836 27810 16838
rect 27866 16836 27890 16838
rect 27946 16836 27952 16838
rect 27644 16827 27952 16836
rect 27252 16788 27304 16794
rect 27252 16730 27304 16736
rect 27356 16782 27568 16810
rect 26792 16720 26844 16726
rect 26792 16662 26844 16668
rect 26882 16688 26938 16697
rect 26516 16176 26568 16182
rect 26516 16118 26568 16124
rect 26700 16176 26752 16182
rect 26700 16118 26752 16124
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26436 14958 26464 15506
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 26620 15162 26648 15302
rect 26712 15162 26740 16118
rect 26804 16046 26832 16662
rect 26882 16623 26884 16632
rect 26936 16623 26938 16632
rect 26884 16594 26936 16600
rect 26792 16040 26844 16046
rect 26792 15982 26844 15988
rect 26896 15978 26924 16594
rect 27264 16538 27292 16730
rect 27356 16658 27384 16782
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27264 16510 27384 16538
rect 26984 16348 27292 16357
rect 26984 16346 26990 16348
rect 27046 16346 27070 16348
rect 27126 16346 27150 16348
rect 27206 16346 27230 16348
rect 27286 16346 27292 16348
rect 27046 16294 27048 16346
rect 27228 16294 27230 16346
rect 26984 16292 26990 16294
rect 27046 16292 27070 16294
rect 27126 16292 27150 16294
rect 27206 16292 27230 16294
rect 27286 16292 27292 16294
rect 26984 16283 27292 16292
rect 27356 16046 27384 16510
rect 27448 16250 27476 16594
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27344 16040 27396 16046
rect 27344 15982 27396 15988
rect 26884 15972 26936 15978
rect 26884 15914 26936 15920
rect 26896 15434 26924 15914
rect 27344 15564 27396 15570
rect 27344 15506 27396 15512
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26712 14890 26740 15098
rect 26700 14884 26752 14890
rect 26700 14826 26752 14832
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25240 13802 25268 14214
rect 25516 13870 25544 14470
rect 25964 14476 26016 14482
rect 26240 14476 26292 14482
rect 25964 14418 26016 14424
rect 26160 14436 26240 14464
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25228 13796 25280 13802
rect 25228 13738 25280 13744
rect 24032 13456 24084 13462
rect 24032 13398 24084 13404
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16868 11354 16896 11630
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 18892 11218 18920 12718
rect 18984 12102 19012 13194
rect 19210 13084 19518 13093
rect 19210 13082 19216 13084
rect 19272 13082 19296 13084
rect 19352 13082 19376 13084
rect 19432 13082 19456 13084
rect 19512 13082 19518 13084
rect 19272 13030 19274 13082
rect 19454 13030 19456 13082
rect 19210 13028 19216 13030
rect 19272 13028 19296 13030
rect 19352 13028 19376 13030
rect 19432 13028 19456 13030
rect 19512 13028 19518 13030
rect 19210 13019 19518 13028
rect 25240 12714 25268 13738
rect 25516 13530 25544 13806
rect 25700 13802 25728 13942
rect 25976 13938 26004 14418
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25792 13394 25820 13806
rect 26160 13802 26188 14436
rect 26240 14418 26292 14424
rect 26804 14414 26832 15302
rect 26984 15260 27292 15269
rect 26984 15258 26990 15260
rect 27046 15258 27070 15260
rect 27126 15258 27150 15260
rect 27206 15258 27230 15260
rect 27286 15258 27292 15260
rect 27046 15206 27048 15258
rect 27228 15206 27230 15258
rect 26984 15204 26990 15206
rect 27046 15204 27070 15206
rect 27126 15204 27150 15206
rect 27206 15204 27230 15206
rect 27286 15204 27292 15206
rect 26984 15195 27292 15204
rect 27356 15162 27384 15506
rect 27448 15502 27476 16186
rect 27436 15496 27488 15502
rect 27436 15438 27488 15444
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27448 14958 27476 15438
rect 27540 15366 27568 16782
rect 28000 16658 28028 17682
rect 28736 17678 28764 18022
rect 29012 17882 29040 18158
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 28724 17672 28776 17678
rect 28724 17614 28776 17620
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 27988 16448 28040 16454
rect 27988 16390 28040 16396
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28000 16046 28028 16390
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 27644 15804 27952 15813
rect 27644 15802 27650 15804
rect 27706 15802 27730 15804
rect 27786 15802 27810 15804
rect 27866 15802 27890 15804
rect 27946 15802 27952 15804
rect 27706 15750 27708 15802
rect 27888 15750 27890 15802
rect 27644 15748 27650 15750
rect 27706 15748 27730 15750
rect 27786 15748 27810 15750
rect 27866 15748 27890 15750
rect 27946 15748 27952 15750
rect 27644 15739 27952 15748
rect 28736 15570 28764 16390
rect 29012 16046 29040 16594
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27644 14716 27952 14725
rect 27644 14714 27650 14716
rect 27706 14714 27730 14716
rect 27786 14714 27810 14716
rect 27866 14714 27890 14716
rect 27946 14714 27952 14716
rect 27706 14662 27708 14714
rect 27888 14662 27890 14714
rect 27644 14660 27650 14662
rect 27706 14660 27730 14662
rect 27786 14660 27810 14662
rect 27866 14660 27890 14662
rect 27946 14660 27952 14662
rect 27644 14651 27952 14660
rect 26332 14408 26384 14414
rect 26332 14350 26384 14356
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26148 13796 26200 13802
rect 26148 13738 26200 13744
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 25872 13728 25924 13734
rect 25872 13670 25924 13676
rect 25780 13388 25832 13394
rect 25700 13348 25780 13376
rect 25700 12850 25728 13348
rect 25780 13330 25832 13336
rect 25884 13326 25912 13670
rect 26252 13394 26280 13738
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25792 12782 25820 13126
rect 26344 12918 26372 14350
rect 26984 14172 27292 14181
rect 26984 14170 26990 14172
rect 27046 14170 27070 14172
rect 27126 14170 27150 14172
rect 27206 14170 27230 14172
rect 27286 14170 27292 14172
rect 27046 14118 27048 14170
rect 27228 14118 27230 14170
rect 26984 14116 26990 14118
rect 27046 14116 27070 14118
rect 27126 14116 27150 14118
rect 27206 14116 27230 14118
rect 27286 14116 27292 14118
rect 26984 14107 27292 14116
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26436 13394 26464 13670
rect 27644 13628 27952 13637
rect 27644 13626 27650 13628
rect 27706 13626 27730 13628
rect 27786 13626 27810 13628
rect 27866 13626 27890 13628
rect 27946 13626 27952 13628
rect 27706 13574 27708 13626
rect 27888 13574 27890 13626
rect 27644 13572 27650 13574
rect 27706 13572 27730 13574
rect 27786 13572 27810 13574
rect 27866 13572 27890 13574
rect 27946 13572 27952 13574
rect 27644 13563 27952 13572
rect 28000 13530 28028 13874
rect 27988 13524 28040 13530
rect 27988 13466 28040 13472
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26528 12986 26556 13330
rect 26984 13084 27292 13093
rect 26984 13082 26990 13084
rect 27046 13082 27070 13084
rect 27126 13082 27150 13084
rect 27206 13082 27230 13084
rect 27286 13082 27292 13084
rect 27046 13030 27048 13082
rect 27228 13030 27230 13082
rect 26984 13028 26990 13030
rect 27046 13028 27070 13030
rect 27126 13028 27150 13030
rect 27206 13028 27230 13030
rect 27286 13028 27292 13030
rect 26984 13019 27292 13028
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26332 12912 26384 12918
rect 26332 12854 26384 12860
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 19870 12540 20178 12549
rect 19870 12538 19876 12540
rect 19932 12538 19956 12540
rect 20012 12538 20036 12540
rect 20092 12538 20116 12540
rect 20172 12538 20178 12540
rect 19932 12486 19934 12538
rect 20114 12486 20116 12538
rect 19870 12484 19876 12486
rect 19932 12484 19956 12486
rect 20012 12484 20036 12486
rect 20092 12484 20116 12486
rect 20172 12484 20178 12486
rect 19870 12475 20178 12484
rect 27644 12540 27952 12549
rect 27644 12538 27650 12540
rect 27706 12538 27730 12540
rect 27786 12538 27810 12540
rect 27866 12538 27890 12540
rect 27946 12538 27952 12540
rect 27706 12486 27708 12538
rect 27888 12486 27890 12538
rect 27644 12484 27650 12486
rect 27706 12484 27730 12486
rect 27786 12484 27810 12486
rect 27866 12484 27890 12486
rect 27946 12484 27952 12486
rect 27644 12475 27952 12484
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 19210 11996 19518 12005
rect 19210 11994 19216 11996
rect 19272 11994 19296 11996
rect 19352 11994 19376 11996
rect 19432 11994 19456 11996
rect 19512 11994 19518 11996
rect 19272 11942 19274 11994
rect 19454 11942 19456 11994
rect 19210 11940 19216 11942
rect 19272 11940 19296 11942
rect 19352 11940 19376 11942
rect 19432 11940 19456 11942
rect 19512 11940 19518 11942
rect 19210 11931 19518 11940
rect 26984 11996 27292 12005
rect 26984 11994 26990 11996
rect 27046 11994 27070 11996
rect 27126 11994 27150 11996
rect 27206 11994 27230 11996
rect 27286 11994 27292 11996
rect 27046 11942 27048 11994
rect 27228 11942 27230 11994
rect 26984 11940 26990 11942
rect 27046 11940 27070 11942
rect 27126 11940 27150 11942
rect 27206 11940 27230 11942
rect 27286 11940 27292 11942
rect 26984 11931 27292 11940
rect 19870 11452 20178 11461
rect 19870 11450 19876 11452
rect 19932 11450 19956 11452
rect 20012 11450 20036 11452
rect 20092 11450 20116 11452
rect 20172 11450 20178 11452
rect 19932 11398 19934 11450
rect 20114 11398 20116 11450
rect 19870 11396 19876 11398
rect 19932 11396 19956 11398
rect 20012 11396 20036 11398
rect 20092 11396 20116 11398
rect 20172 11396 20178 11398
rect 19870 11387 20178 11396
rect 27644 11452 27952 11461
rect 27644 11450 27650 11452
rect 27706 11450 27730 11452
rect 27786 11450 27810 11452
rect 27866 11450 27890 11452
rect 27946 11450 27952 11452
rect 27706 11398 27708 11450
rect 27888 11398 27890 11450
rect 27644 11396 27650 11398
rect 27706 11396 27730 11398
rect 27786 11396 27810 11398
rect 27866 11396 27890 11398
rect 27946 11396 27952 11398
rect 27644 11387 27952 11396
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 11436 10908 11744 10917
rect 11436 10906 11442 10908
rect 11498 10906 11522 10908
rect 11578 10906 11602 10908
rect 11658 10906 11682 10908
rect 11738 10906 11744 10908
rect 11498 10854 11500 10906
rect 11680 10854 11682 10906
rect 11436 10852 11442 10854
rect 11498 10852 11522 10854
rect 11578 10852 11602 10854
rect 11658 10852 11682 10854
rect 11738 10852 11744 10854
rect 11436 10843 11744 10852
rect 19210 10908 19518 10917
rect 19210 10906 19216 10908
rect 19272 10906 19296 10908
rect 19352 10906 19376 10908
rect 19432 10906 19456 10908
rect 19512 10906 19518 10908
rect 19272 10854 19274 10906
rect 19454 10854 19456 10906
rect 19210 10852 19216 10854
rect 19272 10852 19296 10854
rect 19352 10852 19376 10854
rect 19432 10852 19456 10854
rect 19512 10852 19518 10854
rect 19210 10843 19518 10852
rect 26984 10908 27292 10917
rect 26984 10906 26990 10908
rect 27046 10906 27070 10908
rect 27126 10906 27150 10908
rect 27206 10906 27230 10908
rect 27286 10906 27292 10908
rect 27046 10854 27048 10906
rect 27228 10854 27230 10906
rect 26984 10852 26990 10854
rect 27046 10852 27070 10854
rect 27126 10852 27150 10854
rect 27206 10852 27230 10854
rect 27286 10852 27292 10854
rect 26984 10843 27292 10852
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 12096 10364 12404 10373
rect 12096 10362 12102 10364
rect 12158 10362 12182 10364
rect 12238 10362 12262 10364
rect 12318 10362 12342 10364
rect 12398 10362 12404 10364
rect 12158 10310 12160 10362
rect 12340 10310 12342 10362
rect 12096 10308 12102 10310
rect 12158 10308 12182 10310
rect 12238 10308 12262 10310
rect 12318 10308 12342 10310
rect 12398 10308 12404 10310
rect 12096 10299 12404 10308
rect 19870 10364 20178 10373
rect 19870 10362 19876 10364
rect 19932 10362 19956 10364
rect 20012 10362 20036 10364
rect 20092 10362 20116 10364
rect 20172 10362 20178 10364
rect 19932 10310 19934 10362
rect 20114 10310 20116 10362
rect 19870 10308 19876 10310
rect 19932 10308 19956 10310
rect 20012 10308 20036 10310
rect 20092 10308 20116 10310
rect 20172 10308 20178 10310
rect 19870 10299 20178 10308
rect 27644 10364 27952 10373
rect 27644 10362 27650 10364
rect 27706 10362 27730 10364
rect 27786 10362 27810 10364
rect 27866 10362 27890 10364
rect 27946 10362 27952 10364
rect 27706 10310 27708 10362
rect 27888 10310 27890 10362
rect 27644 10308 27650 10310
rect 27706 10308 27730 10310
rect 27786 10308 27810 10310
rect 27866 10308 27890 10310
rect 27946 10308 27952 10310
rect 27644 10299 27952 10308
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 11436 9820 11744 9829
rect 11436 9818 11442 9820
rect 11498 9818 11522 9820
rect 11578 9818 11602 9820
rect 11658 9818 11682 9820
rect 11738 9818 11744 9820
rect 11498 9766 11500 9818
rect 11680 9766 11682 9818
rect 11436 9764 11442 9766
rect 11498 9764 11522 9766
rect 11578 9764 11602 9766
rect 11658 9764 11682 9766
rect 11738 9764 11744 9766
rect 11436 9755 11744 9764
rect 19210 9820 19518 9829
rect 19210 9818 19216 9820
rect 19272 9818 19296 9820
rect 19352 9818 19376 9820
rect 19432 9818 19456 9820
rect 19512 9818 19518 9820
rect 19272 9766 19274 9818
rect 19454 9766 19456 9818
rect 19210 9764 19216 9766
rect 19272 9764 19296 9766
rect 19352 9764 19376 9766
rect 19432 9764 19456 9766
rect 19512 9764 19518 9766
rect 19210 9755 19518 9764
rect 26984 9820 27292 9829
rect 26984 9818 26990 9820
rect 27046 9818 27070 9820
rect 27126 9818 27150 9820
rect 27206 9818 27230 9820
rect 27286 9818 27292 9820
rect 27046 9766 27048 9818
rect 27228 9766 27230 9818
rect 26984 9764 26990 9766
rect 27046 9764 27070 9766
rect 27126 9764 27150 9766
rect 27206 9764 27230 9766
rect 27286 9764 27292 9766
rect 26984 9755 27292 9764
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 12096 9276 12404 9285
rect 12096 9274 12102 9276
rect 12158 9274 12182 9276
rect 12238 9274 12262 9276
rect 12318 9274 12342 9276
rect 12398 9274 12404 9276
rect 12158 9222 12160 9274
rect 12340 9222 12342 9274
rect 12096 9220 12102 9222
rect 12158 9220 12182 9222
rect 12238 9220 12262 9222
rect 12318 9220 12342 9222
rect 12398 9220 12404 9222
rect 12096 9211 12404 9220
rect 19870 9276 20178 9285
rect 19870 9274 19876 9276
rect 19932 9274 19956 9276
rect 20012 9274 20036 9276
rect 20092 9274 20116 9276
rect 20172 9274 20178 9276
rect 19932 9222 19934 9274
rect 20114 9222 20116 9274
rect 19870 9220 19876 9222
rect 19932 9220 19956 9222
rect 20012 9220 20036 9222
rect 20092 9220 20116 9222
rect 20172 9220 20178 9222
rect 19870 9211 20178 9220
rect 27644 9276 27952 9285
rect 27644 9274 27650 9276
rect 27706 9274 27730 9276
rect 27786 9274 27810 9276
rect 27866 9274 27890 9276
rect 27946 9274 27952 9276
rect 27706 9222 27708 9274
rect 27888 9222 27890 9274
rect 27644 9220 27650 9222
rect 27706 9220 27730 9222
rect 27786 9220 27810 9222
rect 27866 9220 27890 9222
rect 27946 9220 27952 9222
rect 27644 9211 27952 9220
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 11436 8732 11744 8741
rect 11436 8730 11442 8732
rect 11498 8730 11522 8732
rect 11578 8730 11602 8732
rect 11658 8730 11682 8732
rect 11738 8730 11744 8732
rect 11498 8678 11500 8730
rect 11680 8678 11682 8730
rect 11436 8676 11442 8678
rect 11498 8676 11522 8678
rect 11578 8676 11602 8678
rect 11658 8676 11682 8678
rect 11738 8676 11744 8678
rect 11436 8667 11744 8676
rect 19210 8732 19518 8741
rect 19210 8730 19216 8732
rect 19272 8730 19296 8732
rect 19352 8730 19376 8732
rect 19432 8730 19456 8732
rect 19512 8730 19518 8732
rect 19272 8678 19274 8730
rect 19454 8678 19456 8730
rect 19210 8676 19216 8678
rect 19272 8676 19296 8678
rect 19352 8676 19376 8678
rect 19432 8676 19456 8678
rect 19512 8676 19518 8678
rect 19210 8667 19518 8676
rect 26984 8732 27292 8741
rect 26984 8730 26990 8732
rect 27046 8730 27070 8732
rect 27126 8730 27150 8732
rect 27206 8730 27230 8732
rect 27286 8730 27292 8732
rect 27046 8678 27048 8730
rect 27228 8678 27230 8730
rect 26984 8676 26990 8678
rect 27046 8676 27070 8678
rect 27126 8676 27150 8678
rect 27206 8676 27230 8678
rect 27286 8676 27292 8678
rect 26984 8667 27292 8676
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 12096 8188 12404 8197
rect 12096 8186 12102 8188
rect 12158 8186 12182 8188
rect 12238 8186 12262 8188
rect 12318 8186 12342 8188
rect 12398 8186 12404 8188
rect 12158 8134 12160 8186
rect 12340 8134 12342 8186
rect 12096 8132 12102 8134
rect 12158 8132 12182 8134
rect 12238 8132 12262 8134
rect 12318 8132 12342 8134
rect 12398 8132 12404 8134
rect 12096 8123 12404 8132
rect 19870 8188 20178 8197
rect 19870 8186 19876 8188
rect 19932 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20178 8188
rect 19932 8134 19934 8186
rect 20114 8134 20116 8186
rect 19870 8132 19876 8134
rect 19932 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20178 8134
rect 19870 8123 20178 8132
rect 27644 8188 27952 8197
rect 27644 8186 27650 8188
rect 27706 8186 27730 8188
rect 27786 8186 27810 8188
rect 27866 8186 27890 8188
rect 27946 8186 27952 8188
rect 27706 8134 27708 8186
rect 27888 8134 27890 8186
rect 27644 8132 27650 8134
rect 27706 8132 27730 8134
rect 27786 8132 27810 8134
rect 27866 8132 27890 8134
rect 27946 8132 27952 8134
rect 27644 8123 27952 8132
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 11436 7644 11744 7653
rect 11436 7642 11442 7644
rect 11498 7642 11522 7644
rect 11578 7642 11602 7644
rect 11658 7642 11682 7644
rect 11738 7642 11744 7644
rect 11498 7590 11500 7642
rect 11680 7590 11682 7642
rect 11436 7588 11442 7590
rect 11498 7588 11522 7590
rect 11578 7588 11602 7590
rect 11658 7588 11682 7590
rect 11738 7588 11744 7590
rect 11436 7579 11744 7588
rect 19210 7644 19518 7653
rect 19210 7642 19216 7644
rect 19272 7642 19296 7644
rect 19352 7642 19376 7644
rect 19432 7642 19456 7644
rect 19512 7642 19518 7644
rect 19272 7590 19274 7642
rect 19454 7590 19456 7642
rect 19210 7588 19216 7590
rect 19272 7588 19296 7590
rect 19352 7588 19376 7590
rect 19432 7588 19456 7590
rect 19512 7588 19518 7590
rect 19210 7579 19518 7588
rect 26984 7644 27292 7653
rect 26984 7642 26990 7644
rect 27046 7642 27070 7644
rect 27126 7642 27150 7644
rect 27206 7642 27230 7644
rect 27286 7642 27292 7644
rect 27046 7590 27048 7642
rect 27228 7590 27230 7642
rect 26984 7588 26990 7590
rect 27046 7588 27070 7590
rect 27126 7588 27150 7590
rect 27206 7588 27230 7590
rect 27286 7588 27292 7590
rect 26984 7579 27292 7588
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 12096 7100 12404 7109
rect 12096 7098 12102 7100
rect 12158 7098 12182 7100
rect 12238 7098 12262 7100
rect 12318 7098 12342 7100
rect 12398 7098 12404 7100
rect 12158 7046 12160 7098
rect 12340 7046 12342 7098
rect 12096 7044 12102 7046
rect 12158 7044 12182 7046
rect 12238 7044 12262 7046
rect 12318 7044 12342 7046
rect 12398 7044 12404 7046
rect 12096 7035 12404 7044
rect 19870 7100 20178 7109
rect 19870 7098 19876 7100
rect 19932 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20178 7100
rect 19932 7046 19934 7098
rect 20114 7046 20116 7098
rect 19870 7044 19876 7046
rect 19932 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20178 7046
rect 19870 7035 20178 7044
rect 27644 7100 27952 7109
rect 27644 7098 27650 7100
rect 27706 7098 27730 7100
rect 27786 7098 27810 7100
rect 27866 7098 27890 7100
rect 27946 7098 27952 7100
rect 27706 7046 27708 7098
rect 27888 7046 27890 7098
rect 27644 7044 27650 7046
rect 27706 7044 27730 7046
rect 27786 7044 27810 7046
rect 27866 7044 27890 7046
rect 27946 7044 27952 7046
rect 27644 7035 27952 7044
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 11436 6556 11744 6565
rect 11436 6554 11442 6556
rect 11498 6554 11522 6556
rect 11578 6554 11602 6556
rect 11658 6554 11682 6556
rect 11738 6554 11744 6556
rect 11498 6502 11500 6554
rect 11680 6502 11682 6554
rect 11436 6500 11442 6502
rect 11498 6500 11522 6502
rect 11578 6500 11602 6502
rect 11658 6500 11682 6502
rect 11738 6500 11744 6502
rect 11436 6491 11744 6500
rect 19210 6556 19518 6565
rect 19210 6554 19216 6556
rect 19272 6554 19296 6556
rect 19352 6554 19376 6556
rect 19432 6554 19456 6556
rect 19512 6554 19518 6556
rect 19272 6502 19274 6554
rect 19454 6502 19456 6554
rect 19210 6500 19216 6502
rect 19272 6500 19296 6502
rect 19352 6500 19376 6502
rect 19432 6500 19456 6502
rect 19512 6500 19518 6502
rect 19210 6491 19518 6500
rect 26984 6556 27292 6565
rect 26984 6554 26990 6556
rect 27046 6554 27070 6556
rect 27126 6554 27150 6556
rect 27206 6554 27230 6556
rect 27286 6554 27292 6556
rect 27046 6502 27048 6554
rect 27228 6502 27230 6554
rect 26984 6500 26990 6502
rect 27046 6500 27070 6502
rect 27126 6500 27150 6502
rect 27206 6500 27230 6502
rect 27286 6500 27292 6502
rect 26984 6491 27292 6500
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 12096 6012 12404 6021
rect 12096 6010 12102 6012
rect 12158 6010 12182 6012
rect 12238 6010 12262 6012
rect 12318 6010 12342 6012
rect 12398 6010 12404 6012
rect 12158 5958 12160 6010
rect 12340 5958 12342 6010
rect 12096 5956 12102 5958
rect 12158 5956 12182 5958
rect 12238 5956 12262 5958
rect 12318 5956 12342 5958
rect 12398 5956 12404 5958
rect 12096 5947 12404 5956
rect 19870 6012 20178 6021
rect 19870 6010 19876 6012
rect 19932 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20178 6012
rect 19932 5958 19934 6010
rect 20114 5958 20116 6010
rect 19870 5956 19876 5958
rect 19932 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20178 5958
rect 19870 5947 20178 5956
rect 27644 6012 27952 6021
rect 27644 6010 27650 6012
rect 27706 6010 27730 6012
rect 27786 6010 27810 6012
rect 27866 6010 27890 6012
rect 27946 6010 27952 6012
rect 27706 5958 27708 6010
rect 27888 5958 27890 6010
rect 27644 5956 27650 5958
rect 27706 5956 27730 5958
rect 27786 5956 27810 5958
rect 27866 5956 27890 5958
rect 27946 5956 27952 5958
rect 27644 5947 27952 5956
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 11436 5468 11744 5477
rect 11436 5466 11442 5468
rect 11498 5466 11522 5468
rect 11578 5466 11602 5468
rect 11658 5466 11682 5468
rect 11738 5466 11744 5468
rect 11498 5414 11500 5466
rect 11680 5414 11682 5466
rect 11436 5412 11442 5414
rect 11498 5412 11522 5414
rect 11578 5412 11602 5414
rect 11658 5412 11682 5414
rect 11738 5412 11744 5414
rect 11436 5403 11744 5412
rect 19210 5468 19518 5477
rect 19210 5466 19216 5468
rect 19272 5466 19296 5468
rect 19352 5466 19376 5468
rect 19432 5466 19456 5468
rect 19512 5466 19518 5468
rect 19272 5414 19274 5466
rect 19454 5414 19456 5466
rect 19210 5412 19216 5414
rect 19272 5412 19296 5414
rect 19352 5412 19376 5414
rect 19432 5412 19456 5414
rect 19512 5412 19518 5414
rect 19210 5403 19518 5412
rect 26984 5468 27292 5477
rect 26984 5466 26990 5468
rect 27046 5466 27070 5468
rect 27126 5466 27150 5468
rect 27206 5466 27230 5468
rect 27286 5466 27292 5468
rect 27046 5414 27048 5466
rect 27228 5414 27230 5466
rect 26984 5412 26990 5414
rect 27046 5412 27070 5414
rect 27126 5412 27150 5414
rect 27206 5412 27230 5414
rect 27286 5412 27292 5414
rect 26984 5403 27292 5412
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 12096 4924 12404 4933
rect 12096 4922 12102 4924
rect 12158 4922 12182 4924
rect 12238 4922 12262 4924
rect 12318 4922 12342 4924
rect 12398 4922 12404 4924
rect 12158 4870 12160 4922
rect 12340 4870 12342 4922
rect 12096 4868 12102 4870
rect 12158 4868 12182 4870
rect 12238 4868 12262 4870
rect 12318 4868 12342 4870
rect 12398 4868 12404 4870
rect 12096 4859 12404 4868
rect 19870 4924 20178 4933
rect 19870 4922 19876 4924
rect 19932 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20178 4924
rect 19932 4870 19934 4922
rect 20114 4870 20116 4922
rect 19870 4868 19876 4870
rect 19932 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20178 4870
rect 19870 4859 20178 4868
rect 27644 4924 27952 4933
rect 27644 4922 27650 4924
rect 27706 4922 27730 4924
rect 27786 4922 27810 4924
rect 27866 4922 27890 4924
rect 27946 4922 27952 4924
rect 27706 4870 27708 4922
rect 27888 4870 27890 4922
rect 27644 4868 27650 4870
rect 27706 4868 27730 4870
rect 27786 4868 27810 4870
rect 27866 4868 27890 4870
rect 27946 4868 27952 4870
rect 27644 4859 27952 4868
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 11436 4380 11744 4389
rect 11436 4378 11442 4380
rect 11498 4378 11522 4380
rect 11578 4378 11602 4380
rect 11658 4378 11682 4380
rect 11738 4378 11744 4380
rect 11498 4326 11500 4378
rect 11680 4326 11682 4378
rect 11436 4324 11442 4326
rect 11498 4324 11522 4326
rect 11578 4324 11602 4326
rect 11658 4324 11682 4326
rect 11738 4324 11744 4326
rect 11436 4315 11744 4324
rect 19210 4380 19518 4389
rect 19210 4378 19216 4380
rect 19272 4378 19296 4380
rect 19352 4378 19376 4380
rect 19432 4378 19456 4380
rect 19512 4378 19518 4380
rect 19272 4326 19274 4378
rect 19454 4326 19456 4378
rect 19210 4324 19216 4326
rect 19272 4324 19296 4326
rect 19352 4324 19376 4326
rect 19432 4324 19456 4326
rect 19512 4324 19518 4326
rect 19210 4315 19518 4324
rect 26984 4380 27292 4389
rect 26984 4378 26990 4380
rect 27046 4378 27070 4380
rect 27126 4378 27150 4380
rect 27206 4378 27230 4380
rect 27286 4378 27292 4380
rect 27046 4326 27048 4378
rect 27228 4326 27230 4378
rect 26984 4324 26990 4326
rect 27046 4324 27070 4326
rect 27126 4324 27150 4326
rect 27206 4324 27230 4326
rect 27286 4324 27292 4326
rect 26984 4315 27292 4324
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 12096 3836 12404 3845
rect 12096 3834 12102 3836
rect 12158 3834 12182 3836
rect 12238 3834 12262 3836
rect 12318 3834 12342 3836
rect 12398 3834 12404 3836
rect 12158 3782 12160 3834
rect 12340 3782 12342 3834
rect 12096 3780 12102 3782
rect 12158 3780 12182 3782
rect 12238 3780 12262 3782
rect 12318 3780 12342 3782
rect 12398 3780 12404 3782
rect 12096 3771 12404 3780
rect 19870 3836 20178 3845
rect 19870 3834 19876 3836
rect 19932 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20178 3836
rect 19932 3782 19934 3834
rect 20114 3782 20116 3834
rect 19870 3780 19876 3782
rect 19932 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20178 3782
rect 19870 3771 20178 3780
rect 27644 3836 27952 3845
rect 27644 3834 27650 3836
rect 27706 3834 27730 3836
rect 27786 3834 27810 3836
rect 27866 3834 27890 3836
rect 27946 3834 27952 3836
rect 27706 3782 27708 3834
rect 27888 3782 27890 3834
rect 27644 3780 27650 3782
rect 27706 3780 27730 3782
rect 27786 3780 27810 3782
rect 27866 3780 27890 3782
rect 27946 3780 27952 3782
rect 27644 3771 27952 3780
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 11436 3292 11744 3301
rect 11436 3290 11442 3292
rect 11498 3290 11522 3292
rect 11578 3290 11602 3292
rect 11658 3290 11682 3292
rect 11738 3290 11744 3292
rect 11498 3238 11500 3290
rect 11680 3238 11682 3290
rect 11436 3236 11442 3238
rect 11498 3236 11522 3238
rect 11578 3236 11602 3238
rect 11658 3236 11682 3238
rect 11738 3236 11744 3238
rect 11436 3227 11744 3236
rect 19210 3292 19518 3301
rect 19210 3290 19216 3292
rect 19272 3290 19296 3292
rect 19352 3290 19376 3292
rect 19432 3290 19456 3292
rect 19512 3290 19518 3292
rect 19272 3238 19274 3290
rect 19454 3238 19456 3290
rect 19210 3236 19216 3238
rect 19272 3236 19296 3238
rect 19352 3236 19376 3238
rect 19432 3236 19456 3238
rect 19512 3236 19518 3238
rect 19210 3227 19518 3236
rect 26984 3292 27292 3301
rect 26984 3290 26990 3292
rect 27046 3290 27070 3292
rect 27126 3290 27150 3292
rect 27206 3290 27230 3292
rect 27286 3290 27292 3292
rect 27046 3238 27048 3290
rect 27228 3238 27230 3290
rect 26984 3236 26990 3238
rect 27046 3236 27070 3238
rect 27126 3236 27150 3238
rect 27206 3236 27230 3238
rect 27286 3236 27292 3238
rect 26984 3227 27292 3236
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 12096 2748 12404 2757
rect 12096 2746 12102 2748
rect 12158 2746 12182 2748
rect 12238 2746 12262 2748
rect 12318 2746 12342 2748
rect 12398 2746 12404 2748
rect 12158 2694 12160 2746
rect 12340 2694 12342 2746
rect 12096 2692 12102 2694
rect 12158 2692 12182 2694
rect 12238 2692 12262 2694
rect 12318 2692 12342 2694
rect 12398 2692 12404 2694
rect 12096 2683 12404 2692
rect 19870 2748 20178 2757
rect 19870 2746 19876 2748
rect 19932 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20178 2748
rect 19932 2694 19934 2746
rect 20114 2694 20116 2746
rect 19870 2692 19876 2694
rect 19932 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20178 2694
rect 19870 2683 20178 2692
rect 27644 2748 27952 2757
rect 27644 2746 27650 2748
rect 27706 2746 27730 2748
rect 27786 2746 27810 2748
rect 27866 2746 27890 2748
rect 27946 2746 27952 2748
rect 27706 2694 27708 2746
rect 27888 2694 27890 2746
rect 27644 2692 27650 2694
rect 27706 2692 27730 2694
rect 27786 2692 27810 2694
rect 27866 2692 27890 2694
rect 27946 2692 27952 2694
rect 27644 2683 27952 2692
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 11436 2204 11744 2213
rect 11436 2202 11442 2204
rect 11498 2202 11522 2204
rect 11578 2202 11602 2204
rect 11658 2202 11682 2204
rect 11738 2202 11744 2204
rect 11498 2150 11500 2202
rect 11680 2150 11682 2202
rect 11436 2148 11442 2150
rect 11498 2148 11522 2150
rect 11578 2148 11602 2150
rect 11658 2148 11682 2150
rect 11738 2148 11744 2150
rect 11436 2139 11744 2148
rect 19210 2204 19518 2213
rect 19210 2202 19216 2204
rect 19272 2202 19296 2204
rect 19352 2202 19376 2204
rect 19432 2202 19456 2204
rect 19512 2202 19518 2204
rect 19272 2150 19274 2202
rect 19454 2150 19456 2202
rect 19210 2148 19216 2150
rect 19272 2148 19296 2150
rect 19352 2148 19376 2150
rect 19432 2148 19456 2150
rect 19512 2148 19518 2150
rect 19210 2139 19518 2148
rect 26984 2204 27292 2213
rect 26984 2202 26990 2204
rect 27046 2202 27070 2204
rect 27126 2202 27150 2204
rect 27206 2202 27230 2204
rect 27286 2202 27292 2204
rect 27046 2150 27048 2202
rect 27228 2150 27230 2202
rect 26984 2148 26990 2150
rect 27046 2148 27070 2150
rect 27126 2148 27150 2150
rect 27206 2148 27230 2150
rect 27286 2148 27292 2150
rect 26984 2139 27292 2148
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 12096 1660 12404 1669
rect 12096 1658 12102 1660
rect 12158 1658 12182 1660
rect 12238 1658 12262 1660
rect 12318 1658 12342 1660
rect 12398 1658 12404 1660
rect 12158 1606 12160 1658
rect 12340 1606 12342 1658
rect 12096 1604 12102 1606
rect 12158 1604 12182 1606
rect 12238 1604 12262 1606
rect 12318 1604 12342 1606
rect 12398 1604 12404 1606
rect 12096 1595 12404 1604
rect 19870 1660 20178 1669
rect 19870 1658 19876 1660
rect 19932 1658 19956 1660
rect 20012 1658 20036 1660
rect 20092 1658 20116 1660
rect 20172 1658 20178 1660
rect 19932 1606 19934 1658
rect 20114 1606 20116 1658
rect 19870 1604 19876 1606
rect 19932 1604 19956 1606
rect 20012 1604 20036 1606
rect 20092 1604 20116 1606
rect 20172 1604 20178 1606
rect 19870 1595 20178 1604
rect 27644 1660 27952 1669
rect 27644 1658 27650 1660
rect 27706 1658 27730 1660
rect 27786 1658 27810 1660
rect 27866 1658 27890 1660
rect 27946 1658 27952 1660
rect 27706 1606 27708 1658
rect 27888 1606 27890 1658
rect 27644 1604 27650 1606
rect 27706 1604 27730 1606
rect 27786 1604 27810 1606
rect 27866 1604 27890 1606
rect 27946 1604 27952 1606
rect 27644 1595 27952 1604
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 11436 1116 11744 1125
rect 11436 1114 11442 1116
rect 11498 1114 11522 1116
rect 11578 1114 11602 1116
rect 11658 1114 11682 1116
rect 11738 1114 11744 1116
rect 11498 1062 11500 1114
rect 11680 1062 11682 1114
rect 11436 1060 11442 1062
rect 11498 1060 11522 1062
rect 11578 1060 11602 1062
rect 11658 1060 11682 1062
rect 11738 1060 11744 1062
rect 11436 1051 11744 1060
rect 19210 1116 19518 1125
rect 19210 1114 19216 1116
rect 19272 1114 19296 1116
rect 19352 1114 19376 1116
rect 19432 1114 19456 1116
rect 19512 1114 19518 1116
rect 19272 1062 19274 1114
rect 19454 1062 19456 1114
rect 19210 1060 19216 1062
rect 19272 1060 19296 1062
rect 19352 1060 19376 1062
rect 19432 1060 19456 1062
rect 19512 1060 19518 1062
rect 19210 1051 19518 1060
rect 26984 1116 27292 1125
rect 26984 1114 26990 1116
rect 27046 1114 27070 1116
rect 27126 1114 27150 1116
rect 27206 1114 27230 1116
rect 27286 1114 27292 1116
rect 27046 1062 27048 1114
rect 27228 1062 27230 1114
rect 26984 1060 26990 1062
rect 27046 1060 27070 1062
rect 27126 1060 27150 1062
rect 27206 1060 27230 1062
rect 27286 1060 27292 1062
rect 26984 1051 27292 1060
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 12096 572 12404 581
rect 12096 570 12102 572
rect 12158 570 12182 572
rect 12238 570 12262 572
rect 12318 570 12342 572
rect 12398 570 12404 572
rect 12158 518 12160 570
rect 12340 518 12342 570
rect 12096 516 12102 518
rect 12158 516 12182 518
rect 12238 516 12262 518
rect 12318 516 12342 518
rect 12398 516 12404 518
rect 12096 507 12404 516
rect 19870 572 20178 581
rect 19870 570 19876 572
rect 19932 570 19956 572
rect 20012 570 20036 572
rect 20092 570 20116 572
rect 20172 570 20178 572
rect 19932 518 19934 570
rect 20114 518 20116 570
rect 19870 516 19876 518
rect 19932 516 19956 518
rect 20012 516 20036 518
rect 20092 516 20116 518
rect 20172 516 20178 518
rect 19870 507 20178 516
rect 27644 572 27952 581
rect 27644 570 27650 572
rect 27706 570 27730 572
rect 27786 570 27810 572
rect 27866 570 27890 572
rect 27946 570 27952 572
rect 27706 518 27708 570
rect 27888 518 27890 570
rect 27644 516 27650 518
rect 27706 516 27730 518
rect 27786 516 27810 518
rect 27866 516 27890 518
rect 27946 516 27952 518
rect 27644 507 27952 516
<< via2 >>
rect 11794 44784 11850 44840
rect 13082 44784 13138 44840
rect 21638 44784 21694 44840
rect 27434 44784 27490 44840
rect 28170 44784 28226 44840
rect 3668 44634 3724 44636
rect 3748 44634 3804 44636
rect 3828 44634 3884 44636
rect 3908 44634 3964 44636
rect 3668 44582 3714 44634
rect 3714 44582 3724 44634
rect 3748 44582 3778 44634
rect 3778 44582 3790 44634
rect 3790 44582 3804 44634
rect 3828 44582 3842 44634
rect 3842 44582 3854 44634
rect 3854 44582 3884 44634
rect 3908 44582 3918 44634
rect 3918 44582 3964 44634
rect 3668 44580 3724 44582
rect 3748 44580 3804 44582
rect 3828 44580 3884 44582
rect 3908 44580 3964 44582
rect 11442 44634 11498 44636
rect 11522 44634 11578 44636
rect 11602 44634 11658 44636
rect 11682 44634 11738 44636
rect 11442 44582 11488 44634
rect 11488 44582 11498 44634
rect 11522 44582 11552 44634
rect 11552 44582 11564 44634
rect 11564 44582 11578 44634
rect 11602 44582 11616 44634
rect 11616 44582 11628 44634
rect 11628 44582 11658 44634
rect 11682 44582 11692 44634
rect 11692 44582 11738 44634
rect 11442 44580 11498 44582
rect 11522 44580 11578 44582
rect 11602 44580 11658 44582
rect 11682 44580 11738 44582
rect 7194 44532 7250 44568
rect 7194 44512 7196 44532
rect 7196 44512 7248 44532
rect 7248 44512 7250 44532
rect 7654 44532 7710 44568
rect 7654 44512 7656 44532
rect 7656 44512 7708 44532
rect 7708 44512 7710 44532
rect 8298 44532 8354 44568
rect 8298 44512 8300 44532
rect 8300 44512 8352 44532
rect 8352 44512 8354 44532
rect 8758 44532 8814 44568
rect 8758 44512 8760 44532
rect 8760 44512 8812 44532
rect 8812 44512 8814 44532
rect 9310 44532 9366 44568
rect 9310 44512 9312 44532
rect 9312 44512 9364 44532
rect 9364 44512 9366 44532
rect 12806 44532 12862 44568
rect 19216 44634 19272 44636
rect 19296 44634 19352 44636
rect 19376 44634 19432 44636
rect 19456 44634 19512 44636
rect 19216 44582 19262 44634
rect 19262 44582 19272 44634
rect 19296 44582 19326 44634
rect 19326 44582 19338 44634
rect 19338 44582 19352 44634
rect 19376 44582 19390 44634
rect 19390 44582 19402 44634
rect 19402 44582 19432 44634
rect 19456 44582 19466 44634
rect 19466 44582 19512 44634
rect 19216 44580 19272 44582
rect 19296 44580 19352 44582
rect 19376 44580 19432 44582
rect 19456 44580 19512 44582
rect 12806 44512 12808 44532
rect 12808 44512 12860 44532
rect 12860 44512 12862 44532
rect 4328 44090 4384 44092
rect 4408 44090 4464 44092
rect 4488 44090 4544 44092
rect 4568 44090 4624 44092
rect 4328 44038 4374 44090
rect 4374 44038 4384 44090
rect 4408 44038 4438 44090
rect 4438 44038 4450 44090
rect 4450 44038 4464 44090
rect 4488 44038 4502 44090
rect 4502 44038 4514 44090
rect 4514 44038 4544 44090
rect 4568 44038 4578 44090
rect 4578 44038 4624 44090
rect 4328 44036 4384 44038
rect 4408 44036 4464 44038
rect 4488 44036 4544 44038
rect 4568 44036 4624 44038
rect 6550 43988 6606 44024
rect 6550 43968 6552 43988
rect 6552 43968 6604 43988
rect 6604 43968 6606 43988
rect 6918 43988 6974 44024
rect 6918 43968 6920 43988
rect 6920 43968 6972 43988
rect 6972 43968 6974 43988
rect 10690 43988 10746 44024
rect 10690 43968 10692 43988
rect 10692 43968 10744 43988
rect 10744 43968 10746 43988
rect 3668 43546 3724 43548
rect 3748 43546 3804 43548
rect 3828 43546 3884 43548
rect 3908 43546 3964 43548
rect 3668 43494 3714 43546
rect 3714 43494 3724 43546
rect 3748 43494 3778 43546
rect 3778 43494 3790 43546
rect 3790 43494 3804 43546
rect 3828 43494 3842 43546
rect 3842 43494 3854 43546
rect 3854 43494 3884 43546
rect 3908 43494 3918 43546
rect 3918 43494 3964 43546
rect 3668 43492 3724 43494
rect 3748 43492 3804 43494
rect 3828 43492 3884 43494
rect 3908 43492 3964 43494
rect 4328 43002 4384 43004
rect 4408 43002 4464 43004
rect 4488 43002 4544 43004
rect 4568 43002 4624 43004
rect 4328 42950 4374 43002
rect 4374 42950 4384 43002
rect 4408 42950 4438 43002
rect 4438 42950 4450 43002
rect 4450 42950 4464 43002
rect 4488 42950 4502 43002
rect 4502 42950 4514 43002
rect 4514 42950 4544 43002
rect 4568 42950 4578 43002
rect 4578 42950 4624 43002
rect 4328 42948 4384 42950
rect 4408 42948 4464 42950
rect 4488 42948 4544 42950
rect 4568 42948 4624 42950
rect 3668 42458 3724 42460
rect 3748 42458 3804 42460
rect 3828 42458 3884 42460
rect 3908 42458 3964 42460
rect 3668 42406 3714 42458
rect 3714 42406 3724 42458
rect 3748 42406 3778 42458
rect 3778 42406 3790 42458
rect 3790 42406 3804 42458
rect 3828 42406 3842 42458
rect 3842 42406 3854 42458
rect 3854 42406 3884 42458
rect 3908 42406 3918 42458
rect 3918 42406 3964 42458
rect 3668 42404 3724 42406
rect 3748 42404 3804 42406
rect 3828 42404 3884 42406
rect 3908 42404 3964 42406
rect 4328 41914 4384 41916
rect 4408 41914 4464 41916
rect 4488 41914 4544 41916
rect 4568 41914 4624 41916
rect 4328 41862 4374 41914
rect 4374 41862 4384 41914
rect 4408 41862 4438 41914
rect 4438 41862 4450 41914
rect 4450 41862 4464 41914
rect 4488 41862 4502 41914
rect 4502 41862 4514 41914
rect 4514 41862 4544 41914
rect 4568 41862 4578 41914
rect 4578 41862 4624 41914
rect 4328 41860 4384 41862
rect 4408 41860 4464 41862
rect 4488 41860 4544 41862
rect 4568 41860 4624 41862
rect 11334 43832 11390 43888
rect 3668 41370 3724 41372
rect 3748 41370 3804 41372
rect 3828 41370 3884 41372
rect 3908 41370 3964 41372
rect 3668 41318 3714 41370
rect 3714 41318 3724 41370
rect 3748 41318 3778 41370
rect 3778 41318 3790 41370
rect 3790 41318 3804 41370
rect 3828 41318 3842 41370
rect 3842 41318 3854 41370
rect 3854 41318 3884 41370
rect 3908 41318 3918 41370
rect 3918 41318 3964 41370
rect 3668 41316 3724 41318
rect 3748 41316 3804 41318
rect 3828 41316 3884 41318
rect 3908 41316 3964 41318
rect 4328 40826 4384 40828
rect 4408 40826 4464 40828
rect 4488 40826 4544 40828
rect 4568 40826 4624 40828
rect 4328 40774 4374 40826
rect 4374 40774 4384 40826
rect 4408 40774 4438 40826
rect 4438 40774 4450 40826
rect 4450 40774 4464 40826
rect 4488 40774 4502 40826
rect 4502 40774 4514 40826
rect 4514 40774 4544 40826
rect 4568 40774 4578 40826
rect 4578 40774 4624 40826
rect 4328 40772 4384 40774
rect 4408 40772 4464 40774
rect 4488 40772 4544 40774
rect 4568 40772 4624 40774
rect 3668 40282 3724 40284
rect 3748 40282 3804 40284
rect 3828 40282 3884 40284
rect 3908 40282 3964 40284
rect 3668 40230 3714 40282
rect 3714 40230 3724 40282
rect 3748 40230 3778 40282
rect 3778 40230 3790 40282
rect 3790 40230 3804 40282
rect 3828 40230 3842 40282
rect 3842 40230 3854 40282
rect 3854 40230 3884 40282
rect 3908 40230 3918 40282
rect 3918 40230 3964 40282
rect 3668 40228 3724 40230
rect 3748 40228 3804 40230
rect 3828 40228 3884 40230
rect 3908 40228 3964 40230
rect 4328 39738 4384 39740
rect 4408 39738 4464 39740
rect 4488 39738 4544 39740
rect 4568 39738 4624 39740
rect 4328 39686 4374 39738
rect 4374 39686 4384 39738
rect 4408 39686 4438 39738
rect 4438 39686 4450 39738
rect 4450 39686 4464 39738
rect 4488 39686 4502 39738
rect 4502 39686 4514 39738
rect 4514 39686 4544 39738
rect 4568 39686 4578 39738
rect 4578 39686 4624 39738
rect 4328 39684 4384 39686
rect 4408 39684 4464 39686
rect 4488 39684 4544 39686
rect 4568 39684 4624 39686
rect 3668 39194 3724 39196
rect 3748 39194 3804 39196
rect 3828 39194 3884 39196
rect 3908 39194 3964 39196
rect 3668 39142 3714 39194
rect 3714 39142 3724 39194
rect 3748 39142 3778 39194
rect 3778 39142 3790 39194
rect 3790 39142 3804 39194
rect 3828 39142 3842 39194
rect 3842 39142 3854 39194
rect 3854 39142 3884 39194
rect 3908 39142 3918 39194
rect 3918 39142 3964 39194
rect 3668 39140 3724 39142
rect 3748 39140 3804 39142
rect 3828 39140 3884 39142
rect 3908 39140 3964 39142
rect 4328 38650 4384 38652
rect 4408 38650 4464 38652
rect 4488 38650 4544 38652
rect 4568 38650 4624 38652
rect 4328 38598 4374 38650
rect 4374 38598 4384 38650
rect 4408 38598 4438 38650
rect 4438 38598 4450 38650
rect 4450 38598 4464 38650
rect 4488 38598 4502 38650
rect 4502 38598 4514 38650
rect 4514 38598 4544 38650
rect 4568 38598 4578 38650
rect 4578 38598 4624 38650
rect 4328 38596 4384 38598
rect 4408 38596 4464 38598
rect 4488 38596 4544 38598
rect 4568 38596 4624 38598
rect 3668 38106 3724 38108
rect 3748 38106 3804 38108
rect 3828 38106 3884 38108
rect 3908 38106 3964 38108
rect 3668 38054 3714 38106
rect 3714 38054 3724 38106
rect 3748 38054 3778 38106
rect 3778 38054 3790 38106
rect 3790 38054 3804 38106
rect 3828 38054 3842 38106
rect 3842 38054 3854 38106
rect 3854 38054 3884 38106
rect 3908 38054 3918 38106
rect 3918 38054 3964 38106
rect 3668 38052 3724 38054
rect 3748 38052 3804 38054
rect 3828 38052 3884 38054
rect 3908 38052 3964 38054
rect 4328 37562 4384 37564
rect 4408 37562 4464 37564
rect 4488 37562 4544 37564
rect 4568 37562 4624 37564
rect 4328 37510 4374 37562
rect 4374 37510 4384 37562
rect 4408 37510 4438 37562
rect 4438 37510 4450 37562
rect 4450 37510 4464 37562
rect 4488 37510 4502 37562
rect 4502 37510 4514 37562
rect 4514 37510 4544 37562
rect 4568 37510 4578 37562
rect 4578 37510 4624 37562
rect 4328 37508 4384 37510
rect 4408 37508 4464 37510
rect 4488 37508 4544 37510
rect 4568 37508 4624 37510
rect 3668 37018 3724 37020
rect 3748 37018 3804 37020
rect 3828 37018 3884 37020
rect 3908 37018 3964 37020
rect 3668 36966 3714 37018
rect 3714 36966 3724 37018
rect 3748 36966 3778 37018
rect 3778 36966 3790 37018
rect 3790 36966 3804 37018
rect 3828 36966 3842 37018
rect 3842 36966 3854 37018
rect 3854 36966 3884 37018
rect 3908 36966 3918 37018
rect 3918 36966 3964 37018
rect 3668 36964 3724 36966
rect 3748 36964 3804 36966
rect 3828 36964 3884 36966
rect 3908 36964 3964 36966
rect 4328 36474 4384 36476
rect 4408 36474 4464 36476
rect 4488 36474 4544 36476
rect 4568 36474 4624 36476
rect 4328 36422 4374 36474
rect 4374 36422 4384 36474
rect 4408 36422 4438 36474
rect 4438 36422 4450 36474
rect 4450 36422 4464 36474
rect 4488 36422 4502 36474
rect 4502 36422 4514 36474
rect 4514 36422 4544 36474
rect 4568 36422 4578 36474
rect 4578 36422 4624 36474
rect 4328 36420 4384 36422
rect 4408 36420 4464 36422
rect 4488 36420 4544 36422
rect 4568 36420 4624 36422
rect 3668 35930 3724 35932
rect 3748 35930 3804 35932
rect 3828 35930 3884 35932
rect 3908 35930 3964 35932
rect 3668 35878 3714 35930
rect 3714 35878 3724 35930
rect 3748 35878 3778 35930
rect 3778 35878 3790 35930
rect 3790 35878 3804 35930
rect 3828 35878 3842 35930
rect 3842 35878 3854 35930
rect 3854 35878 3884 35930
rect 3908 35878 3918 35930
rect 3918 35878 3964 35930
rect 3668 35876 3724 35878
rect 3748 35876 3804 35878
rect 3828 35876 3884 35878
rect 3908 35876 3964 35878
rect 4328 35386 4384 35388
rect 4408 35386 4464 35388
rect 4488 35386 4544 35388
rect 4568 35386 4624 35388
rect 4328 35334 4374 35386
rect 4374 35334 4384 35386
rect 4408 35334 4438 35386
rect 4438 35334 4450 35386
rect 4450 35334 4464 35386
rect 4488 35334 4502 35386
rect 4502 35334 4514 35386
rect 4514 35334 4544 35386
rect 4568 35334 4578 35386
rect 4578 35334 4624 35386
rect 4328 35332 4384 35334
rect 4408 35332 4464 35334
rect 4488 35332 4544 35334
rect 4568 35332 4624 35334
rect 3668 34842 3724 34844
rect 3748 34842 3804 34844
rect 3828 34842 3884 34844
rect 3908 34842 3964 34844
rect 3668 34790 3714 34842
rect 3714 34790 3724 34842
rect 3748 34790 3778 34842
rect 3778 34790 3790 34842
rect 3790 34790 3804 34842
rect 3828 34790 3842 34842
rect 3842 34790 3854 34842
rect 3854 34790 3884 34842
rect 3908 34790 3918 34842
rect 3918 34790 3964 34842
rect 3668 34788 3724 34790
rect 3748 34788 3804 34790
rect 3828 34788 3884 34790
rect 3908 34788 3964 34790
rect 4328 34298 4384 34300
rect 4408 34298 4464 34300
rect 4488 34298 4544 34300
rect 4568 34298 4624 34300
rect 4328 34246 4374 34298
rect 4374 34246 4384 34298
rect 4408 34246 4438 34298
rect 4438 34246 4450 34298
rect 4450 34246 4464 34298
rect 4488 34246 4502 34298
rect 4502 34246 4514 34298
rect 4514 34246 4544 34298
rect 4568 34246 4578 34298
rect 4578 34246 4624 34298
rect 4328 34244 4384 34246
rect 4408 34244 4464 34246
rect 4488 34244 4544 34246
rect 4568 34244 4624 34246
rect 3668 33754 3724 33756
rect 3748 33754 3804 33756
rect 3828 33754 3884 33756
rect 3908 33754 3964 33756
rect 3668 33702 3714 33754
rect 3714 33702 3724 33754
rect 3748 33702 3778 33754
rect 3778 33702 3790 33754
rect 3790 33702 3804 33754
rect 3828 33702 3842 33754
rect 3842 33702 3854 33754
rect 3854 33702 3884 33754
rect 3908 33702 3918 33754
rect 3918 33702 3964 33754
rect 3668 33700 3724 33702
rect 3748 33700 3804 33702
rect 3828 33700 3884 33702
rect 3908 33700 3964 33702
rect 4328 33210 4384 33212
rect 4408 33210 4464 33212
rect 4488 33210 4544 33212
rect 4568 33210 4624 33212
rect 4328 33158 4374 33210
rect 4374 33158 4384 33210
rect 4408 33158 4438 33210
rect 4438 33158 4450 33210
rect 4450 33158 4464 33210
rect 4488 33158 4502 33210
rect 4502 33158 4514 33210
rect 4514 33158 4544 33210
rect 4568 33158 4578 33210
rect 4578 33158 4624 33210
rect 4328 33156 4384 33158
rect 4408 33156 4464 33158
rect 4488 33156 4544 33158
rect 4568 33156 4624 33158
rect 3668 32666 3724 32668
rect 3748 32666 3804 32668
rect 3828 32666 3884 32668
rect 3908 32666 3964 32668
rect 3668 32614 3714 32666
rect 3714 32614 3724 32666
rect 3748 32614 3778 32666
rect 3778 32614 3790 32666
rect 3790 32614 3804 32666
rect 3828 32614 3842 32666
rect 3842 32614 3854 32666
rect 3854 32614 3884 32666
rect 3908 32614 3918 32666
rect 3918 32614 3964 32666
rect 3668 32612 3724 32614
rect 3748 32612 3804 32614
rect 3828 32612 3884 32614
rect 3908 32612 3964 32614
rect 4328 32122 4384 32124
rect 4408 32122 4464 32124
rect 4488 32122 4544 32124
rect 4568 32122 4624 32124
rect 4328 32070 4374 32122
rect 4374 32070 4384 32122
rect 4408 32070 4438 32122
rect 4438 32070 4450 32122
rect 4450 32070 4464 32122
rect 4488 32070 4502 32122
rect 4502 32070 4514 32122
rect 4514 32070 4544 32122
rect 4568 32070 4578 32122
rect 4578 32070 4624 32122
rect 4328 32068 4384 32070
rect 4408 32068 4464 32070
rect 4488 32068 4544 32070
rect 4568 32068 4624 32070
rect 3668 31578 3724 31580
rect 3748 31578 3804 31580
rect 3828 31578 3884 31580
rect 3908 31578 3964 31580
rect 3668 31526 3714 31578
rect 3714 31526 3724 31578
rect 3748 31526 3778 31578
rect 3778 31526 3790 31578
rect 3790 31526 3804 31578
rect 3828 31526 3842 31578
rect 3842 31526 3854 31578
rect 3854 31526 3884 31578
rect 3908 31526 3918 31578
rect 3918 31526 3964 31578
rect 3668 31524 3724 31526
rect 3748 31524 3804 31526
rect 3828 31524 3884 31526
rect 3908 31524 3964 31526
rect 4328 31034 4384 31036
rect 4408 31034 4464 31036
rect 4488 31034 4544 31036
rect 4568 31034 4624 31036
rect 4328 30982 4374 31034
rect 4374 30982 4384 31034
rect 4408 30982 4438 31034
rect 4438 30982 4450 31034
rect 4450 30982 4464 31034
rect 4488 30982 4502 31034
rect 4502 30982 4514 31034
rect 4514 30982 4544 31034
rect 4568 30982 4578 31034
rect 4578 30982 4624 31034
rect 4328 30980 4384 30982
rect 4408 30980 4464 30982
rect 4488 30980 4544 30982
rect 4568 30980 4624 30982
rect 3668 30490 3724 30492
rect 3748 30490 3804 30492
rect 3828 30490 3884 30492
rect 3908 30490 3964 30492
rect 3668 30438 3714 30490
rect 3714 30438 3724 30490
rect 3748 30438 3778 30490
rect 3778 30438 3790 30490
rect 3790 30438 3804 30490
rect 3828 30438 3842 30490
rect 3842 30438 3854 30490
rect 3854 30438 3884 30490
rect 3908 30438 3918 30490
rect 3918 30438 3964 30490
rect 3668 30436 3724 30438
rect 3748 30436 3804 30438
rect 3828 30436 3884 30438
rect 3908 30436 3964 30438
rect 11442 43546 11498 43548
rect 11522 43546 11578 43548
rect 11602 43546 11658 43548
rect 11682 43546 11738 43548
rect 11442 43494 11488 43546
rect 11488 43494 11498 43546
rect 11522 43494 11552 43546
rect 11552 43494 11564 43546
rect 11564 43494 11578 43546
rect 11602 43494 11616 43546
rect 11616 43494 11628 43546
rect 11628 43494 11658 43546
rect 11682 43494 11692 43546
rect 11692 43494 11738 43546
rect 11442 43492 11498 43494
rect 11522 43492 11578 43494
rect 11602 43492 11658 43494
rect 11682 43492 11738 43494
rect 24030 44648 24086 44704
rect 24398 44648 24454 44704
rect 24950 44648 25006 44704
rect 25502 44648 25558 44704
rect 26054 44648 26110 44704
rect 26514 44648 26570 44704
rect 12102 44090 12158 44092
rect 12182 44090 12238 44092
rect 12262 44090 12318 44092
rect 12342 44090 12398 44092
rect 12102 44038 12148 44090
rect 12148 44038 12158 44090
rect 12182 44038 12212 44090
rect 12212 44038 12224 44090
rect 12224 44038 12238 44090
rect 12262 44038 12276 44090
rect 12276 44038 12288 44090
rect 12288 44038 12318 44090
rect 12342 44038 12352 44090
rect 12352 44038 12398 44090
rect 12102 44036 12158 44038
rect 12182 44036 12238 44038
rect 12262 44036 12318 44038
rect 12342 44036 12398 44038
rect 10966 39888 11022 39944
rect 11442 42458 11498 42460
rect 11522 42458 11578 42460
rect 11602 42458 11658 42460
rect 11682 42458 11738 42460
rect 11442 42406 11488 42458
rect 11488 42406 11498 42458
rect 11522 42406 11552 42458
rect 11552 42406 11564 42458
rect 11564 42406 11578 42458
rect 11602 42406 11616 42458
rect 11616 42406 11628 42458
rect 11628 42406 11658 42458
rect 11682 42406 11692 42458
rect 11692 42406 11738 42458
rect 11442 42404 11498 42406
rect 11522 42404 11578 42406
rect 11602 42404 11658 42406
rect 11682 42404 11738 42406
rect 11442 41370 11498 41372
rect 11522 41370 11578 41372
rect 11602 41370 11658 41372
rect 11682 41370 11738 41372
rect 11442 41318 11488 41370
rect 11488 41318 11498 41370
rect 11522 41318 11552 41370
rect 11552 41318 11564 41370
rect 11564 41318 11578 41370
rect 11602 41318 11616 41370
rect 11616 41318 11628 41370
rect 11628 41318 11658 41370
rect 11682 41318 11692 41370
rect 11692 41318 11738 41370
rect 11442 41316 11498 41318
rect 11522 41316 11578 41318
rect 11602 41316 11658 41318
rect 11682 41316 11738 41318
rect 11442 40282 11498 40284
rect 11522 40282 11578 40284
rect 11602 40282 11658 40284
rect 11682 40282 11738 40284
rect 11442 40230 11488 40282
rect 11488 40230 11498 40282
rect 11522 40230 11552 40282
rect 11552 40230 11564 40282
rect 11564 40230 11578 40282
rect 11602 40230 11616 40282
rect 11616 40230 11628 40282
rect 11628 40230 11658 40282
rect 11682 40230 11692 40282
rect 11692 40230 11738 40282
rect 11442 40228 11498 40230
rect 11522 40228 11578 40230
rect 11602 40228 11658 40230
rect 11682 40228 11738 40230
rect 12102 43002 12158 43004
rect 12182 43002 12238 43004
rect 12262 43002 12318 43004
rect 12342 43002 12398 43004
rect 12102 42950 12148 43002
rect 12148 42950 12158 43002
rect 12182 42950 12212 43002
rect 12212 42950 12224 43002
rect 12224 42950 12238 43002
rect 12262 42950 12276 43002
rect 12276 42950 12288 43002
rect 12288 42950 12318 43002
rect 12342 42950 12352 43002
rect 12352 42950 12398 43002
rect 12102 42948 12158 42950
rect 12182 42948 12238 42950
rect 12262 42948 12318 42950
rect 12342 42948 12398 42950
rect 13266 43988 13322 44024
rect 13266 43968 13268 43988
rect 13268 43968 13320 43988
rect 13320 43968 13322 43988
rect 13818 43696 13874 43752
rect 14370 43444 14426 43480
rect 14370 43424 14372 43444
rect 14372 43424 14424 43444
rect 14424 43424 14426 43444
rect 12102 41914 12158 41916
rect 12182 41914 12238 41916
rect 12262 41914 12318 41916
rect 12342 41914 12398 41916
rect 12102 41862 12148 41914
rect 12148 41862 12158 41914
rect 12182 41862 12212 41914
rect 12212 41862 12224 41914
rect 12224 41862 12238 41914
rect 12262 41862 12276 41914
rect 12276 41862 12288 41914
rect 12288 41862 12318 41914
rect 12342 41862 12352 41914
rect 12352 41862 12398 41914
rect 12102 41860 12158 41862
rect 12182 41860 12238 41862
rect 12262 41860 12318 41862
rect 12342 41860 12398 41862
rect 13726 41792 13782 41848
rect 12102 40826 12158 40828
rect 12182 40826 12238 40828
rect 12262 40826 12318 40828
rect 12342 40826 12398 40828
rect 12102 40774 12148 40826
rect 12148 40774 12158 40826
rect 12182 40774 12212 40826
rect 12212 40774 12224 40826
rect 12224 40774 12238 40826
rect 12262 40774 12276 40826
rect 12276 40774 12288 40826
rect 12288 40774 12318 40826
rect 12342 40774 12352 40826
rect 12352 40774 12398 40826
rect 12102 40772 12158 40774
rect 12182 40772 12238 40774
rect 12262 40772 12318 40774
rect 12342 40772 12398 40774
rect 11442 39194 11498 39196
rect 11522 39194 11578 39196
rect 11602 39194 11658 39196
rect 11682 39194 11738 39196
rect 11442 39142 11488 39194
rect 11488 39142 11498 39194
rect 11522 39142 11552 39194
rect 11552 39142 11564 39194
rect 11564 39142 11578 39194
rect 11602 39142 11616 39194
rect 11616 39142 11628 39194
rect 11628 39142 11658 39194
rect 11682 39142 11692 39194
rect 11692 39142 11738 39194
rect 11442 39140 11498 39142
rect 11522 39140 11578 39142
rect 11602 39140 11658 39142
rect 11682 39140 11738 39142
rect 11442 38106 11498 38108
rect 11522 38106 11578 38108
rect 11602 38106 11658 38108
rect 11682 38106 11738 38108
rect 11442 38054 11488 38106
rect 11488 38054 11498 38106
rect 11522 38054 11552 38106
rect 11552 38054 11564 38106
rect 11564 38054 11578 38106
rect 11602 38054 11616 38106
rect 11616 38054 11628 38106
rect 11628 38054 11658 38106
rect 11682 38054 11692 38106
rect 11692 38054 11738 38106
rect 11442 38052 11498 38054
rect 11522 38052 11578 38054
rect 11602 38052 11658 38054
rect 11682 38052 11738 38054
rect 11442 37018 11498 37020
rect 11522 37018 11578 37020
rect 11602 37018 11658 37020
rect 11682 37018 11738 37020
rect 11442 36966 11488 37018
rect 11488 36966 11498 37018
rect 11522 36966 11552 37018
rect 11552 36966 11564 37018
rect 11564 36966 11578 37018
rect 11602 36966 11616 37018
rect 11616 36966 11628 37018
rect 11628 36966 11658 37018
rect 11682 36966 11692 37018
rect 11692 36966 11738 37018
rect 11442 36964 11498 36966
rect 11522 36964 11578 36966
rect 11602 36964 11658 36966
rect 11682 36964 11738 36966
rect 11442 35930 11498 35932
rect 11522 35930 11578 35932
rect 11602 35930 11658 35932
rect 11682 35930 11738 35932
rect 11442 35878 11488 35930
rect 11488 35878 11498 35930
rect 11522 35878 11552 35930
rect 11552 35878 11564 35930
rect 11564 35878 11578 35930
rect 11602 35878 11616 35930
rect 11616 35878 11628 35930
rect 11628 35878 11658 35930
rect 11682 35878 11692 35930
rect 11692 35878 11738 35930
rect 11442 35876 11498 35878
rect 11522 35876 11578 35878
rect 11602 35876 11658 35878
rect 11682 35876 11738 35878
rect 12102 39738 12158 39740
rect 12182 39738 12238 39740
rect 12262 39738 12318 39740
rect 12342 39738 12398 39740
rect 12102 39686 12148 39738
rect 12148 39686 12158 39738
rect 12182 39686 12212 39738
rect 12212 39686 12224 39738
rect 12224 39686 12238 39738
rect 12262 39686 12276 39738
rect 12276 39686 12288 39738
rect 12288 39686 12318 39738
rect 12342 39686 12352 39738
rect 12352 39686 12398 39738
rect 12102 39684 12158 39686
rect 12182 39684 12238 39686
rect 12262 39684 12318 39686
rect 12342 39684 12398 39686
rect 12102 38650 12158 38652
rect 12182 38650 12238 38652
rect 12262 38650 12318 38652
rect 12342 38650 12398 38652
rect 12102 38598 12148 38650
rect 12148 38598 12158 38650
rect 12182 38598 12212 38650
rect 12212 38598 12224 38650
rect 12224 38598 12238 38650
rect 12262 38598 12276 38650
rect 12276 38598 12288 38650
rect 12288 38598 12318 38650
rect 12342 38598 12352 38650
rect 12352 38598 12398 38650
rect 12102 38596 12158 38598
rect 12182 38596 12238 38598
rect 12262 38596 12318 38598
rect 12342 38596 12398 38598
rect 12102 37562 12158 37564
rect 12182 37562 12238 37564
rect 12262 37562 12318 37564
rect 12342 37562 12398 37564
rect 12102 37510 12148 37562
rect 12148 37510 12158 37562
rect 12182 37510 12212 37562
rect 12212 37510 12224 37562
rect 12224 37510 12238 37562
rect 12262 37510 12276 37562
rect 12276 37510 12288 37562
rect 12288 37510 12318 37562
rect 12342 37510 12352 37562
rect 12352 37510 12398 37562
rect 12102 37508 12158 37510
rect 12182 37508 12238 37510
rect 12262 37508 12318 37510
rect 12342 37508 12398 37510
rect 12990 39888 13046 39944
rect 12102 36474 12158 36476
rect 12182 36474 12238 36476
rect 12262 36474 12318 36476
rect 12342 36474 12398 36476
rect 12102 36422 12148 36474
rect 12148 36422 12158 36474
rect 12182 36422 12212 36474
rect 12212 36422 12224 36474
rect 12224 36422 12238 36474
rect 12262 36422 12276 36474
rect 12276 36422 12288 36474
rect 12288 36422 12318 36474
rect 12342 36422 12352 36474
rect 12352 36422 12398 36474
rect 12102 36420 12158 36422
rect 12182 36420 12238 36422
rect 12262 36420 12318 36422
rect 12342 36420 12398 36422
rect 12102 35386 12158 35388
rect 12182 35386 12238 35388
rect 12262 35386 12318 35388
rect 12342 35386 12398 35388
rect 12102 35334 12148 35386
rect 12148 35334 12158 35386
rect 12182 35334 12212 35386
rect 12212 35334 12224 35386
rect 12224 35334 12238 35386
rect 12262 35334 12276 35386
rect 12276 35334 12288 35386
rect 12288 35334 12318 35386
rect 12342 35334 12352 35386
rect 12352 35334 12398 35386
rect 12102 35332 12158 35334
rect 12182 35332 12238 35334
rect 12262 35332 12318 35334
rect 12342 35332 12398 35334
rect 11442 34842 11498 34844
rect 11522 34842 11578 34844
rect 11602 34842 11658 34844
rect 11682 34842 11738 34844
rect 11442 34790 11488 34842
rect 11488 34790 11498 34842
rect 11522 34790 11552 34842
rect 11552 34790 11564 34842
rect 11564 34790 11578 34842
rect 11602 34790 11616 34842
rect 11616 34790 11628 34842
rect 11628 34790 11658 34842
rect 11682 34790 11692 34842
rect 11692 34790 11738 34842
rect 11442 34788 11498 34790
rect 11522 34788 11578 34790
rect 11602 34788 11658 34790
rect 11682 34788 11738 34790
rect 11442 33754 11498 33756
rect 11522 33754 11578 33756
rect 11602 33754 11658 33756
rect 11682 33754 11738 33756
rect 11442 33702 11488 33754
rect 11488 33702 11498 33754
rect 11522 33702 11552 33754
rect 11552 33702 11564 33754
rect 11564 33702 11578 33754
rect 11602 33702 11616 33754
rect 11616 33702 11628 33754
rect 11628 33702 11658 33754
rect 11682 33702 11692 33754
rect 11692 33702 11738 33754
rect 11442 33700 11498 33702
rect 11522 33700 11578 33702
rect 11602 33700 11658 33702
rect 11682 33700 11738 33702
rect 11610 33380 11666 33416
rect 11610 33360 11612 33380
rect 11612 33360 11664 33380
rect 11664 33360 11666 33380
rect 11442 32666 11498 32668
rect 11522 32666 11578 32668
rect 11602 32666 11658 32668
rect 11682 32666 11738 32668
rect 11442 32614 11488 32666
rect 11488 32614 11498 32666
rect 11522 32614 11552 32666
rect 11552 32614 11564 32666
rect 11564 32614 11578 32666
rect 11602 32614 11616 32666
rect 11616 32614 11628 32666
rect 11628 32614 11658 32666
rect 11682 32614 11692 32666
rect 11692 32614 11738 32666
rect 11442 32612 11498 32614
rect 11522 32612 11578 32614
rect 11602 32612 11658 32614
rect 11682 32612 11738 32614
rect 11442 31578 11498 31580
rect 11522 31578 11578 31580
rect 11602 31578 11658 31580
rect 11682 31578 11738 31580
rect 11442 31526 11488 31578
rect 11488 31526 11498 31578
rect 11522 31526 11552 31578
rect 11552 31526 11564 31578
rect 11564 31526 11578 31578
rect 11602 31526 11616 31578
rect 11616 31526 11628 31578
rect 11628 31526 11658 31578
rect 11682 31526 11692 31578
rect 11692 31526 11738 31578
rect 11442 31524 11498 31526
rect 11522 31524 11578 31526
rect 11602 31524 11658 31526
rect 11682 31524 11738 31526
rect 11442 30490 11498 30492
rect 11522 30490 11578 30492
rect 11602 30490 11658 30492
rect 11682 30490 11738 30492
rect 11442 30438 11488 30490
rect 11488 30438 11498 30490
rect 11522 30438 11552 30490
rect 11552 30438 11564 30490
rect 11564 30438 11578 30490
rect 11602 30438 11616 30490
rect 11616 30438 11628 30490
rect 11628 30438 11658 30490
rect 11682 30438 11692 30490
rect 11692 30438 11738 30490
rect 11442 30436 11498 30438
rect 11522 30436 11578 30438
rect 11602 30436 11658 30438
rect 11682 30436 11738 30438
rect 12714 35028 12716 35048
rect 12716 35028 12768 35048
rect 12768 35028 12770 35048
rect 12714 34992 12770 35028
rect 12102 34298 12158 34300
rect 12182 34298 12238 34300
rect 12262 34298 12318 34300
rect 12342 34298 12398 34300
rect 12102 34246 12148 34298
rect 12148 34246 12158 34298
rect 12182 34246 12212 34298
rect 12212 34246 12224 34298
rect 12224 34246 12238 34298
rect 12262 34246 12276 34298
rect 12276 34246 12288 34298
rect 12288 34246 12318 34298
rect 12342 34246 12352 34298
rect 12352 34246 12398 34298
rect 12102 34244 12158 34246
rect 12182 34244 12238 34246
rect 12262 34244 12318 34246
rect 12342 34244 12398 34246
rect 12530 33396 12532 33416
rect 12532 33396 12584 33416
rect 12584 33396 12586 33416
rect 12530 33360 12586 33396
rect 12102 33210 12158 33212
rect 12182 33210 12238 33212
rect 12262 33210 12318 33212
rect 12342 33210 12398 33212
rect 12102 33158 12148 33210
rect 12148 33158 12158 33210
rect 12182 33158 12212 33210
rect 12212 33158 12224 33210
rect 12224 33158 12238 33210
rect 12262 33158 12276 33210
rect 12276 33158 12288 33210
rect 12288 33158 12318 33210
rect 12342 33158 12352 33210
rect 12352 33158 12398 33210
rect 12102 33156 12158 33158
rect 12182 33156 12238 33158
rect 12262 33156 12318 33158
rect 12342 33156 12398 33158
rect 13726 34992 13782 35048
rect 12102 32122 12158 32124
rect 12182 32122 12238 32124
rect 12262 32122 12318 32124
rect 12342 32122 12398 32124
rect 12102 32070 12148 32122
rect 12148 32070 12158 32122
rect 12182 32070 12212 32122
rect 12212 32070 12224 32122
rect 12224 32070 12238 32122
rect 12262 32070 12276 32122
rect 12276 32070 12288 32122
rect 12288 32070 12318 32122
rect 12342 32070 12352 32122
rect 12352 32070 12398 32122
rect 12102 32068 12158 32070
rect 12182 32068 12238 32070
rect 12262 32068 12318 32070
rect 12342 32068 12398 32070
rect 14278 35944 14334 36000
rect 12102 31034 12158 31036
rect 12182 31034 12238 31036
rect 12262 31034 12318 31036
rect 12342 31034 12398 31036
rect 12102 30982 12148 31034
rect 12148 30982 12158 31034
rect 12182 30982 12212 31034
rect 12212 30982 12224 31034
rect 12224 30982 12238 31034
rect 12262 30982 12276 31034
rect 12276 30982 12288 31034
rect 12288 30982 12318 31034
rect 12342 30982 12352 31034
rect 12352 30982 12398 31034
rect 12102 30980 12158 30982
rect 12182 30980 12238 30982
rect 12262 30980 12318 30982
rect 12342 30980 12398 30982
rect 4328 29946 4384 29948
rect 4408 29946 4464 29948
rect 4488 29946 4544 29948
rect 4568 29946 4624 29948
rect 4328 29894 4374 29946
rect 4374 29894 4384 29946
rect 4408 29894 4438 29946
rect 4438 29894 4450 29946
rect 4450 29894 4464 29946
rect 4488 29894 4502 29946
rect 4502 29894 4514 29946
rect 4514 29894 4544 29946
rect 4568 29894 4578 29946
rect 4578 29894 4624 29946
rect 4328 29892 4384 29894
rect 4408 29892 4464 29894
rect 4488 29892 4544 29894
rect 4568 29892 4624 29894
rect 3668 29402 3724 29404
rect 3748 29402 3804 29404
rect 3828 29402 3884 29404
rect 3908 29402 3964 29404
rect 3668 29350 3714 29402
rect 3714 29350 3724 29402
rect 3748 29350 3778 29402
rect 3778 29350 3790 29402
rect 3790 29350 3804 29402
rect 3828 29350 3842 29402
rect 3842 29350 3854 29402
rect 3854 29350 3884 29402
rect 3908 29350 3918 29402
rect 3918 29350 3964 29402
rect 3668 29348 3724 29350
rect 3748 29348 3804 29350
rect 3828 29348 3884 29350
rect 3908 29348 3964 29350
rect 11442 29402 11498 29404
rect 11522 29402 11578 29404
rect 11602 29402 11658 29404
rect 11682 29402 11738 29404
rect 11442 29350 11488 29402
rect 11488 29350 11498 29402
rect 11522 29350 11552 29402
rect 11552 29350 11564 29402
rect 11564 29350 11578 29402
rect 11602 29350 11616 29402
rect 11616 29350 11628 29402
rect 11628 29350 11658 29402
rect 11682 29350 11692 29402
rect 11692 29350 11738 29402
rect 11442 29348 11498 29350
rect 11522 29348 11578 29350
rect 11602 29348 11658 29350
rect 11682 29348 11738 29350
rect 4328 28858 4384 28860
rect 4408 28858 4464 28860
rect 4488 28858 4544 28860
rect 4568 28858 4624 28860
rect 4328 28806 4374 28858
rect 4374 28806 4384 28858
rect 4408 28806 4438 28858
rect 4438 28806 4450 28858
rect 4450 28806 4464 28858
rect 4488 28806 4502 28858
rect 4502 28806 4514 28858
rect 4514 28806 4544 28858
rect 4568 28806 4578 28858
rect 4578 28806 4624 28858
rect 4328 28804 4384 28806
rect 4408 28804 4464 28806
rect 4488 28804 4544 28806
rect 4568 28804 4624 28806
rect 3668 28314 3724 28316
rect 3748 28314 3804 28316
rect 3828 28314 3884 28316
rect 3908 28314 3964 28316
rect 3668 28262 3714 28314
rect 3714 28262 3724 28314
rect 3748 28262 3778 28314
rect 3778 28262 3790 28314
rect 3790 28262 3804 28314
rect 3828 28262 3842 28314
rect 3842 28262 3854 28314
rect 3854 28262 3884 28314
rect 3908 28262 3918 28314
rect 3918 28262 3964 28314
rect 3668 28260 3724 28262
rect 3748 28260 3804 28262
rect 3828 28260 3884 28262
rect 3908 28260 3964 28262
rect 12102 29946 12158 29948
rect 12182 29946 12238 29948
rect 12262 29946 12318 29948
rect 12342 29946 12398 29948
rect 12102 29894 12148 29946
rect 12148 29894 12158 29946
rect 12182 29894 12212 29946
rect 12212 29894 12224 29946
rect 12224 29894 12238 29946
rect 12262 29894 12276 29946
rect 12276 29894 12288 29946
rect 12288 29894 12318 29946
rect 12342 29894 12352 29946
rect 12352 29894 12398 29946
rect 12102 29892 12158 29894
rect 12182 29892 12238 29894
rect 12262 29892 12318 29894
rect 12342 29892 12398 29894
rect 12102 28858 12158 28860
rect 12182 28858 12238 28860
rect 12262 28858 12318 28860
rect 12342 28858 12398 28860
rect 12102 28806 12148 28858
rect 12148 28806 12158 28858
rect 12182 28806 12212 28858
rect 12212 28806 12224 28858
rect 12224 28806 12238 28858
rect 12262 28806 12276 28858
rect 12276 28806 12288 28858
rect 12288 28806 12318 28858
rect 12342 28806 12352 28858
rect 12352 28806 12398 28858
rect 12102 28804 12158 28806
rect 12182 28804 12238 28806
rect 12262 28804 12318 28806
rect 12342 28804 12398 28806
rect 11442 28314 11498 28316
rect 11522 28314 11578 28316
rect 11602 28314 11658 28316
rect 11682 28314 11738 28316
rect 11442 28262 11488 28314
rect 11488 28262 11498 28314
rect 11522 28262 11552 28314
rect 11552 28262 11564 28314
rect 11564 28262 11578 28314
rect 11602 28262 11616 28314
rect 11616 28262 11628 28314
rect 11628 28262 11658 28314
rect 11682 28262 11692 28314
rect 11692 28262 11738 28314
rect 11442 28260 11498 28262
rect 11522 28260 11578 28262
rect 11602 28260 11658 28262
rect 11682 28260 11738 28262
rect 4328 27770 4384 27772
rect 4408 27770 4464 27772
rect 4488 27770 4544 27772
rect 4568 27770 4624 27772
rect 4328 27718 4374 27770
rect 4374 27718 4384 27770
rect 4408 27718 4438 27770
rect 4438 27718 4450 27770
rect 4450 27718 4464 27770
rect 4488 27718 4502 27770
rect 4502 27718 4514 27770
rect 4514 27718 4544 27770
rect 4568 27718 4578 27770
rect 4578 27718 4624 27770
rect 4328 27716 4384 27718
rect 4408 27716 4464 27718
rect 4488 27716 4544 27718
rect 4568 27716 4624 27718
rect 12102 27770 12158 27772
rect 12182 27770 12238 27772
rect 12262 27770 12318 27772
rect 12342 27770 12398 27772
rect 12102 27718 12148 27770
rect 12148 27718 12158 27770
rect 12182 27718 12212 27770
rect 12212 27718 12224 27770
rect 12224 27718 12238 27770
rect 12262 27718 12276 27770
rect 12276 27718 12288 27770
rect 12288 27718 12318 27770
rect 12342 27718 12352 27770
rect 12352 27718 12398 27770
rect 12102 27716 12158 27718
rect 12182 27716 12238 27718
rect 12262 27716 12318 27718
rect 12342 27716 12398 27718
rect 3668 27226 3724 27228
rect 3748 27226 3804 27228
rect 3828 27226 3884 27228
rect 3908 27226 3964 27228
rect 3668 27174 3714 27226
rect 3714 27174 3724 27226
rect 3748 27174 3778 27226
rect 3778 27174 3790 27226
rect 3790 27174 3804 27226
rect 3828 27174 3842 27226
rect 3842 27174 3854 27226
rect 3854 27174 3884 27226
rect 3908 27174 3918 27226
rect 3918 27174 3964 27226
rect 3668 27172 3724 27174
rect 3748 27172 3804 27174
rect 3828 27172 3884 27174
rect 3908 27172 3964 27174
rect 11442 27226 11498 27228
rect 11522 27226 11578 27228
rect 11602 27226 11658 27228
rect 11682 27226 11738 27228
rect 11442 27174 11488 27226
rect 11488 27174 11498 27226
rect 11522 27174 11552 27226
rect 11552 27174 11564 27226
rect 11564 27174 11578 27226
rect 11602 27174 11616 27226
rect 11616 27174 11628 27226
rect 11628 27174 11658 27226
rect 11682 27174 11692 27226
rect 11692 27174 11738 27226
rect 11442 27172 11498 27174
rect 11522 27172 11578 27174
rect 11602 27172 11658 27174
rect 11682 27172 11738 27174
rect 15106 43152 15162 43208
rect 14278 28756 14334 28792
rect 14278 28736 14280 28756
rect 14280 28736 14332 28756
rect 14332 28736 14334 28756
rect 4328 26682 4384 26684
rect 4408 26682 4464 26684
rect 4488 26682 4544 26684
rect 4568 26682 4624 26684
rect 4328 26630 4374 26682
rect 4374 26630 4384 26682
rect 4408 26630 4438 26682
rect 4438 26630 4450 26682
rect 4450 26630 4464 26682
rect 4488 26630 4502 26682
rect 4502 26630 4514 26682
rect 4514 26630 4544 26682
rect 4568 26630 4578 26682
rect 4578 26630 4624 26682
rect 4328 26628 4384 26630
rect 4408 26628 4464 26630
rect 4488 26628 4544 26630
rect 4568 26628 4624 26630
rect 3668 26138 3724 26140
rect 3748 26138 3804 26140
rect 3828 26138 3884 26140
rect 3908 26138 3964 26140
rect 3668 26086 3714 26138
rect 3714 26086 3724 26138
rect 3748 26086 3778 26138
rect 3778 26086 3790 26138
rect 3790 26086 3804 26138
rect 3828 26086 3842 26138
rect 3842 26086 3854 26138
rect 3854 26086 3884 26138
rect 3908 26086 3918 26138
rect 3918 26086 3964 26138
rect 3668 26084 3724 26086
rect 3748 26084 3804 26086
rect 3828 26084 3884 26086
rect 3908 26084 3964 26086
rect 12102 26682 12158 26684
rect 12182 26682 12238 26684
rect 12262 26682 12318 26684
rect 12342 26682 12398 26684
rect 12102 26630 12148 26682
rect 12148 26630 12158 26682
rect 12182 26630 12212 26682
rect 12212 26630 12224 26682
rect 12224 26630 12238 26682
rect 12262 26630 12276 26682
rect 12276 26630 12288 26682
rect 12288 26630 12318 26682
rect 12342 26630 12352 26682
rect 12352 26630 12398 26682
rect 12102 26628 12158 26630
rect 12182 26628 12238 26630
rect 12262 26628 12318 26630
rect 12342 26628 12398 26630
rect 15474 42900 15530 42936
rect 15474 42880 15476 42900
rect 15476 42880 15528 42900
rect 15528 42880 15530 42900
rect 16578 43968 16634 44024
rect 17406 43968 17462 44024
rect 18142 43988 18198 44024
rect 18142 43968 18144 43988
rect 18144 43968 18196 43988
rect 18196 43968 18198 43988
rect 16302 41112 16358 41168
rect 19876 44090 19932 44092
rect 19956 44090 20012 44092
rect 20036 44090 20092 44092
rect 20116 44090 20172 44092
rect 19876 44038 19922 44090
rect 19922 44038 19932 44090
rect 19956 44038 19986 44090
rect 19986 44038 19998 44090
rect 19998 44038 20012 44090
rect 20036 44038 20050 44090
rect 20050 44038 20062 44090
rect 20062 44038 20092 44090
rect 20116 44038 20126 44090
rect 20126 44038 20172 44090
rect 19876 44036 19932 44038
rect 19956 44036 20012 44038
rect 20036 44036 20092 44038
rect 20116 44036 20172 44038
rect 19216 43546 19272 43548
rect 19296 43546 19352 43548
rect 19376 43546 19432 43548
rect 19456 43546 19512 43548
rect 19216 43494 19262 43546
rect 19262 43494 19272 43546
rect 19296 43494 19326 43546
rect 19326 43494 19338 43546
rect 19338 43494 19352 43546
rect 19376 43494 19390 43546
rect 19390 43494 19402 43546
rect 19402 43494 19432 43546
rect 19456 43494 19466 43546
rect 19466 43494 19512 43546
rect 19216 43492 19272 43494
rect 19296 43492 19352 43494
rect 19376 43492 19432 43494
rect 19456 43492 19512 43494
rect 19614 43288 19670 43344
rect 17406 42200 17462 42256
rect 17958 42880 18014 42936
rect 18326 42200 18382 42256
rect 19154 43172 19210 43208
rect 19154 43152 19156 43172
rect 19156 43152 19208 43172
rect 19208 43152 19210 43172
rect 19216 42458 19272 42460
rect 19296 42458 19352 42460
rect 19376 42458 19432 42460
rect 19456 42458 19512 42460
rect 19216 42406 19262 42458
rect 19262 42406 19272 42458
rect 19296 42406 19326 42458
rect 19326 42406 19338 42458
rect 19338 42406 19352 42458
rect 19376 42406 19390 42458
rect 19390 42406 19402 42458
rect 19402 42406 19432 42458
rect 19456 42406 19466 42458
rect 19466 42406 19512 42458
rect 19216 42404 19272 42406
rect 19296 42404 19352 42406
rect 19376 42404 19432 42406
rect 19456 42404 19512 42406
rect 19154 42200 19210 42256
rect 19876 43002 19932 43004
rect 19956 43002 20012 43004
rect 20036 43002 20092 43004
rect 20116 43002 20172 43004
rect 19876 42950 19922 43002
rect 19922 42950 19932 43002
rect 19956 42950 19986 43002
rect 19986 42950 19998 43002
rect 19998 42950 20012 43002
rect 20036 42950 20050 43002
rect 20050 42950 20062 43002
rect 20062 42950 20092 43002
rect 20116 42950 20126 43002
rect 20126 42950 20172 43002
rect 19876 42948 19932 42950
rect 19956 42948 20012 42950
rect 20036 42948 20092 42950
rect 20116 42948 20172 42950
rect 19216 41370 19272 41372
rect 19296 41370 19352 41372
rect 19376 41370 19432 41372
rect 19456 41370 19512 41372
rect 19216 41318 19262 41370
rect 19262 41318 19272 41370
rect 19296 41318 19326 41370
rect 19326 41318 19338 41370
rect 19338 41318 19352 41370
rect 19376 41318 19390 41370
rect 19390 41318 19402 41370
rect 19402 41318 19432 41370
rect 19456 41318 19466 41370
rect 19466 41318 19512 41370
rect 19216 41316 19272 41318
rect 19296 41316 19352 41318
rect 19376 41316 19432 41318
rect 19456 41316 19512 41318
rect 19216 40282 19272 40284
rect 19296 40282 19352 40284
rect 19376 40282 19432 40284
rect 19456 40282 19512 40284
rect 19216 40230 19262 40282
rect 19262 40230 19272 40282
rect 19296 40230 19326 40282
rect 19326 40230 19338 40282
rect 19338 40230 19352 40282
rect 19376 40230 19390 40282
rect 19390 40230 19402 40282
rect 19402 40230 19432 40282
rect 19456 40230 19466 40282
rect 19466 40230 19512 40282
rect 19216 40228 19272 40230
rect 19296 40228 19352 40230
rect 19376 40228 19432 40230
rect 19456 40228 19512 40230
rect 19876 41914 19932 41916
rect 19956 41914 20012 41916
rect 20036 41914 20092 41916
rect 20116 41914 20172 41916
rect 19876 41862 19922 41914
rect 19922 41862 19932 41914
rect 19956 41862 19986 41914
rect 19986 41862 19998 41914
rect 19998 41862 20012 41914
rect 20036 41862 20050 41914
rect 20050 41862 20062 41914
rect 20062 41862 20092 41914
rect 20116 41862 20126 41914
rect 20126 41862 20172 41914
rect 19876 41860 19932 41862
rect 19956 41860 20012 41862
rect 20036 41860 20092 41862
rect 20116 41860 20172 41862
rect 19876 40826 19932 40828
rect 19956 40826 20012 40828
rect 20036 40826 20092 40828
rect 20116 40826 20172 40828
rect 19876 40774 19922 40826
rect 19922 40774 19932 40826
rect 19956 40774 19986 40826
rect 19986 40774 19998 40826
rect 19998 40774 20012 40826
rect 20036 40774 20050 40826
rect 20050 40774 20062 40826
rect 20062 40774 20092 40826
rect 20116 40774 20126 40826
rect 20126 40774 20172 40826
rect 19876 40772 19932 40774
rect 19956 40772 20012 40774
rect 20036 40772 20092 40774
rect 20116 40772 20172 40774
rect 19216 39194 19272 39196
rect 19296 39194 19352 39196
rect 19376 39194 19432 39196
rect 19456 39194 19512 39196
rect 19216 39142 19262 39194
rect 19262 39142 19272 39194
rect 19296 39142 19326 39194
rect 19326 39142 19338 39194
rect 19338 39142 19352 39194
rect 19376 39142 19390 39194
rect 19390 39142 19402 39194
rect 19402 39142 19432 39194
rect 19456 39142 19466 39194
rect 19466 39142 19512 39194
rect 19216 39140 19272 39142
rect 19296 39140 19352 39142
rect 19376 39140 19432 39142
rect 19456 39140 19512 39142
rect 16670 31900 16672 31920
rect 16672 31900 16724 31920
rect 16724 31900 16726 31920
rect 16670 31864 16726 31900
rect 11442 26138 11498 26140
rect 11522 26138 11578 26140
rect 11602 26138 11658 26140
rect 11682 26138 11738 26140
rect 11442 26086 11488 26138
rect 11488 26086 11498 26138
rect 11522 26086 11552 26138
rect 11552 26086 11564 26138
rect 11564 26086 11578 26138
rect 11602 26086 11616 26138
rect 11616 26086 11628 26138
rect 11628 26086 11658 26138
rect 11682 26086 11692 26138
rect 11692 26086 11738 26138
rect 11442 26084 11498 26086
rect 11522 26084 11578 26086
rect 11602 26084 11658 26086
rect 11682 26084 11738 26086
rect 4328 25594 4384 25596
rect 4408 25594 4464 25596
rect 4488 25594 4544 25596
rect 4568 25594 4624 25596
rect 4328 25542 4374 25594
rect 4374 25542 4384 25594
rect 4408 25542 4438 25594
rect 4438 25542 4450 25594
rect 4450 25542 4464 25594
rect 4488 25542 4502 25594
rect 4502 25542 4514 25594
rect 4514 25542 4544 25594
rect 4568 25542 4578 25594
rect 4578 25542 4624 25594
rect 4328 25540 4384 25542
rect 4408 25540 4464 25542
rect 4488 25540 4544 25542
rect 4568 25540 4624 25542
rect 3668 25050 3724 25052
rect 3748 25050 3804 25052
rect 3828 25050 3884 25052
rect 3908 25050 3964 25052
rect 3668 24998 3714 25050
rect 3714 24998 3724 25050
rect 3748 24998 3778 25050
rect 3778 24998 3790 25050
rect 3790 24998 3804 25050
rect 3828 24998 3842 25050
rect 3842 24998 3854 25050
rect 3854 24998 3884 25050
rect 3908 24998 3918 25050
rect 3918 24998 3964 25050
rect 3668 24996 3724 24998
rect 3748 24996 3804 24998
rect 3828 24996 3884 24998
rect 3908 24996 3964 24998
rect 12102 25594 12158 25596
rect 12182 25594 12238 25596
rect 12262 25594 12318 25596
rect 12342 25594 12398 25596
rect 12102 25542 12148 25594
rect 12148 25542 12158 25594
rect 12182 25542 12212 25594
rect 12212 25542 12224 25594
rect 12224 25542 12238 25594
rect 12262 25542 12276 25594
rect 12276 25542 12288 25594
rect 12288 25542 12318 25594
rect 12342 25542 12352 25594
rect 12352 25542 12398 25594
rect 12102 25540 12158 25542
rect 12182 25540 12238 25542
rect 12262 25540 12318 25542
rect 12342 25540 12398 25542
rect 11442 25050 11498 25052
rect 11522 25050 11578 25052
rect 11602 25050 11658 25052
rect 11682 25050 11738 25052
rect 11442 24998 11488 25050
rect 11488 24998 11498 25050
rect 11522 24998 11552 25050
rect 11552 24998 11564 25050
rect 11564 24998 11578 25050
rect 11602 24998 11616 25050
rect 11616 24998 11628 25050
rect 11628 24998 11658 25050
rect 11682 24998 11692 25050
rect 11692 24998 11738 25050
rect 11442 24996 11498 24998
rect 11522 24996 11578 24998
rect 11602 24996 11658 24998
rect 11682 24996 11738 24998
rect 4328 24506 4384 24508
rect 4408 24506 4464 24508
rect 4488 24506 4544 24508
rect 4568 24506 4624 24508
rect 4328 24454 4374 24506
rect 4374 24454 4384 24506
rect 4408 24454 4438 24506
rect 4438 24454 4450 24506
rect 4450 24454 4464 24506
rect 4488 24454 4502 24506
rect 4502 24454 4514 24506
rect 4514 24454 4544 24506
rect 4568 24454 4578 24506
rect 4578 24454 4624 24506
rect 4328 24452 4384 24454
rect 4408 24452 4464 24454
rect 4488 24452 4544 24454
rect 4568 24452 4624 24454
rect 3668 23962 3724 23964
rect 3748 23962 3804 23964
rect 3828 23962 3884 23964
rect 3908 23962 3964 23964
rect 3668 23910 3714 23962
rect 3714 23910 3724 23962
rect 3748 23910 3778 23962
rect 3778 23910 3790 23962
rect 3790 23910 3804 23962
rect 3828 23910 3842 23962
rect 3842 23910 3854 23962
rect 3854 23910 3884 23962
rect 3908 23910 3918 23962
rect 3918 23910 3964 23962
rect 3668 23908 3724 23910
rect 3748 23908 3804 23910
rect 3828 23908 3884 23910
rect 3908 23908 3964 23910
rect 12102 24506 12158 24508
rect 12182 24506 12238 24508
rect 12262 24506 12318 24508
rect 12342 24506 12398 24508
rect 12102 24454 12148 24506
rect 12148 24454 12158 24506
rect 12182 24454 12212 24506
rect 12212 24454 12224 24506
rect 12224 24454 12238 24506
rect 12262 24454 12276 24506
rect 12276 24454 12288 24506
rect 12288 24454 12318 24506
rect 12342 24454 12352 24506
rect 12352 24454 12398 24506
rect 12102 24452 12158 24454
rect 12182 24452 12238 24454
rect 12262 24452 12318 24454
rect 12342 24452 12398 24454
rect 11442 23962 11498 23964
rect 11522 23962 11578 23964
rect 11602 23962 11658 23964
rect 11682 23962 11738 23964
rect 11442 23910 11488 23962
rect 11488 23910 11498 23962
rect 11522 23910 11552 23962
rect 11552 23910 11564 23962
rect 11564 23910 11578 23962
rect 11602 23910 11616 23962
rect 11616 23910 11628 23962
rect 11628 23910 11658 23962
rect 11682 23910 11692 23962
rect 11692 23910 11738 23962
rect 11442 23908 11498 23910
rect 11522 23908 11578 23910
rect 11602 23908 11658 23910
rect 11682 23908 11738 23910
rect 4328 23418 4384 23420
rect 4408 23418 4464 23420
rect 4488 23418 4544 23420
rect 4568 23418 4624 23420
rect 4328 23366 4374 23418
rect 4374 23366 4384 23418
rect 4408 23366 4438 23418
rect 4438 23366 4450 23418
rect 4450 23366 4464 23418
rect 4488 23366 4502 23418
rect 4502 23366 4514 23418
rect 4514 23366 4544 23418
rect 4568 23366 4578 23418
rect 4578 23366 4624 23418
rect 4328 23364 4384 23366
rect 4408 23364 4464 23366
rect 4488 23364 4544 23366
rect 4568 23364 4624 23366
rect 12102 23418 12158 23420
rect 12182 23418 12238 23420
rect 12262 23418 12318 23420
rect 12342 23418 12398 23420
rect 12102 23366 12148 23418
rect 12148 23366 12158 23418
rect 12182 23366 12212 23418
rect 12212 23366 12224 23418
rect 12224 23366 12238 23418
rect 12262 23366 12276 23418
rect 12276 23366 12288 23418
rect 12288 23366 12318 23418
rect 12342 23366 12352 23418
rect 12352 23366 12398 23418
rect 12102 23364 12158 23366
rect 12182 23364 12238 23366
rect 12262 23364 12318 23366
rect 12342 23364 12398 23366
rect 3668 22874 3724 22876
rect 3748 22874 3804 22876
rect 3828 22874 3884 22876
rect 3908 22874 3964 22876
rect 3668 22822 3714 22874
rect 3714 22822 3724 22874
rect 3748 22822 3778 22874
rect 3778 22822 3790 22874
rect 3790 22822 3804 22874
rect 3828 22822 3842 22874
rect 3842 22822 3854 22874
rect 3854 22822 3884 22874
rect 3908 22822 3918 22874
rect 3918 22822 3964 22874
rect 3668 22820 3724 22822
rect 3748 22820 3804 22822
rect 3828 22820 3884 22822
rect 3908 22820 3964 22822
rect 11442 22874 11498 22876
rect 11522 22874 11578 22876
rect 11602 22874 11658 22876
rect 11682 22874 11738 22876
rect 11442 22822 11488 22874
rect 11488 22822 11498 22874
rect 11522 22822 11552 22874
rect 11552 22822 11564 22874
rect 11564 22822 11578 22874
rect 11602 22822 11616 22874
rect 11616 22822 11628 22874
rect 11628 22822 11658 22874
rect 11682 22822 11692 22874
rect 11692 22822 11738 22874
rect 11442 22820 11498 22822
rect 11522 22820 11578 22822
rect 11602 22820 11658 22822
rect 11682 22820 11738 22822
rect 4328 22330 4384 22332
rect 4408 22330 4464 22332
rect 4488 22330 4544 22332
rect 4568 22330 4624 22332
rect 4328 22278 4374 22330
rect 4374 22278 4384 22330
rect 4408 22278 4438 22330
rect 4438 22278 4450 22330
rect 4450 22278 4464 22330
rect 4488 22278 4502 22330
rect 4502 22278 4514 22330
rect 4514 22278 4544 22330
rect 4568 22278 4578 22330
rect 4578 22278 4624 22330
rect 4328 22276 4384 22278
rect 4408 22276 4464 22278
rect 4488 22276 4544 22278
rect 4568 22276 4624 22278
rect 12102 22330 12158 22332
rect 12182 22330 12238 22332
rect 12262 22330 12318 22332
rect 12342 22330 12398 22332
rect 12102 22278 12148 22330
rect 12148 22278 12158 22330
rect 12182 22278 12212 22330
rect 12212 22278 12224 22330
rect 12224 22278 12238 22330
rect 12262 22278 12276 22330
rect 12276 22278 12288 22330
rect 12288 22278 12318 22330
rect 12342 22278 12352 22330
rect 12352 22278 12398 22330
rect 12102 22276 12158 22278
rect 12182 22276 12238 22278
rect 12262 22276 12318 22278
rect 12342 22276 12398 22278
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 11442 21786 11498 21788
rect 11522 21786 11578 21788
rect 11602 21786 11658 21788
rect 11682 21786 11738 21788
rect 11442 21734 11488 21786
rect 11488 21734 11498 21786
rect 11522 21734 11552 21786
rect 11552 21734 11564 21786
rect 11564 21734 11578 21786
rect 11602 21734 11616 21786
rect 11616 21734 11628 21786
rect 11628 21734 11658 21786
rect 11682 21734 11692 21786
rect 11692 21734 11738 21786
rect 11442 21732 11498 21734
rect 11522 21732 11578 21734
rect 11602 21732 11658 21734
rect 11682 21732 11738 21734
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 12102 21242 12158 21244
rect 12182 21242 12238 21244
rect 12262 21242 12318 21244
rect 12342 21242 12398 21244
rect 12102 21190 12148 21242
rect 12148 21190 12158 21242
rect 12182 21190 12212 21242
rect 12212 21190 12224 21242
rect 12224 21190 12238 21242
rect 12262 21190 12276 21242
rect 12276 21190 12288 21242
rect 12288 21190 12318 21242
rect 12342 21190 12352 21242
rect 12352 21190 12398 21242
rect 12102 21188 12158 21190
rect 12182 21188 12238 21190
rect 12262 21188 12318 21190
rect 12342 21188 12398 21190
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 11442 20698 11498 20700
rect 11522 20698 11578 20700
rect 11602 20698 11658 20700
rect 11682 20698 11738 20700
rect 11442 20646 11488 20698
rect 11488 20646 11498 20698
rect 11522 20646 11552 20698
rect 11552 20646 11564 20698
rect 11564 20646 11578 20698
rect 11602 20646 11616 20698
rect 11616 20646 11628 20698
rect 11628 20646 11658 20698
rect 11682 20646 11692 20698
rect 11692 20646 11738 20698
rect 11442 20644 11498 20646
rect 11522 20644 11578 20646
rect 11602 20644 11658 20646
rect 11682 20644 11738 20646
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 12102 20154 12158 20156
rect 12182 20154 12238 20156
rect 12262 20154 12318 20156
rect 12342 20154 12398 20156
rect 12102 20102 12148 20154
rect 12148 20102 12158 20154
rect 12182 20102 12212 20154
rect 12212 20102 12224 20154
rect 12224 20102 12238 20154
rect 12262 20102 12276 20154
rect 12276 20102 12288 20154
rect 12288 20102 12318 20154
rect 12342 20102 12352 20154
rect 12352 20102 12398 20154
rect 12102 20100 12158 20102
rect 12182 20100 12238 20102
rect 12262 20100 12318 20102
rect 12342 20100 12398 20102
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 11442 19610 11498 19612
rect 11522 19610 11578 19612
rect 11602 19610 11658 19612
rect 11682 19610 11738 19612
rect 11442 19558 11488 19610
rect 11488 19558 11498 19610
rect 11522 19558 11552 19610
rect 11552 19558 11564 19610
rect 11564 19558 11578 19610
rect 11602 19558 11616 19610
rect 11616 19558 11628 19610
rect 11628 19558 11658 19610
rect 11682 19558 11692 19610
rect 11692 19558 11738 19610
rect 11442 19556 11498 19558
rect 11522 19556 11578 19558
rect 11602 19556 11658 19558
rect 11682 19556 11738 19558
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 12102 19066 12158 19068
rect 12182 19066 12238 19068
rect 12262 19066 12318 19068
rect 12342 19066 12398 19068
rect 12102 19014 12148 19066
rect 12148 19014 12158 19066
rect 12182 19014 12212 19066
rect 12212 19014 12224 19066
rect 12224 19014 12238 19066
rect 12262 19014 12276 19066
rect 12276 19014 12288 19066
rect 12288 19014 12318 19066
rect 12342 19014 12352 19066
rect 12352 19014 12398 19066
rect 12102 19012 12158 19014
rect 12182 19012 12238 19014
rect 12262 19012 12318 19014
rect 12342 19012 12398 19014
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 11442 18522 11498 18524
rect 11522 18522 11578 18524
rect 11602 18522 11658 18524
rect 11682 18522 11738 18524
rect 11442 18470 11488 18522
rect 11488 18470 11498 18522
rect 11522 18470 11552 18522
rect 11552 18470 11564 18522
rect 11564 18470 11578 18522
rect 11602 18470 11616 18522
rect 11616 18470 11628 18522
rect 11628 18470 11658 18522
rect 11682 18470 11692 18522
rect 11692 18470 11738 18522
rect 11442 18468 11498 18470
rect 11522 18468 11578 18470
rect 11602 18468 11658 18470
rect 11682 18468 11738 18470
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 12102 17978 12158 17980
rect 12182 17978 12238 17980
rect 12262 17978 12318 17980
rect 12342 17978 12398 17980
rect 12102 17926 12148 17978
rect 12148 17926 12158 17978
rect 12182 17926 12212 17978
rect 12212 17926 12224 17978
rect 12224 17926 12238 17978
rect 12262 17926 12276 17978
rect 12276 17926 12288 17978
rect 12288 17926 12318 17978
rect 12342 17926 12352 17978
rect 12352 17926 12398 17978
rect 12102 17924 12158 17926
rect 12182 17924 12238 17926
rect 12262 17924 12318 17926
rect 12342 17924 12398 17926
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 11442 17434 11498 17436
rect 11522 17434 11578 17436
rect 11602 17434 11658 17436
rect 11682 17434 11738 17436
rect 11442 17382 11488 17434
rect 11488 17382 11498 17434
rect 11522 17382 11552 17434
rect 11552 17382 11564 17434
rect 11564 17382 11578 17434
rect 11602 17382 11616 17434
rect 11616 17382 11628 17434
rect 11628 17382 11658 17434
rect 11682 17382 11692 17434
rect 11692 17382 11738 17434
rect 11442 17380 11498 17382
rect 11522 17380 11578 17382
rect 11602 17380 11658 17382
rect 11682 17380 11738 17382
rect 19430 38256 19486 38312
rect 19876 39738 19932 39740
rect 19956 39738 20012 39740
rect 20036 39738 20092 39740
rect 20116 39738 20172 39740
rect 19876 39686 19922 39738
rect 19922 39686 19932 39738
rect 19956 39686 19986 39738
rect 19986 39686 19998 39738
rect 19998 39686 20012 39738
rect 20036 39686 20050 39738
rect 20050 39686 20062 39738
rect 20062 39686 20092 39738
rect 20116 39686 20126 39738
rect 20126 39686 20172 39738
rect 19876 39684 19932 39686
rect 19956 39684 20012 39686
rect 20036 39684 20092 39686
rect 20116 39684 20172 39686
rect 20350 39344 20406 39400
rect 19614 38392 19670 38448
rect 20166 38800 20222 38856
rect 19876 38650 19932 38652
rect 19956 38650 20012 38652
rect 20036 38650 20092 38652
rect 20116 38650 20172 38652
rect 19876 38598 19922 38650
rect 19922 38598 19932 38650
rect 19956 38598 19986 38650
rect 19986 38598 19998 38650
rect 19998 38598 20012 38650
rect 20036 38598 20050 38650
rect 20050 38598 20062 38650
rect 20062 38598 20092 38650
rect 20116 38598 20126 38650
rect 20126 38598 20172 38650
rect 19876 38596 19932 38598
rect 19956 38596 20012 38598
rect 20036 38596 20092 38598
rect 20116 38596 20172 38598
rect 20166 38392 20222 38448
rect 19216 38106 19272 38108
rect 19296 38106 19352 38108
rect 19376 38106 19432 38108
rect 19456 38106 19512 38108
rect 19216 38054 19262 38106
rect 19262 38054 19272 38106
rect 19296 38054 19326 38106
rect 19326 38054 19338 38106
rect 19338 38054 19352 38106
rect 19376 38054 19390 38106
rect 19390 38054 19402 38106
rect 19402 38054 19432 38106
rect 19456 38054 19466 38106
rect 19466 38054 19512 38106
rect 19216 38052 19272 38054
rect 19296 38052 19352 38054
rect 19376 38052 19432 38054
rect 19456 38052 19512 38054
rect 19338 37868 19394 37904
rect 19338 37848 19340 37868
rect 19340 37848 19392 37868
rect 19392 37848 19394 37868
rect 19338 37304 19394 37360
rect 19522 37168 19578 37224
rect 19216 37018 19272 37020
rect 19296 37018 19352 37020
rect 19376 37018 19432 37020
rect 19456 37018 19512 37020
rect 19216 36966 19262 37018
rect 19262 36966 19272 37018
rect 19296 36966 19326 37018
rect 19326 36966 19338 37018
rect 19338 36966 19352 37018
rect 19376 36966 19390 37018
rect 19390 36966 19402 37018
rect 19402 36966 19432 37018
rect 19456 36966 19466 37018
rect 19466 36966 19512 37018
rect 19216 36964 19272 36966
rect 19296 36964 19352 36966
rect 19376 36964 19432 36966
rect 19456 36964 19512 36966
rect 19522 36760 19578 36816
rect 19062 36216 19118 36272
rect 18510 34060 18566 34096
rect 18510 34040 18512 34060
rect 18512 34040 18564 34060
rect 18564 34040 18566 34060
rect 19216 35930 19272 35932
rect 19296 35930 19352 35932
rect 19376 35930 19432 35932
rect 19456 35930 19512 35932
rect 19216 35878 19262 35930
rect 19262 35878 19272 35930
rect 19296 35878 19326 35930
rect 19326 35878 19338 35930
rect 19338 35878 19352 35930
rect 19376 35878 19390 35930
rect 19390 35878 19402 35930
rect 19402 35878 19432 35930
rect 19456 35878 19466 35930
rect 19466 35878 19512 35930
rect 19216 35876 19272 35878
rect 19296 35876 19352 35878
rect 19376 35876 19432 35878
rect 19456 35876 19512 35878
rect 19890 38120 19946 38176
rect 19798 37984 19854 38040
rect 20166 37984 20222 38040
rect 20074 37748 20076 37768
rect 20076 37748 20128 37768
rect 20128 37748 20130 37768
rect 20074 37712 20130 37748
rect 20534 38256 20590 38312
rect 19876 37562 19932 37564
rect 19956 37562 20012 37564
rect 20036 37562 20092 37564
rect 20116 37562 20172 37564
rect 19876 37510 19922 37562
rect 19922 37510 19932 37562
rect 19956 37510 19986 37562
rect 19986 37510 19998 37562
rect 19998 37510 20012 37562
rect 20036 37510 20050 37562
rect 20050 37510 20062 37562
rect 20062 37510 20092 37562
rect 20116 37510 20126 37562
rect 20126 37510 20172 37562
rect 19876 37508 19932 37510
rect 19956 37508 20012 37510
rect 20036 37508 20092 37510
rect 20116 37508 20172 37510
rect 20166 37324 20222 37360
rect 20166 37304 20168 37324
rect 20168 37304 20220 37324
rect 20220 37304 20222 37324
rect 19876 36474 19932 36476
rect 19956 36474 20012 36476
rect 20036 36474 20092 36476
rect 20116 36474 20172 36476
rect 19876 36422 19922 36474
rect 19922 36422 19932 36474
rect 19956 36422 19986 36474
rect 19986 36422 19998 36474
rect 19998 36422 20012 36474
rect 20036 36422 20050 36474
rect 20050 36422 20062 36474
rect 20062 36422 20092 36474
rect 20116 36422 20126 36474
rect 20126 36422 20172 36474
rect 19876 36420 19932 36422
rect 19956 36420 20012 36422
rect 20036 36420 20092 36422
rect 20116 36420 20172 36422
rect 19876 35386 19932 35388
rect 19956 35386 20012 35388
rect 20036 35386 20092 35388
rect 20116 35386 20172 35388
rect 19876 35334 19922 35386
rect 19922 35334 19932 35386
rect 19956 35334 19986 35386
rect 19986 35334 19998 35386
rect 19998 35334 20012 35386
rect 20036 35334 20050 35386
rect 20050 35334 20062 35386
rect 20062 35334 20092 35386
rect 20116 35334 20126 35386
rect 20126 35334 20172 35386
rect 19876 35332 19932 35334
rect 19956 35332 20012 35334
rect 20036 35332 20092 35334
rect 20116 35332 20172 35334
rect 19216 34842 19272 34844
rect 19296 34842 19352 34844
rect 19376 34842 19432 34844
rect 19456 34842 19512 34844
rect 19216 34790 19262 34842
rect 19262 34790 19272 34842
rect 19296 34790 19326 34842
rect 19326 34790 19338 34842
rect 19338 34790 19352 34842
rect 19376 34790 19390 34842
rect 19390 34790 19402 34842
rect 19402 34790 19432 34842
rect 19456 34790 19466 34842
rect 19466 34790 19512 34842
rect 19216 34788 19272 34790
rect 19296 34788 19352 34790
rect 19376 34788 19432 34790
rect 19456 34788 19512 34790
rect 18602 33904 18658 33960
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 12102 16890 12158 16892
rect 12182 16890 12238 16892
rect 12262 16890 12318 16892
rect 12342 16890 12398 16892
rect 12102 16838 12148 16890
rect 12148 16838 12158 16890
rect 12182 16838 12212 16890
rect 12212 16838 12224 16890
rect 12224 16838 12238 16890
rect 12262 16838 12276 16890
rect 12276 16838 12288 16890
rect 12288 16838 12318 16890
rect 12342 16838 12352 16890
rect 12352 16838 12398 16890
rect 12102 16836 12158 16838
rect 12182 16836 12238 16838
rect 12262 16836 12318 16838
rect 12342 16836 12398 16838
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 11442 16346 11498 16348
rect 11522 16346 11578 16348
rect 11602 16346 11658 16348
rect 11682 16346 11738 16348
rect 11442 16294 11488 16346
rect 11488 16294 11498 16346
rect 11522 16294 11552 16346
rect 11552 16294 11564 16346
rect 11564 16294 11578 16346
rect 11602 16294 11616 16346
rect 11616 16294 11628 16346
rect 11628 16294 11658 16346
rect 11682 16294 11692 16346
rect 11692 16294 11738 16346
rect 11442 16292 11498 16294
rect 11522 16292 11578 16294
rect 11602 16292 11658 16294
rect 11682 16292 11738 16294
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 12102 15802 12158 15804
rect 12182 15802 12238 15804
rect 12262 15802 12318 15804
rect 12342 15802 12398 15804
rect 12102 15750 12148 15802
rect 12148 15750 12158 15802
rect 12182 15750 12212 15802
rect 12212 15750 12224 15802
rect 12224 15750 12238 15802
rect 12262 15750 12276 15802
rect 12276 15750 12288 15802
rect 12288 15750 12318 15802
rect 12342 15750 12352 15802
rect 12352 15750 12398 15802
rect 12102 15748 12158 15750
rect 12182 15748 12238 15750
rect 12262 15748 12318 15750
rect 12342 15748 12398 15750
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 11442 15258 11498 15260
rect 11522 15258 11578 15260
rect 11602 15258 11658 15260
rect 11682 15258 11738 15260
rect 11442 15206 11488 15258
rect 11488 15206 11498 15258
rect 11522 15206 11552 15258
rect 11552 15206 11564 15258
rect 11564 15206 11578 15258
rect 11602 15206 11616 15258
rect 11616 15206 11628 15258
rect 11628 15206 11658 15258
rect 11682 15206 11692 15258
rect 11692 15206 11738 15258
rect 11442 15204 11498 15206
rect 11522 15204 11578 15206
rect 11602 15204 11658 15206
rect 11682 15204 11738 15206
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 12102 14714 12158 14716
rect 12182 14714 12238 14716
rect 12262 14714 12318 14716
rect 12342 14714 12398 14716
rect 12102 14662 12148 14714
rect 12148 14662 12158 14714
rect 12182 14662 12212 14714
rect 12212 14662 12224 14714
rect 12224 14662 12238 14714
rect 12262 14662 12276 14714
rect 12276 14662 12288 14714
rect 12288 14662 12318 14714
rect 12342 14662 12352 14714
rect 12352 14662 12398 14714
rect 12102 14660 12158 14662
rect 12182 14660 12238 14662
rect 12262 14660 12318 14662
rect 12342 14660 12398 14662
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 11442 14170 11498 14172
rect 11522 14170 11578 14172
rect 11602 14170 11658 14172
rect 11682 14170 11738 14172
rect 11442 14118 11488 14170
rect 11488 14118 11498 14170
rect 11522 14118 11552 14170
rect 11552 14118 11564 14170
rect 11564 14118 11578 14170
rect 11602 14118 11616 14170
rect 11616 14118 11628 14170
rect 11628 14118 11658 14170
rect 11682 14118 11692 14170
rect 11692 14118 11738 14170
rect 11442 14116 11498 14118
rect 11522 14116 11578 14118
rect 11602 14116 11658 14118
rect 11682 14116 11738 14118
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 12102 13626 12158 13628
rect 12182 13626 12238 13628
rect 12262 13626 12318 13628
rect 12342 13626 12398 13628
rect 12102 13574 12148 13626
rect 12148 13574 12158 13626
rect 12182 13574 12212 13626
rect 12212 13574 12224 13626
rect 12224 13574 12238 13626
rect 12262 13574 12276 13626
rect 12276 13574 12288 13626
rect 12288 13574 12318 13626
rect 12342 13574 12352 13626
rect 12352 13574 12398 13626
rect 12102 13572 12158 13574
rect 12182 13572 12238 13574
rect 12262 13572 12318 13574
rect 12342 13572 12398 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 11442 13082 11498 13084
rect 11522 13082 11578 13084
rect 11602 13082 11658 13084
rect 11682 13082 11738 13084
rect 11442 13030 11488 13082
rect 11488 13030 11498 13082
rect 11522 13030 11552 13082
rect 11552 13030 11564 13082
rect 11564 13030 11578 13082
rect 11602 13030 11616 13082
rect 11616 13030 11628 13082
rect 11628 13030 11658 13082
rect 11682 13030 11692 13082
rect 11692 13030 11738 13082
rect 11442 13028 11498 13030
rect 11522 13028 11578 13030
rect 11602 13028 11658 13030
rect 11682 13028 11738 13030
rect 17222 16632 17278 16688
rect 16946 15156 17002 15192
rect 16946 15136 16948 15156
rect 16948 15136 17000 15156
rect 17000 15136 17002 15156
rect 19154 33904 19210 33960
rect 19876 34298 19932 34300
rect 19956 34298 20012 34300
rect 20036 34298 20092 34300
rect 20116 34298 20172 34300
rect 19876 34246 19922 34298
rect 19922 34246 19932 34298
rect 19956 34246 19986 34298
rect 19986 34246 19998 34298
rect 19998 34246 20012 34298
rect 20036 34246 20050 34298
rect 20050 34246 20062 34298
rect 20062 34246 20092 34298
rect 20116 34246 20126 34298
rect 20126 34246 20172 34298
rect 19876 34244 19932 34246
rect 19956 34244 20012 34246
rect 20036 34244 20092 34246
rect 20116 34244 20172 34246
rect 19216 33754 19272 33756
rect 19296 33754 19352 33756
rect 19376 33754 19432 33756
rect 19456 33754 19512 33756
rect 19216 33702 19262 33754
rect 19262 33702 19272 33754
rect 19296 33702 19326 33754
rect 19326 33702 19338 33754
rect 19338 33702 19352 33754
rect 19376 33702 19390 33754
rect 19390 33702 19402 33754
rect 19402 33702 19432 33754
rect 19456 33702 19466 33754
rect 19466 33702 19512 33754
rect 19216 33700 19272 33702
rect 19296 33700 19352 33702
rect 19376 33700 19432 33702
rect 19456 33700 19512 33702
rect 19216 32666 19272 32668
rect 19296 32666 19352 32668
rect 19376 32666 19432 32668
rect 19456 32666 19512 32668
rect 19216 32614 19262 32666
rect 19262 32614 19272 32666
rect 19296 32614 19326 32666
rect 19326 32614 19338 32666
rect 19338 32614 19352 32666
rect 19376 32614 19390 32666
rect 19390 32614 19402 32666
rect 19402 32614 19432 32666
rect 19456 32614 19466 32666
rect 19466 32614 19512 32666
rect 19216 32612 19272 32614
rect 19296 32612 19352 32614
rect 19376 32612 19432 32614
rect 19456 32612 19512 32614
rect 19216 31578 19272 31580
rect 19296 31578 19352 31580
rect 19376 31578 19432 31580
rect 19456 31578 19512 31580
rect 19216 31526 19262 31578
rect 19262 31526 19272 31578
rect 19296 31526 19326 31578
rect 19326 31526 19338 31578
rect 19338 31526 19352 31578
rect 19376 31526 19390 31578
rect 19390 31526 19402 31578
rect 19402 31526 19432 31578
rect 19456 31526 19466 31578
rect 19466 31526 19512 31578
rect 19216 31524 19272 31526
rect 19296 31524 19352 31526
rect 19376 31524 19432 31526
rect 19456 31524 19512 31526
rect 19216 30490 19272 30492
rect 19296 30490 19352 30492
rect 19376 30490 19432 30492
rect 19456 30490 19512 30492
rect 19216 30438 19262 30490
rect 19262 30438 19272 30490
rect 19296 30438 19326 30490
rect 19326 30438 19338 30490
rect 19338 30438 19352 30490
rect 19376 30438 19390 30490
rect 19390 30438 19402 30490
rect 19402 30438 19432 30490
rect 19456 30438 19466 30490
rect 19466 30438 19512 30490
rect 19216 30436 19272 30438
rect 19296 30436 19352 30438
rect 19376 30436 19432 30438
rect 19456 30436 19512 30438
rect 19876 33210 19932 33212
rect 19956 33210 20012 33212
rect 20036 33210 20092 33212
rect 20116 33210 20172 33212
rect 19876 33158 19922 33210
rect 19922 33158 19932 33210
rect 19956 33158 19986 33210
rect 19986 33158 19998 33210
rect 19998 33158 20012 33210
rect 20036 33158 20050 33210
rect 20050 33158 20062 33210
rect 20062 33158 20092 33210
rect 20116 33158 20126 33210
rect 20126 33158 20172 33210
rect 19876 33156 19932 33158
rect 19956 33156 20012 33158
rect 20036 33156 20092 33158
rect 20116 33156 20172 33158
rect 19216 29402 19272 29404
rect 19296 29402 19352 29404
rect 19376 29402 19432 29404
rect 19456 29402 19512 29404
rect 19216 29350 19262 29402
rect 19262 29350 19272 29402
rect 19296 29350 19326 29402
rect 19326 29350 19338 29402
rect 19338 29350 19352 29402
rect 19376 29350 19390 29402
rect 19390 29350 19402 29402
rect 19402 29350 19432 29402
rect 19456 29350 19466 29402
rect 19466 29350 19512 29402
rect 19216 29348 19272 29350
rect 19296 29348 19352 29350
rect 19376 29348 19432 29350
rect 19456 29348 19512 29350
rect 19522 29144 19578 29200
rect 19216 28314 19272 28316
rect 19296 28314 19352 28316
rect 19376 28314 19432 28316
rect 19456 28314 19512 28316
rect 19216 28262 19262 28314
rect 19262 28262 19272 28314
rect 19296 28262 19326 28314
rect 19326 28262 19338 28314
rect 19338 28262 19352 28314
rect 19376 28262 19390 28314
rect 19390 28262 19402 28314
rect 19402 28262 19432 28314
rect 19456 28262 19466 28314
rect 19466 28262 19512 28314
rect 19216 28260 19272 28262
rect 19296 28260 19352 28262
rect 19376 28260 19432 28262
rect 19456 28260 19512 28262
rect 19216 27226 19272 27228
rect 19296 27226 19352 27228
rect 19376 27226 19432 27228
rect 19456 27226 19512 27228
rect 19216 27174 19262 27226
rect 19262 27174 19272 27226
rect 19296 27174 19326 27226
rect 19326 27174 19338 27226
rect 19338 27174 19352 27226
rect 19376 27174 19390 27226
rect 19390 27174 19402 27226
rect 19402 27174 19432 27226
rect 19456 27174 19466 27226
rect 19466 27174 19512 27226
rect 19216 27172 19272 27174
rect 19296 27172 19352 27174
rect 19376 27172 19432 27174
rect 19456 27172 19512 27174
rect 20074 32408 20130 32464
rect 20166 32308 20168 32328
rect 20168 32308 20220 32328
rect 20220 32308 20222 32328
rect 20166 32272 20222 32308
rect 19876 32122 19932 32124
rect 19956 32122 20012 32124
rect 20036 32122 20092 32124
rect 20116 32122 20172 32124
rect 19876 32070 19922 32122
rect 19922 32070 19932 32122
rect 19956 32070 19986 32122
rect 19986 32070 19998 32122
rect 19998 32070 20012 32122
rect 20036 32070 20050 32122
rect 20050 32070 20062 32122
rect 20062 32070 20092 32122
rect 20116 32070 20126 32122
rect 20126 32070 20172 32122
rect 19876 32068 19932 32070
rect 19956 32068 20012 32070
rect 20036 32068 20092 32070
rect 20116 32068 20172 32070
rect 21822 37304 21878 37360
rect 20810 37168 20866 37224
rect 20350 31864 20406 31920
rect 20350 31592 20406 31648
rect 19876 31034 19932 31036
rect 19956 31034 20012 31036
rect 20036 31034 20092 31036
rect 20116 31034 20172 31036
rect 19876 30982 19922 31034
rect 19922 30982 19932 31034
rect 19956 30982 19986 31034
rect 19986 30982 19998 31034
rect 19998 30982 20012 31034
rect 20036 30982 20050 31034
rect 20050 30982 20062 31034
rect 20062 30982 20092 31034
rect 20116 30982 20126 31034
rect 20126 30982 20172 31034
rect 19876 30980 19932 30982
rect 19956 30980 20012 30982
rect 20036 30980 20092 30982
rect 20116 30980 20172 30982
rect 19876 29946 19932 29948
rect 19956 29946 20012 29948
rect 20036 29946 20092 29948
rect 20116 29946 20172 29948
rect 19876 29894 19922 29946
rect 19922 29894 19932 29946
rect 19956 29894 19986 29946
rect 19986 29894 19998 29946
rect 19998 29894 20012 29946
rect 20036 29894 20050 29946
rect 20050 29894 20062 29946
rect 20062 29894 20092 29946
rect 20116 29894 20126 29946
rect 20126 29894 20172 29946
rect 19876 29892 19932 29894
rect 19956 29892 20012 29894
rect 20036 29892 20092 29894
rect 20116 29892 20172 29894
rect 19876 28858 19932 28860
rect 19956 28858 20012 28860
rect 20036 28858 20092 28860
rect 20116 28858 20172 28860
rect 19876 28806 19922 28858
rect 19922 28806 19932 28858
rect 19956 28806 19986 28858
rect 19986 28806 19998 28858
rect 19998 28806 20012 28858
rect 20036 28806 20050 28858
rect 20050 28806 20062 28858
rect 20062 28806 20092 28858
rect 20116 28806 20126 28858
rect 20126 28806 20172 28858
rect 19876 28804 19932 28806
rect 19956 28804 20012 28806
rect 20036 28804 20092 28806
rect 20116 28804 20172 28806
rect 21914 36660 21916 36680
rect 21916 36660 21968 36680
rect 21968 36660 21970 36680
rect 21914 36624 21970 36660
rect 20902 32444 20904 32464
rect 20904 32444 20956 32464
rect 20956 32444 20958 32464
rect 20902 32408 20958 32444
rect 23662 42236 23664 42256
rect 23664 42236 23716 42256
rect 23716 42236 23718 42256
rect 23662 42200 23718 42236
rect 26990 44634 27046 44636
rect 27070 44634 27126 44636
rect 27150 44634 27206 44636
rect 27230 44634 27286 44636
rect 26990 44582 27036 44634
rect 27036 44582 27046 44634
rect 27070 44582 27100 44634
rect 27100 44582 27112 44634
rect 27112 44582 27126 44634
rect 27150 44582 27164 44634
rect 27164 44582 27176 44634
rect 27176 44582 27206 44634
rect 27230 44582 27240 44634
rect 27240 44582 27286 44634
rect 26990 44580 27046 44582
rect 27070 44580 27126 44582
rect 27150 44580 27206 44582
rect 27230 44580 27286 44582
rect 28998 44648 29054 44704
rect 27650 44090 27706 44092
rect 27730 44090 27786 44092
rect 27810 44090 27866 44092
rect 27890 44090 27946 44092
rect 27650 44038 27696 44090
rect 27696 44038 27706 44090
rect 27730 44038 27760 44090
rect 27760 44038 27772 44090
rect 27772 44038 27786 44090
rect 27810 44038 27824 44090
rect 27824 44038 27836 44090
rect 27836 44038 27866 44090
rect 27890 44038 27900 44090
rect 27900 44038 27946 44090
rect 27650 44036 27706 44038
rect 27730 44036 27786 44038
rect 27810 44036 27866 44038
rect 27890 44036 27946 44038
rect 26990 43546 27046 43548
rect 27070 43546 27126 43548
rect 27150 43546 27206 43548
rect 27230 43546 27286 43548
rect 26990 43494 27036 43546
rect 27036 43494 27046 43546
rect 27070 43494 27100 43546
rect 27100 43494 27112 43546
rect 27112 43494 27126 43546
rect 27150 43494 27164 43546
rect 27164 43494 27176 43546
rect 27176 43494 27206 43546
rect 27230 43494 27240 43546
rect 27240 43494 27286 43546
rect 26990 43492 27046 43494
rect 27070 43492 27126 43494
rect 27150 43492 27206 43494
rect 27230 43492 27286 43494
rect 22098 36216 22154 36272
rect 22282 36100 22338 36136
rect 22282 36080 22284 36100
rect 22284 36080 22336 36100
rect 22336 36080 22338 36100
rect 19876 27770 19932 27772
rect 19956 27770 20012 27772
rect 20036 27770 20092 27772
rect 20116 27770 20172 27772
rect 19876 27718 19922 27770
rect 19922 27718 19932 27770
rect 19956 27718 19986 27770
rect 19986 27718 19998 27770
rect 19998 27718 20012 27770
rect 20036 27718 20050 27770
rect 20050 27718 20062 27770
rect 20062 27718 20092 27770
rect 20116 27718 20126 27770
rect 20126 27718 20172 27770
rect 19876 27716 19932 27718
rect 19956 27716 20012 27718
rect 20036 27716 20092 27718
rect 20116 27716 20172 27718
rect 18786 23604 18788 23624
rect 18788 23604 18840 23624
rect 18840 23604 18842 23624
rect 18786 23568 18842 23604
rect 19216 26138 19272 26140
rect 19296 26138 19352 26140
rect 19376 26138 19432 26140
rect 19456 26138 19512 26140
rect 19216 26086 19262 26138
rect 19262 26086 19272 26138
rect 19296 26086 19326 26138
rect 19326 26086 19338 26138
rect 19338 26086 19352 26138
rect 19376 26086 19390 26138
rect 19390 26086 19402 26138
rect 19402 26086 19432 26138
rect 19456 26086 19466 26138
rect 19466 26086 19512 26138
rect 19216 26084 19272 26086
rect 19296 26084 19352 26086
rect 19376 26084 19432 26086
rect 19456 26084 19512 26086
rect 19216 25050 19272 25052
rect 19296 25050 19352 25052
rect 19376 25050 19432 25052
rect 19456 25050 19512 25052
rect 19216 24998 19262 25050
rect 19262 24998 19272 25050
rect 19296 24998 19326 25050
rect 19326 24998 19338 25050
rect 19338 24998 19352 25050
rect 19376 24998 19390 25050
rect 19390 24998 19402 25050
rect 19402 24998 19432 25050
rect 19456 24998 19466 25050
rect 19466 24998 19512 25050
rect 19216 24996 19272 24998
rect 19296 24996 19352 24998
rect 19376 24996 19432 24998
rect 19456 24996 19512 24998
rect 19216 23962 19272 23964
rect 19296 23962 19352 23964
rect 19376 23962 19432 23964
rect 19456 23962 19512 23964
rect 19216 23910 19262 23962
rect 19262 23910 19272 23962
rect 19296 23910 19326 23962
rect 19326 23910 19338 23962
rect 19338 23910 19352 23962
rect 19376 23910 19390 23962
rect 19390 23910 19402 23962
rect 19402 23910 19432 23962
rect 19456 23910 19466 23962
rect 19466 23910 19512 23962
rect 19216 23908 19272 23910
rect 19296 23908 19352 23910
rect 19376 23908 19432 23910
rect 19456 23908 19512 23910
rect 19246 23588 19302 23624
rect 19246 23568 19248 23588
rect 19248 23568 19300 23588
rect 19300 23568 19302 23588
rect 19876 26682 19932 26684
rect 19956 26682 20012 26684
rect 20036 26682 20092 26684
rect 20116 26682 20172 26684
rect 19876 26630 19922 26682
rect 19922 26630 19932 26682
rect 19956 26630 19986 26682
rect 19986 26630 19998 26682
rect 19998 26630 20012 26682
rect 20036 26630 20050 26682
rect 20050 26630 20062 26682
rect 20062 26630 20092 26682
rect 20116 26630 20126 26682
rect 20126 26630 20172 26682
rect 19876 26628 19932 26630
rect 19956 26628 20012 26630
rect 20036 26628 20092 26630
rect 20116 26628 20172 26630
rect 20534 27376 20590 27432
rect 19876 25594 19932 25596
rect 19956 25594 20012 25596
rect 20036 25594 20092 25596
rect 20116 25594 20172 25596
rect 19876 25542 19922 25594
rect 19922 25542 19932 25594
rect 19956 25542 19986 25594
rect 19986 25542 19998 25594
rect 19998 25542 20012 25594
rect 20036 25542 20050 25594
rect 20050 25542 20062 25594
rect 20062 25542 20092 25594
rect 20116 25542 20126 25594
rect 20126 25542 20172 25594
rect 19876 25540 19932 25542
rect 19956 25540 20012 25542
rect 20036 25540 20092 25542
rect 20116 25540 20172 25542
rect 19876 24506 19932 24508
rect 19956 24506 20012 24508
rect 20036 24506 20092 24508
rect 20116 24506 20172 24508
rect 19876 24454 19922 24506
rect 19922 24454 19932 24506
rect 19956 24454 19986 24506
rect 19986 24454 19998 24506
rect 19998 24454 20012 24506
rect 20036 24454 20050 24506
rect 20050 24454 20062 24506
rect 20062 24454 20092 24506
rect 20116 24454 20126 24506
rect 20126 24454 20172 24506
rect 19876 24452 19932 24454
rect 19956 24452 20012 24454
rect 20036 24452 20092 24454
rect 20116 24452 20172 24454
rect 20258 24384 20314 24440
rect 20350 23860 20406 23896
rect 20350 23840 20352 23860
rect 20352 23840 20404 23860
rect 20404 23840 20406 23860
rect 19876 23418 19932 23420
rect 19956 23418 20012 23420
rect 20036 23418 20092 23420
rect 20116 23418 20172 23420
rect 19876 23366 19922 23418
rect 19922 23366 19932 23418
rect 19956 23366 19986 23418
rect 19986 23366 19998 23418
rect 19998 23366 20012 23418
rect 20036 23366 20050 23418
rect 20050 23366 20062 23418
rect 20062 23366 20092 23418
rect 20116 23366 20126 23418
rect 20126 23366 20172 23418
rect 19876 23364 19932 23366
rect 19956 23364 20012 23366
rect 20036 23364 20092 23366
rect 20116 23364 20172 23366
rect 19216 22874 19272 22876
rect 19296 22874 19352 22876
rect 19376 22874 19432 22876
rect 19456 22874 19512 22876
rect 19216 22822 19262 22874
rect 19262 22822 19272 22874
rect 19296 22822 19326 22874
rect 19326 22822 19338 22874
rect 19338 22822 19352 22874
rect 19376 22822 19390 22874
rect 19390 22822 19402 22874
rect 19402 22822 19432 22874
rect 19456 22822 19466 22874
rect 19466 22822 19512 22874
rect 19216 22820 19272 22822
rect 19296 22820 19352 22822
rect 19376 22820 19432 22822
rect 19456 22820 19512 22822
rect 19876 22330 19932 22332
rect 19956 22330 20012 22332
rect 20036 22330 20092 22332
rect 20116 22330 20172 22332
rect 19876 22278 19922 22330
rect 19922 22278 19932 22330
rect 19956 22278 19986 22330
rect 19986 22278 19998 22330
rect 19998 22278 20012 22330
rect 20036 22278 20050 22330
rect 20050 22278 20062 22330
rect 20062 22278 20092 22330
rect 20116 22278 20126 22330
rect 20126 22278 20172 22330
rect 19876 22276 19932 22278
rect 19956 22276 20012 22278
rect 20036 22276 20092 22278
rect 20116 22276 20172 22278
rect 19216 21786 19272 21788
rect 19296 21786 19352 21788
rect 19376 21786 19432 21788
rect 19456 21786 19512 21788
rect 19216 21734 19262 21786
rect 19262 21734 19272 21786
rect 19296 21734 19326 21786
rect 19326 21734 19338 21786
rect 19338 21734 19352 21786
rect 19376 21734 19390 21786
rect 19390 21734 19402 21786
rect 19402 21734 19432 21786
rect 19456 21734 19466 21786
rect 19466 21734 19512 21786
rect 19216 21732 19272 21734
rect 19296 21732 19352 21734
rect 19376 21732 19432 21734
rect 19456 21732 19512 21734
rect 19216 20698 19272 20700
rect 19296 20698 19352 20700
rect 19376 20698 19432 20700
rect 19456 20698 19512 20700
rect 19216 20646 19262 20698
rect 19262 20646 19272 20698
rect 19296 20646 19326 20698
rect 19326 20646 19338 20698
rect 19338 20646 19352 20698
rect 19376 20646 19390 20698
rect 19390 20646 19402 20698
rect 19402 20646 19432 20698
rect 19456 20646 19466 20698
rect 19466 20646 19512 20698
rect 19216 20644 19272 20646
rect 19296 20644 19352 20646
rect 19376 20644 19432 20646
rect 19456 20644 19512 20646
rect 19216 19610 19272 19612
rect 19296 19610 19352 19612
rect 19376 19610 19432 19612
rect 19456 19610 19512 19612
rect 19216 19558 19262 19610
rect 19262 19558 19272 19610
rect 19296 19558 19326 19610
rect 19326 19558 19338 19610
rect 19338 19558 19352 19610
rect 19376 19558 19390 19610
rect 19390 19558 19402 19610
rect 19402 19558 19432 19610
rect 19456 19558 19466 19610
rect 19466 19558 19512 19610
rect 19216 19556 19272 19558
rect 19296 19556 19352 19558
rect 19376 19556 19432 19558
rect 19456 19556 19512 19558
rect 19876 21242 19932 21244
rect 19956 21242 20012 21244
rect 20036 21242 20092 21244
rect 20116 21242 20172 21244
rect 19876 21190 19922 21242
rect 19922 21190 19932 21242
rect 19956 21190 19986 21242
rect 19986 21190 19998 21242
rect 19998 21190 20012 21242
rect 20036 21190 20050 21242
rect 20050 21190 20062 21242
rect 20062 21190 20092 21242
rect 20116 21190 20126 21242
rect 20126 21190 20172 21242
rect 19876 21188 19932 21190
rect 19956 21188 20012 21190
rect 20036 21188 20092 21190
rect 20116 21188 20172 21190
rect 19876 20154 19932 20156
rect 19956 20154 20012 20156
rect 20036 20154 20092 20156
rect 20116 20154 20172 20156
rect 19876 20102 19922 20154
rect 19922 20102 19932 20154
rect 19956 20102 19986 20154
rect 19986 20102 19998 20154
rect 19998 20102 20012 20154
rect 20036 20102 20050 20154
rect 20050 20102 20062 20154
rect 20062 20102 20092 20154
rect 20116 20102 20126 20154
rect 20126 20102 20172 20154
rect 19876 20100 19932 20102
rect 19956 20100 20012 20102
rect 20036 20100 20092 20102
rect 20116 20100 20172 20102
rect 19876 19066 19932 19068
rect 19956 19066 20012 19068
rect 20036 19066 20092 19068
rect 20116 19066 20172 19068
rect 19876 19014 19922 19066
rect 19922 19014 19932 19066
rect 19956 19014 19986 19066
rect 19986 19014 19998 19066
rect 19998 19014 20012 19066
rect 20036 19014 20050 19066
rect 20050 19014 20062 19066
rect 20062 19014 20092 19066
rect 20116 19014 20126 19066
rect 20126 19014 20172 19066
rect 19876 19012 19932 19014
rect 19956 19012 20012 19014
rect 20036 19012 20092 19014
rect 20116 19012 20172 19014
rect 19216 18522 19272 18524
rect 19296 18522 19352 18524
rect 19376 18522 19432 18524
rect 19456 18522 19512 18524
rect 19216 18470 19262 18522
rect 19262 18470 19272 18522
rect 19296 18470 19326 18522
rect 19326 18470 19338 18522
rect 19338 18470 19352 18522
rect 19376 18470 19390 18522
rect 19390 18470 19402 18522
rect 19402 18470 19432 18522
rect 19456 18470 19466 18522
rect 19466 18470 19512 18522
rect 19216 18468 19272 18470
rect 19296 18468 19352 18470
rect 19376 18468 19432 18470
rect 19456 18468 19512 18470
rect 19216 17434 19272 17436
rect 19296 17434 19352 17436
rect 19376 17434 19432 17436
rect 19456 17434 19512 17436
rect 19216 17382 19262 17434
rect 19262 17382 19272 17434
rect 19296 17382 19326 17434
rect 19326 17382 19338 17434
rect 19338 17382 19352 17434
rect 19376 17382 19390 17434
rect 19390 17382 19402 17434
rect 19402 17382 19432 17434
rect 19456 17382 19466 17434
rect 19466 17382 19512 17434
rect 19216 17380 19272 17382
rect 19296 17380 19352 17382
rect 19376 17380 19432 17382
rect 19456 17380 19512 17382
rect 19876 17978 19932 17980
rect 19956 17978 20012 17980
rect 20036 17978 20092 17980
rect 20116 17978 20172 17980
rect 19876 17926 19922 17978
rect 19922 17926 19932 17978
rect 19956 17926 19986 17978
rect 19986 17926 19998 17978
rect 19998 17926 20012 17978
rect 20036 17926 20050 17978
rect 20050 17926 20062 17978
rect 20062 17926 20092 17978
rect 20116 17926 20126 17978
rect 20126 17926 20172 17978
rect 19876 17924 19932 17926
rect 19956 17924 20012 17926
rect 20036 17924 20092 17926
rect 20116 17924 20172 17926
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 12102 12538 12158 12540
rect 12182 12538 12238 12540
rect 12262 12538 12318 12540
rect 12342 12538 12398 12540
rect 12102 12486 12148 12538
rect 12148 12486 12158 12538
rect 12182 12486 12212 12538
rect 12212 12486 12224 12538
rect 12224 12486 12238 12538
rect 12262 12486 12276 12538
rect 12276 12486 12288 12538
rect 12288 12486 12318 12538
rect 12342 12486 12352 12538
rect 12352 12486 12398 12538
rect 12102 12484 12158 12486
rect 12182 12484 12238 12486
rect 12262 12484 12318 12486
rect 12342 12484 12398 12486
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 11442 11994 11498 11996
rect 11522 11994 11578 11996
rect 11602 11994 11658 11996
rect 11682 11994 11738 11996
rect 11442 11942 11488 11994
rect 11488 11942 11498 11994
rect 11522 11942 11552 11994
rect 11552 11942 11564 11994
rect 11564 11942 11578 11994
rect 11602 11942 11616 11994
rect 11616 11942 11628 11994
rect 11628 11942 11658 11994
rect 11682 11942 11692 11994
rect 11692 11942 11738 11994
rect 11442 11940 11498 11942
rect 11522 11940 11578 11942
rect 11602 11940 11658 11942
rect 11682 11940 11738 11942
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 12102 11450 12158 11452
rect 12182 11450 12238 11452
rect 12262 11450 12318 11452
rect 12342 11450 12398 11452
rect 12102 11398 12148 11450
rect 12148 11398 12158 11450
rect 12182 11398 12212 11450
rect 12212 11398 12224 11450
rect 12224 11398 12238 11450
rect 12262 11398 12276 11450
rect 12276 11398 12288 11450
rect 12288 11398 12318 11450
rect 12342 11398 12352 11450
rect 12352 11398 12398 11450
rect 12102 11396 12158 11398
rect 12182 11396 12238 11398
rect 12262 11396 12318 11398
rect 12342 11396 12398 11398
rect 19876 16890 19932 16892
rect 19956 16890 20012 16892
rect 20036 16890 20092 16892
rect 20116 16890 20172 16892
rect 19876 16838 19922 16890
rect 19922 16838 19932 16890
rect 19956 16838 19986 16890
rect 19986 16838 19998 16890
rect 19998 16838 20012 16890
rect 20036 16838 20050 16890
rect 20050 16838 20062 16890
rect 20062 16838 20092 16890
rect 20116 16838 20126 16890
rect 20126 16838 20172 16890
rect 19876 16836 19932 16838
rect 19956 16836 20012 16838
rect 20036 16836 20092 16838
rect 20116 16836 20172 16838
rect 19614 16632 19670 16688
rect 19216 16346 19272 16348
rect 19296 16346 19352 16348
rect 19376 16346 19432 16348
rect 19456 16346 19512 16348
rect 19216 16294 19262 16346
rect 19262 16294 19272 16346
rect 19296 16294 19326 16346
rect 19326 16294 19338 16346
rect 19338 16294 19352 16346
rect 19376 16294 19390 16346
rect 19390 16294 19402 16346
rect 19402 16294 19432 16346
rect 19456 16294 19466 16346
rect 19466 16294 19512 16346
rect 19216 16292 19272 16294
rect 19296 16292 19352 16294
rect 19376 16292 19432 16294
rect 19456 16292 19512 16294
rect 20902 28464 20958 28520
rect 23938 41540 23994 41576
rect 23938 41520 23940 41540
rect 23940 41520 23992 41540
rect 23992 41520 23994 41540
rect 27650 43002 27706 43004
rect 27730 43002 27786 43004
rect 27810 43002 27866 43004
rect 27890 43002 27946 43004
rect 27650 42950 27696 43002
rect 27696 42950 27706 43002
rect 27730 42950 27760 43002
rect 27760 42950 27772 43002
rect 27772 42950 27786 43002
rect 27810 42950 27824 43002
rect 27824 42950 27836 43002
rect 27836 42950 27866 43002
rect 27890 42950 27900 43002
rect 27900 42950 27946 43002
rect 27650 42948 27706 42950
rect 27730 42948 27786 42950
rect 27810 42948 27866 42950
rect 27890 42948 27946 42950
rect 26990 42458 27046 42460
rect 27070 42458 27126 42460
rect 27150 42458 27206 42460
rect 27230 42458 27286 42460
rect 26990 42406 27036 42458
rect 27036 42406 27046 42458
rect 27070 42406 27100 42458
rect 27100 42406 27112 42458
rect 27112 42406 27126 42458
rect 27150 42406 27164 42458
rect 27164 42406 27176 42458
rect 27176 42406 27206 42458
rect 27230 42406 27240 42458
rect 27240 42406 27286 42458
rect 26990 42404 27046 42406
rect 27070 42404 27126 42406
rect 27150 42404 27206 42406
rect 27230 42404 27286 42406
rect 21638 24556 21640 24576
rect 21640 24556 21692 24576
rect 21692 24556 21694 24576
rect 21638 24520 21694 24556
rect 20810 17876 20866 17912
rect 20810 17856 20812 17876
rect 20812 17856 20864 17876
rect 20864 17856 20866 17876
rect 21914 28620 21970 28656
rect 21914 28600 21916 28620
rect 21916 28600 21968 28620
rect 21968 28600 21970 28620
rect 22558 32308 22560 32328
rect 22560 32308 22612 32328
rect 22612 32308 22614 32328
rect 22558 32272 22614 32308
rect 27650 41914 27706 41916
rect 27730 41914 27786 41916
rect 27810 41914 27866 41916
rect 27890 41914 27946 41916
rect 27650 41862 27696 41914
rect 27696 41862 27706 41914
rect 27730 41862 27760 41914
rect 27760 41862 27772 41914
rect 27772 41862 27786 41914
rect 27810 41862 27824 41914
rect 27824 41862 27836 41914
rect 27836 41862 27866 41914
rect 27890 41862 27900 41914
rect 27900 41862 27946 41914
rect 27650 41860 27706 41862
rect 27730 41860 27786 41862
rect 27810 41860 27866 41862
rect 27890 41860 27946 41862
rect 26990 41370 27046 41372
rect 27070 41370 27126 41372
rect 27150 41370 27206 41372
rect 27230 41370 27286 41372
rect 26990 41318 27036 41370
rect 27036 41318 27046 41370
rect 27070 41318 27100 41370
rect 27100 41318 27112 41370
rect 27112 41318 27126 41370
rect 27150 41318 27164 41370
rect 27164 41318 27176 41370
rect 27176 41318 27206 41370
rect 27230 41318 27240 41370
rect 27240 41318 27286 41370
rect 26990 41316 27046 41318
rect 27070 41316 27126 41318
rect 27150 41316 27206 41318
rect 27230 41316 27286 41318
rect 25870 38956 25926 38992
rect 25870 38936 25872 38956
rect 25872 38936 25924 38956
rect 25924 38936 25926 38956
rect 26990 40282 27046 40284
rect 27070 40282 27126 40284
rect 27150 40282 27206 40284
rect 27230 40282 27286 40284
rect 26990 40230 27036 40282
rect 27036 40230 27046 40282
rect 27070 40230 27100 40282
rect 27100 40230 27112 40282
rect 27112 40230 27126 40282
rect 27150 40230 27164 40282
rect 27164 40230 27176 40282
rect 27176 40230 27206 40282
rect 27230 40230 27240 40282
rect 27240 40230 27286 40282
rect 26990 40228 27046 40230
rect 27070 40228 27126 40230
rect 27150 40228 27206 40230
rect 27230 40228 27286 40230
rect 27650 40826 27706 40828
rect 27730 40826 27786 40828
rect 27810 40826 27866 40828
rect 27890 40826 27946 40828
rect 27650 40774 27696 40826
rect 27696 40774 27706 40826
rect 27730 40774 27760 40826
rect 27760 40774 27772 40826
rect 27772 40774 27786 40826
rect 27810 40774 27824 40826
rect 27824 40774 27836 40826
rect 27836 40774 27866 40826
rect 27890 40774 27900 40826
rect 27900 40774 27946 40826
rect 27650 40772 27706 40774
rect 27730 40772 27786 40774
rect 27810 40772 27866 40774
rect 27890 40772 27946 40774
rect 27650 39738 27706 39740
rect 27730 39738 27786 39740
rect 27810 39738 27866 39740
rect 27890 39738 27946 39740
rect 27650 39686 27696 39738
rect 27696 39686 27706 39738
rect 27730 39686 27760 39738
rect 27760 39686 27772 39738
rect 27772 39686 27786 39738
rect 27810 39686 27824 39738
rect 27824 39686 27836 39738
rect 27836 39686 27866 39738
rect 27890 39686 27900 39738
rect 27900 39686 27946 39738
rect 27650 39684 27706 39686
rect 27730 39684 27786 39686
rect 27810 39684 27866 39686
rect 27890 39684 27946 39686
rect 26990 39194 27046 39196
rect 27070 39194 27126 39196
rect 27150 39194 27206 39196
rect 27230 39194 27286 39196
rect 26990 39142 27036 39194
rect 27036 39142 27046 39194
rect 27070 39142 27100 39194
rect 27100 39142 27112 39194
rect 27112 39142 27126 39194
rect 27150 39142 27164 39194
rect 27164 39142 27176 39194
rect 27176 39142 27206 39194
rect 27230 39142 27240 39194
rect 27240 39142 27286 39194
rect 26990 39140 27046 39142
rect 27070 39140 27126 39142
rect 27150 39140 27206 39142
rect 27230 39140 27286 39142
rect 26990 38106 27046 38108
rect 27070 38106 27126 38108
rect 27150 38106 27206 38108
rect 27230 38106 27286 38108
rect 26990 38054 27036 38106
rect 27036 38054 27046 38106
rect 27070 38054 27100 38106
rect 27100 38054 27112 38106
rect 27112 38054 27126 38106
rect 27150 38054 27164 38106
rect 27164 38054 27176 38106
rect 27176 38054 27206 38106
rect 27230 38054 27240 38106
rect 27240 38054 27286 38106
rect 26990 38052 27046 38054
rect 27070 38052 27126 38054
rect 27150 38052 27206 38054
rect 27230 38052 27286 38054
rect 26990 37018 27046 37020
rect 27070 37018 27126 37020
rect 27150 37018 27206 37020
rect 27230 37018 27286 37020
rect 26990 36966 27036 37018
rect 27036 36966 27046 37018
rect 27070 36966 27100 37018
rect 27100 36966 27112 37018
rect 27112 36966 27126 37018
rect 27150 36966 27164 37018
rect 27164 36966 27176 37018
rect 27176 36966 27206 37018
rect 27230 36966 27240 37018
rect 27240 36966 27286 37018
rect 26990 36964 27046 36966
rect 27070 36964 27126 36966
rect 27150 36964 27206 36966
rect 27230 36964 27286 36966
rect 27710 38936 27766 38992
rect 27650 38650 27706 38652
rect 27730 38650 27786 38652
rect 27810 38650 27866 38652
rect 27890 38650 27946 38652
rect 27650 38598 27696 38650
rect 27696 38598 27706 38650
rect 27730 38598 27760 38650
rect 27760 38598 27772 38650
rect 27772 38598 27786 38650
rect 27810 38598 27824 38650
rect 27824 38598 27836 38650
rect 27836 38598 27866 38650
rect 27890 38598 27900 38650
rect 27900 38598 27946 38650
rect 27650 38596 27706 38598
rect 27730 38596 27786 38598
rect 27810 38596 27866 38598
rect 27890 38596 27946 38598
rect 27650 37562 27706 37564
rect 27730 37562 27786 37564
rect 27810 37562 27866 37564
rect 27890 37562 27946 37564
rect 27650 37510 27696 37562
rect 27696 37510 27706 37562
rect 27730 37510 27760 37562
rect 27760 37510 27772 37562
rect 27772 37510 27786 37562
rect 27810 37510 27824 37562
rect 27824 37510 27836 37562
rect 27836 37510 27866 37562
rect 27890 37510 27900 37562
rect 27900 37510 27946 37562
rect 27650 37508 27706 37510
rect 27730 37508 27786 37510
rect 27810 37508 27866 37510
rect 27890 37508 27946 37510
rect 27650 36474 27706 36476
rect 27730 36474 27786 36476
rect 27810 36474 27866 36476
rect 27890 36474 27946 36476
rect 27650 36422 27696 36474
rect 27696 36422 27706 36474
rect 27730 36422 27760 36474
rect 27760 36422 27772 36474
rect 27772 36422 27786 36474
rect 27810 36422 27824 36474
rect 27824 36422 27836 36474
rect 27836 36422 27866 36474
rect 27890 36422 27900 36474
rect 27900 36422 27946 36474
rect 27650 36420 27706 36422
rect 27730 36420 27786 36422
rect 27810 36420 27866 36422
rect 27890 36420 27946 36422
rect 26990 35930 27046 35932
rect 27070 35930 27126 35932
rect 27150 35930 27206 35932
rect 27230 35930 27286 35932
rect 26990 35878 27036 35930
rect 27036 35878 27046 35930
rect 27070 35878 27100 35930
rect 27100 35878 27112 35930
rect 27112 35878 27126 35930
rect 27150 35878 27164 35930
rect 27164 35878 27176 35930
rect 27176 35878 27206 35930
rect 27230 35878 27240 35930
rect 27240 35878 27286 35930
rect 26990 35876 27046 35878
rect 27070 35876 27126 35878
rect 27150 35876 27206 35878
rect 27230 35876 27286 35878
rect 27650 35386 27706 35388
rect 27730 35386 27786 35388
rect 27810 35386 27866 35388
rect 27890 35386 27946 35388
rect 27650 35334 27696 35386
rect 27696 35334 27706 35386
rect 27730 35334 27760 35386
rect 27760 35334 27772 35386
rect 27772 35334 27786 35386
rect 27810 35334 27824 35386
rect 27824 35334 27836 35386
rect 27836 35334 27866 35386
rect 27890 35334 27900 35386
rect 27900 35334 27946 35386
rect 27650 35332 27706 35334
rect 27730 35332 27786 35334
rect 27810 35332 27866 35334
rect 27890 35332 27946 35334
rect 26990 34842 27046 34844
rect 27070 34842 27126 34844
rect 27150 34842 27206 34844
rect 27230 34842 27286 34844
rect 26990 34790 27036 34842
rect 27036 34790 27046 34842
rect 27070 34790 27100 34842
rect 27100 34790 27112 34842
rect 27112 34790 27126 34842
rect 27150 34790 27164 34842
rect 27164 34790 27176 34842
rect 27176 34790 27206 34842
rect 27230 34790 27240 34842
rect 27240 34790 27286 34842
rect 26990 34788 27046 34790
rect 27070 34788 27126 34790
rect 27150 34788 27206 34790
rect 27230 34788 27286 34790
rect 27650 34298 27706 34300
rect 27730 34298 27786 34300
rect 27810 34298 27866 34300
rect 27890 34298 27946 34300
rect 27650 34246 27696 34298
rect 27696 34246 27706 34298
rect 27730 34246 27760 34298
rect 27760 34246 27772 34298
rect 27772 34246 27786 34298
rect 27810 34246 27824 34298
rect 27824 34246 27836 34298
rect 27836 34246 27866 34298
rect 27890 34246 27900 34298
rect 27900 34246 27946 34298
rect 27650 34244 27706 34246
rect 27730 34244 27786 34246
rect 27810 34244 27866 34246
rect 27890 34244 27946 34246
rect 23570 30232 23626 30288
rect 21914 24384 21970 24440
rect 22466 24384 22522 24440
rect 19876 15802 19932 15804
rect 19956 15802 20012 15804
rect 20036 15802 20092 15804
rect 20116 15802 20172 15804
rect 19876 15750 19922 15802
rect 19922 15750 19932 15802
rect 19956 15750 19986 15802
rect 19986 15750 19998 15802
rect 19998 15750 20012 15802
rect 20036 15750 20050 15802
rect 20050 15750 20062 15802
rect 20062 15750 20092 15802
rect 20116 15750 20126 15802
rect 20126 15750 20172 15802
rect 19876 15748 19932 15750
rect 19956 15748 20012 15750
rect 20036 15748 20092 15750
rect 20116 15748 20172 15750
rect 19216 15258 19272 15260
rect 19296 15258 19352 15260
rect 19376 15258 19432 15260
rect 19456 15258 19512 15260
rect 19216 15206 19262 15258
rect 19262 15206 19272 15258
rect 19296 15206 19326 15258
rect 19326 15206 19338 15258
rect 19338 15206 19352 15258
rect 19376 15206 19390 15258
rect 19390 15206 19402 15258
rect 19402 15206 19432 15258
rect 19456 15206 19466 15258
rect 19466 15206 19512 15258
rect 19216 15204 19272 15206
rect 19296 15204 19352 15206
rect 19376 15204 19432 15206
rect 19456 15204 19512 15206
rect 19876 14714 19932 14716
rect 19956 14714 20012 14716
rect 20036 14714 20092 14716
rect 20116 14714 20172 14716
rect 19876 14662 19922 14714
rect 19922 14662 19932 14714
rect 19956 14662 19986 14714
rect 19986 14662 19998 14714
rect 19998 14662 20012 14714
rect 20036 14662 20050 14714
rect 20050 14662 20062 14714
rect 20062 14662 20092 14714
rect 20116 14662 20126 14714
rect 20126 14662 20172 14714
rect 19876 14660 19932 14662
rect 19956 14660 20012 14662
rect 20036 14660 20092 14662
rect 20116 14660 20172 14662
rect 22098 17312 22154 17368
rect 23662 27376 23718 27432
rect 23202 22208 23258 22264
rect 23202 21428 23204 21448
rect 23204 21428 23256 21448
rect 23256 21428 23258 21448
rect 23202 21392 23258 21428
rect 23570 22208 23626 22264
rect 23754 21392 23810 21448
rect 24490 28056 24546 28112
rect 24122 24520 24178 24576
rect 24306 17312 24362 17368
rect 19216 14170 19272 14172
rect 19296 14170 19352 14172
rect 19376 14170 19432 14172
rect 19456 14170 19512 14172
rect 19216 14118 19262 14170
rect 19262 14118 19272 14170
rect 19296 14118 19326 14170
rect 19326 14118 19338 14170
rect 19338 14118 19352 14170
rect 19376 14118 19390 14170
rect 19390 14118 19402 14170
rect 19402 14118 19432 14170
rect 19456 14118 19466 14170
rect 19466 14118 19512 14170
rect 19216 14116 19272 14118
rect 19296 14116 19352 14118
rect 19376 14116 19432 14118
rect 19456 14116 19512 14118
rect 19876 13626 19932 13628
rect 19956 13626 20012 13628
rect 20036 13626 20092 13628
rect 20116 13626 20172 13628
rect 19876 13574 19922 13626
rect 19922 13574 19932 13626
rect 19956 13574 19986 13626
rect 19986 13574 19998 13626
rect 19998 13574 20012 13626
rect 20036 13574 20050 13626
rect 20050 13574 20062 13626
rect 20062 13574 20092 13626
rect 20116 13574 20126 13626
rect 20126 13574 20172 13626
rect 19876 13572 19932 13574
rect 19956 13572 20012 13574
rect 20036 13572 20092 13574
rect 20116 13572 20172 13574
rect 26698 30640 26754 30696
rect 26990 33754 27046 33756
rect 27070 33754 27126 33756
rect 27150 33754 27206 33756
rect 27230 33754 27286 33756
rect 26990 33702 27036 33754
rect 27036 33702 27046 33754
rect 27070 33702 27100 33754
rect 27100 33702 27112 33754
rect 27112 33702 27126 33754
rect 27150 33702 27164 33754
rect 27164 33702 27176 33754
rect 27176 33702 27206 33754
rect 27230 33702 27240 33754
rect 27240 33702 27286 33754
rect 26990 33700 27046 33702
rect 27070 33700 27126 33702
rect 27150 33700 27206 33702
rect 27230 33700 27286 33702
rect 27650 33210 27706 33212
rect 27730 33210 27786 33212
rect 27810 33210 27866 33212
rect 27890 33210 27946 33212
rect 27650 33158 27696 33210
rect 27696 33158 27706 33210
rect 27730 33158 27760 33210
rect 27760 33158 27772 33210
rect 27772 33158 27786 33210
rect 27810 33158 27824 33210
rect 27824 33158 27836 33210
rect 27836 33158 27866 33210
rect 27890 33158 27900 33210
rect 27900 33158 27946 33210
rect 27650 33156 27706 33158
rect 27730 33156 27786 33158
rect 27810 33156 27866 33158
rect 27890 33156 27946 33158
rect 26990 32666 27046 32668
rect 27070 32666 27126 32668
rect 27150 32666 27206 32668
rect 27230 32666 27286 32668
rect 26990 32614 27036 32666
rect 27036 32614 27046 32666
rect 27070 32614 27100 32666
rect 27100 32614 27112 32666
rect 27112 32614 27126 32666
rect 27150 32614 27164 32666
rect 27164 32614 27176 32666
rect 27176 32614 27206 32666
rect 27230 32614 27240 32666
rect 27240 32614 27286 32666
rect 26990 32612 27046 32614
rect 27070 32612 27126 32614
rect 27150 32612 27206 32614
rect 27230 32612 27286 32614
rect 26990 31578 27046 31580
rect 27070 31578 27126 31580
rect 27150 31578 27206 31580
rect 27230 31578 27286 31580
rect 26990 31526 27036 31578
rect 27036 31526 27046 31578
rect 27070 31526 27100 31578
rect 27100 31526 27112 31578
rect 27112 31526 27126 31578
rect 27150 31526 27164 31578
rect 27164 31526 27176 31578
rect 27176 31526 27206 31578
rect 27230 31526 27240 31578
rect 27240 31526 27286 31578
rect 26990 31524 27046 31526
rect 27070 31524 27126 31526
rect 27150 31524 27206 31526
rect 27230 31524 27286 31526
rect 26990 30490 27046 30492
rect 27070 30490 27126 30492
rect 27150 30490 27206 30492
rect 27230 30490 27286 30492
rect 26990 30438 27036 30490
rect 27036 30438 27046 30490
rect 27070 30438 27100 30490
rect 27100 30438 27112 30490
rect 27112 30438 27126 30490
rect 27150 30438 27164 30490
rect 27164 30438 27176 30490
rect 27176 30438 27206 30490
rect 27230 30438 27240 30490
rect 27240 30438 27286 30490
rect 26990 30436 27046 30438
rect 27070 30436 27126 30438
rect 27150 30436 27206 30438
rect 27230 30436 27286 30438
rect 27650 32122 27706 32124
rect 27730 32122 27786 32124
rect 27810 32122 27866 32124
rect 27890 32122 27946 32124
rect 27650 32070 27696 32122
rect 27696 32070 27706 32122
rect 27730 32070 27760 32122
rect 27760 32070 27772 32122
rect 27772 32070 27786 32122
rect 27810 32070 27824 32122
rect 27824 32070 27836 32122
rect 27836 32070 27866 32122
rect 27890 32070 27900 32122
rect 27900 32070 27946 32122
rect 27650 32068 27706 32070
rect 27730 32068 27786 32070
rect 27810 32068 27866 32070
rect 27890 32068 27946 32070
rect 27650 31034 27706 31036
rect 27730 31034 27786 31036
rect 27810 31034 27866 31036
rect 27890 31034 27946 31036
rect 27650 30982 27696 31034
rect 27696 30982 27706 31034
rect 27730 30982 27760 31034
rect 27760 30982 27772 31034
rect 27772 30982 27786 31034
rect 27810 30982 27824 31034
rect 27824 30982 27836 31034
rect 27836 30982 27866 31034
rect 27890 30982 27900 31034
rect 27900 30982 27946 31034
rect 27650 30980 27706 30982
rect 27730 30980 27786 30982
rect 27810 30980 27866 30982
rect 27890 30980 27946 30982
rect 26990 29402 27046 29404
rect 27070 29402 27126 29404
rect 27150 29402 27206 29404
rect 27230 29402 27286 29404
rect 26990 29350 27036 29402
rect 27036 29350 27046 29402
rect 27070 29350 27100 29402
rect 27100 29350 27112 29402
rect 27112 29350 27126 29402
rect 27150 29350 27164 29402
rect 27164 29350 27176 29402
rect 27176 29350 27206 29402
rect 27230 29350 27240 29402
rect 27240 29350 27286 29402
rect 26990 29348 27046 29350
rect 27070 29348 27126 29350
rect 27150 29348 27206 29350
rect 27230 29348 27286 29350
rect 27650 29946 27706 29948
rect 27730 29946 27786 29948
rect 27810 29946 27866 29948
rect 27890 29946 27946 29948
rect 27650 29894 27696 29946
rect 27696 29894 27706 29946
rect 27730 29894 27760 29946
rect 27760 29894 27772 29946
rect 27772 29894 27786 29946
rect 27810 29894 27824 29946
rect 27824 29894 27836 29946
rect 27836 29894 27866 29946
rect 27890 29894 27900 29946
rect 27900 29894 27946 29946
rect 27650 29892 27706 29894
rect 27730 29892 27786 29894
rect 27810 29892 27866 29894
rect 27890 29892 27946 29894
rect 26990 28314 27046 28316
rect 27070 28314 27126 28316
rect 27150 28314 27206 28316
rect 27230 28314 27286 28316
rect 26990 28262 27036 28314
rect 27036 28262 27046 28314
rect 27070 28262 27100 28314
rect 27100 28262 27112 28314
rect 27112 28262 27126 28314
rect 27150 28262 27164 28314
rect 27164 28262 27176 28314
rect 27176 28262 27206 28314
rect 27230 28262 27240 28314
rect 27240 28262 27286 28314
rect 26990 28260 27046 28262
rect 27070 28260 27126 28262
rect 27150 28260 27206 28262
rect 27230 28260 27286 28262
rect 26990 27226 27046 27228
rect 27070 27226 27126 27228
rect 27150 27226 27206 27228
rect 27230 27226 27286 27228
rect 26990 27174 27036 27226
rect 27036 27174 27046 27226
rect 27070 27174 27100 27226
rect 27100 27174 27112 27226
rect 27112 27174 27126 27226
rect 27150 27174 27164 27226
rect 27164 27174 27176 27226
rect 27176 27174 27206 27226
rect 27230 27174 27240 27226
rect 27240 27174 27286 27226
rect 26990 27172 27046 27174
rect 27070 27172 27126 27174
rect 27150 27172 27206 27174
rect 27230 27172 27286 27174
rect 26238 22072 26294 22128
rect 26422 22208 26478 22264
rect 25686 17856 25742 17912
rect 26422 22072 26478 22128
rect 26990 26138 27046 26140
rect 27070 26138 27126 26140
rect 27150 26138 27206 26140
rect 27230 26138 27286 26140
rect 26990 26086 27036 26138
rect 27036 26086 27046 26138
rect 27070 26086 27100 26138
rect 27100 26086 27112 26138
rect 27112 26086 27126 26138
rect 27150 26086 27164 26138
rect 27164 26086 27176 26138
rect 27176 26086 27206 26138
rect 27230 26086 27240 26138
rect 27240 26086 27286 26138
rect 26990 26084 27046 26086
rect 27070 26084 27126 26086
rect 27150 26084 27206 26086
rect 27230 26084 27286 26086
rect 26990 25050 27046 25052
rect 27070 25050 27126 25052
rect 27150 25050 27206 25052
rect 27230 25050 27286 25052
rect 26990 24998 27036 25050
rect 27036 24998 27046 25050
rect 27070 24998 27100 25050
rect 27100 24998 27112 25050
rect 27112 24998 27126 25050
rect 27150 24998 27164 25050
rect 27164 24998 27176 25050
rect 27176 24998 27206 25050
rect 27230 24998 27240 25050
rect 27240 24998 27286 25050
rect 26990 24996 27046 24998
rect 27070 24996 27126 24998
rect 27150 24996 27206 24998
rect 27230 24996 27286 24998
rect 27650 28858 27706 28860
rect 27730 28858 27786 28860
rect 27810 28858 27866 28860
rect 27890 28858 27946 28860
rect 27650 28806 27696 28858
rect 27696 28806 27706 28858
rect 27730 28806 27760 28858
rect 27760 28806 27772 28858
rect 27772 28806 27786 28858
rect 27810 28806 27824 28858
rect 27824 28806 27836 28858
rect 27836 28806 27866 28858
rect 27890 28806 27900 28858
rect 27900 28806 27946 28858
rect 27650 28804 27706 28806
rect 27730 28804 27786 28806
rect 27810 28804 27866 28806
rect 27890 28804 27946 28806
rect 27650 27770 27706 27772
rect 27730 27770 27786 27772
rect 27810 27770 27866 27772
rect 27890 27770 27946 27772
rect 27650 27718 27696 27770
rect 27696 27718 27706 27770
rect 27730 27718 27760 27770
rect 27760 27718 27772 27770
rect 27772 27718 27786 27770
rect 27810 27718 27824 27770
rect 27824 27718 27836 27770
rect 27836 27718 27866 27770
rect 27890 27718 27900 27770
rect 27900 27718 27946 27770
rect 27650 27716 27706 27718
rect 27730 27716 27786 27718
rect 27810 27716 27866 27718
rect 27890 27716 27946 27718
rect 27650 26682 27706 26684
rect 27730 26682 27786 26684
rect 27810 26682 27866 26684
rect 27890 26682 27946 26684
rect 27650 26630 27696 26682
rect 27696 26630 27706 26682
rect 27730 26630 27760 26682
rect 27760 26630 27772 26682
rect 27772 26630 27786 26682
rect 27810 26630 27824 26682
rect 27824 26630 27836 26682
rect 27836 26630 27866 26682
rect 27890 26630 27900 26682
rect 27900 26630 27946 26682
rect 27650 26628 27706 26630
rect 27730 26628 27786 26630
rect 27810 26628 27866 26630
rect 27890 26628 27946 26630
rect 27710 25744 27766 25800
rect 27650 25594 27706 25596
rect 27730 25594 27786 25596
rect 27810 25594 27866 25596
rect 27890 25594 27946 25596
rect 27650 25542 27696 25594
rect 27696 25542 27706 25594
rect 27730 25542 27760 25594
rect 27760 25542 27772 25594
rect 27772 25542 27786 25594
rect 27810 25542 27824 25594
rect 27824 25542 27836 25594
rect 27836 25542 27866 25594
rect 27890 25542 27900 25594
rect 27900 25542 27946 25594
rect 27650 25540 27706 25542
rect 27730 25540 27786 25542
rect 27810 25540 27866 25542
rect 27890 25540 27946 25542
rect 28078 25608 28134 25664
rect 26990 23962 27046 23964
rect 27070 23962 27126 23964
rect 27150 23962 27206 23964
rect 27230 23962 27286 23964
rect 26990 23910 27036 23962
rect 27036 23910 27046 23962
rect 27070 23910 27100 23962
rect 27100 23910 27112 23962
rect 27112 23910 27126 23962
rect 27150 23910 27164 23962
rect 27164 23910 27176 23962
rect 27176 23910 27206 23962
rect 27230 23910 27240 23962
rect 27240 23910 27286 23962
rect 26990 23908 27046 23910
rect 27070 23908 27126 23910
rect 27150 23908 27206 23910
rect 27230 23908 27286 23910
rect 26990 22874 27046 22876
rect 27070 22874 27126 22876
rect 27150 22874 27206 22876
rect 27230 22874 27286 22876
rect 26990 22822 27036 22874
rect 27036 22822 27046 22874
rect 27070 22822 27100 22874
rect 27100 22822 27112 22874
rect 27112 22822 27126 22874
rect 27150 22822 27164 22874
rect 27164 22822 27176 22874
rect 27176 22822 27206 22874
rect 27230 22822 27240 22874
rect 27240 22822 27286 22874
rect 26990 22820 27046 22822
rect 27070 22820 27126 22822
rect 27150 22820 27206 22822
rect 27230 22820 27286 22822
rect 27158 22636 27214 22672
rect 27158 22616 27160 22636
rect 27160 22616 27212 22636
rect 27212 22616 27214 22636
rect 26990 21786 27046 21788
rect 27070 21786 27126 21788
rect 27150 21786 27206 21788
rect 27230 21786 27286 21788
rect 26990 21734 27036 21786
rect 27036 21734 27046 21786
rect 27070 21734 27100 21786
rect 27100 21734 27112 21786
rect 27112 21734 27126 21786
rect 27150 21734 27164 21786
rect 27164 21734 27176 21786
rect 27176 21734 27206 21786
rect 27230 21734 27240 21786
rect 27240 21734 27286 21786
rect 26990 21732 27046 21734
rect 27070 21732 27126 21734
rect 27150 21732 27206 21734
rect 27230 21732 27286 21734
rect 27650 24506 27706 24508
rect 27730 24506 27786 24508
rect 27810 24506 27866 24508
rect 27890 24506 27946 24508
rect 27650 24454 27696 24506
rect 27696 24454 27706 24506
rect 27730 24454 27760 24506
rect 27760 24454 27772 24506
rect 27772 24454 27786 24506
rect 27810 24454 27824 24506
rect 27824 24454 27836 24506
rect 27836 24454 27866 24506
rect 27890 24454 27900 24506
rect 27900 24454 27946 24506
rect 27650 24452 27706 24454
rect 27730 24452 27786 24454
rect 27810 24452 27866 24454
rect 27890 24452 27946 24454
rect 27650 23418 27706 23420
rect 27730 23418 27786 23420
rect 27810 23418 27866 23420
rect 27890 23418 27946 23420
rect 27650 23366 27696 23418
rect 27696 23366 27706 23418
rect 27730 23366 27760 23418
rect 27760 23366 27772 23418
rect 27772 23366 27786 23418
rect 27810 23366 27824 23418
rect 27824 23366 27836 23418
rect 27836 23366 27866 23418
rect 27890 23366 27900 23418
rect 27900 23366 27946 23418
rect 27650 23364 27706 23366
rect 27730 23364 27786 23366
rect 27810 23364 27866 23366
rect 27890 23364 27946 23366
rect 28538 25744 28594 25800
rect 27618 22480 27674 22536
rect 27650 22330 27706 22332
rect 27730 22330 27786 22332
rect 27810 22330 27866 22332
rect 27890 22330 27946 22332
rect 27650 22278 27696 22330
rect 27696 22278 27706 22330
rect 27730 22278 27760 22330
rect 27760 22278 27772 22330
rect 27772 22278 27786 22330
rect 27810 22278 27824 22330
rect 27824 22278 27836 22330
rect 27836 22278 27866 22330
rect 27890 22278 27900 22330
rect 27900 22278 27946 22330
rect 27650 22276 27706 22278
rect 27730 22276 27786 22278
rect 27810 22276 27866 22278
rect 27890 22276 27946 22278
rect 26990 20698 27046 20700
rect 27070 20698 27126 20700
rect 27150 20698 27206 20700
rect 27230 20698 27286 20700
rect 26990 20646 27036 20698
rect 27036 20646 27046 20698
rect 27070 20646 27100 20698
rect 27100 20646 27112 20698
rect 27112 20646 27126 20698
rect 27150 20646 27164 20698
rect 27164 20646 27176 20698
rect 27176 20646 27206 20698
rect 27230 20646 27240 20698
rect 27240 20646 27286 20698
rect 26990 20644 27046 20646
rect 27070 20644 27126 20646
rect 27150 20644 27206 20646
rect 27230 20644 27286 20646
rect 26990 19610 27046 19612
rect 27070 19610 27126 19612
rect 27150 19610 27206 19612
rect 27230 19610 27286 19612
rect 26990 19558 27036 19610
rect 27036 19558 27046 19610
rect 27070 19558 27100 19610
rect 27100 19558 27112 19610
rect 27112 19558 27126 19610
rect 27150 19558 27164 19610
rect 27164 19558 27176 19610
rect 27176 19558 27206 19610
rect 27230 19558 27240 19610
rect 27240 19558 27286 19610
rect 26990 19556 27046 19558
rect 27070 19556 27126 19558
rect 27150 19556 27206 19558
rect 27230 19556 27286 19558
rect 26990 18522 27046 18524
rect 27070 18522 27126 18524
rect 27150 18522 27206 18524
rect 27230 18522 27286 18524
rect 26990 18470 27036 18522
rect 27036 18470 27046 18522
rect 27070 18470 27100 18522
rect 27100 18470 27112 18522
rect 27112 18470 27126 18522
rect 27150 18470 27164 18522
rect 27164 18470 27176 18522
rect 27176 18470 27206 18522
rect 27230 18470 27240 18522
rect 27240 18470 27286 18522
rect 26990 18468 27046 18470
rect 27070 18468 27126 18470
rect 27150 18468 27206 18470
rect 27230 18468 27286 18470
rect 26990 17434 27046 17436
rect 27070 17434 27126 17436
rect 27150 17434 27206 17436
rect 27230 17434 27286 17436
rect 26990 17382 27036 17434
rect 27036 17382 27046 17434
rect 27070 17382 27100 17434
rect 27100 17382 27112 17434
rect 27112 17382 27126 17434
rect 27150 17382 27164 17434
rect 27164 17382 27176 17434
rect 27176 17382 27206 17434
rect 27230 17382 27240 17434
rect 27240 17382 27286 17434
rect 26990 17380 27046 17382
rect 27070 17380 27126 17382
rect 27150 17380 27206 17382
rect 27230 17380 27286 17382
rect 27650 21242 27706 21244
rect 27730 21242 27786 21244
rect 27810 21242 27866 21244
rect 27890 21242 27946 21244
rect 27650 21190 27696 21242
rect 27696 21190 27706 21242
rect 27730 21190 27760 21242
rect 27760 21190 27772 21242
rect 27772 21190 27786 21242
rect 27810 21190 27824 21242
rect 27824 21190 27836 21242
rect 27836 21190 27866 21242
rect 27890 21190 27900 21242
rect 27900 21190 27946 21242
rect 27650 21188 27706 21190
rect 27730 21188 27786 21190
rect 27810 21188 27866 21190
rect 27890 21188 27946 21190
rect 27650 20154 27706 20156
rect 27730 20154 27786 20156
rect 27810 20154 27866 20156
rect 27890 20154 27946 20156
rect 27650 20102 27696 20154
rect 27696 20102 27706 20154
rect 27730 20102 27760 20154
rect 27760 20102 27772 20154
rect 27772 20102 27786 20154
rect 27810 20102 27824 20154
rect 27824 20102 27836 20154
rect 27836 20102 27866 20154
rect 27890 20102 27900 20154
rect 27900 20102 27946 20154
rect 27650 20100 27706 20102
rect 27730 20100 27786 20102
rect 27810 20100 27866 20102
rect 27890 20100 27946 20102
rect 27650 19066 27706 19068
rect 27730 19066 27786 19068
rect 27810 19066 27866 19068
rect 27890 19066 27946 19068
rect 27650 19014 27696 19066
rect 27696 19014 27706 19066
rect 27730 19014 27760 19066
rect 27760 19014 27772 19066
rect 27772 19014 27786 19066
rect 27810 19014 27824 19066
rect 27824 19014 27836 19066
rect 27836 19014 27866 19066
rect 27890 19014 27900 19066
rect 27900 19014 27946 19066
rect 27650 19012 27706 19014
rect 27730 19012 27786 19014
rect 27810 19012 27866 19014
rect 27890 19012 27946 19014
rect 28630 22616 28686 22672
rect 27650 17978 27706 17980
rect 27730 17978 27786 17980
rect 27810 17978 27866 17980
rect 27890 17978 27946 17980
rect 27650 17926 27696 17978
rect 27696 17926 27706 17978
rect 27730 17926 27760 17978
rect 27760 17926 27772 17978
rect 27772 17926 27786 17978
rect 27810 17926 27824 17978
rect 27824 17926 27836 17978
rect 27836 17926 27866 17978
rect 27890 17926 27900 17978
rect 27900 17926 27946 17978
rect 27650 17924 27706 17926
rect 27730 17924 27786 17926
rect 27810 17924 27866 17926
rect 27890 17924 27946 17926
rect 27650 16890 27706 16892
rect 27730 16890 27786 16892
rect 27810 16890 27866 16892
rect 27890 16890 27946 16892
rect 27650 16838 27696 16890
rect 27696 16838 27706 16890
rect 27730 16838 27760 16890
rect 27760 16838 27772 16890
rect 27772 16838 27786 16890
rect 27810 16838 27824 16890
rect 27824 16838 27836 16890
rect 27836 16838 27866 16890
rect 27890 16838 27900 16890
rect 27900 16838 27946 16890
rect 27650 16836 27706 16838
rect 27730 16836 27786 16838
rect 27810 16836 27866 16838
rect 27890 16836 27946 16838
rect 26882 16652 26938 16688
rect 26882 16632 26884 16652
rect 26884 16632 26936 16652
rect 26936 16632 26938 16652
rect 26990 16346 27046 16348
rect 27070 16346 27126 16348
rect 27150 16346 27206 16348
rect 27230 16346 27286 16348
rect 26990 16294 27036 16346
rect 27036 16294 27046 16346
rect 27070 16294 27100 16346
rect 27100 16294 27112 16346
rect 27112 16294 27126 16346
rect 27150 16294 27164 16346
rect 27164 16294 27176 16346
rect 27176 16294 27206 16346
rect 27230 16294 27240 16346
rect 27240 16294 27286 16346
rect 26990 16292 27046 16294
rect 27070 16292 27126 16294
rect 27150 16292 27206 16294
rect 27230 16292 27286 16294
rect 19216 13082 19272 13084
rect 19296 13082 19352 13084
rect 19376 13082 19432 13084
rect 19456 13082 19512 13084
rect 19216 13030 19262 13082
rect 19262 13030 19272 13082
rect 19296 13030 19326 13082
rect 19326 13030 19338 13082
rect 19338 13030 19352 13082
rect 19376 13030 19390 13082
rect 19390 13030 19402 13082
rect 19402 13030 19432 13082
rect 19456 13030 19466 13082
rect 19466 13030 19512 13082
rect 19216 13028 19272 13030
rect 19296 13028 19352 13030
rect 19376 13028 19432 13030
rect 19456 13028 19512 13030
rect 26990 15258 27046 15260
rect 27070 15258 27126 15260
rect 27150 15258 27206 15260
rect 27230 15258 27286 15260
rect 26990 15206 27036 15258
rect 27036 15206 27046 15258
rect 27070 15206 27100 15258
rect 27100 15206 27112 15258
rect 27112 15206 27126 15258
rect 27150 15206 27164 15258
rect 27164 15206 27176 15258
rect 27176 15206 27206 15258
rect 27230 15206 27240 15258
rect 27240 15206 27286 15258
rect 26990 15204 27046 15206
rect 27070 15204 27126 15206
rect 27150 15204 27206 15206
rect 27230 15204 27286 15206
rect 27650 15802 27706 15804
rect 27730 15802 27786 15804
rect 27810 15802 27866 15804
rect 27890 15802 27946 15804
rect 27650 15750 27696 15802
rect 27696 15750 27706 15802
rect 27730 15750 27760 15802
rect 27760 15750 27772 15802
rect 27772 15750 27786 15802
rect 27810 15750 27824 15802
rect 27824 15750 27836 15802
rect 27836 15750 27866 15802
rect 27890 15750 27900 15802
rect 27900 15750 27946 15802
rect 27650 15748 27706 15750
rect 27730 15748 27786 15750
rect 27810 15748 27866 15750
rect 27890 15748 27946 15750
rect 27650 14714 27706 14716
rect 27730 14714 27786 14716
rect 27810 14714 27866 14716
rect 27890 14714 27946 14716
rect 27650 14662 27696 14714
rect 27696 14662 27706 14714
rect 27730 14662 27760 14714
rect 27760 14662 27772 14714
rect 27772 14662 27786 14714
rect 27810 14662 27824 14714
rect 27824 14662 27836 14714
rect 27836 14662 27866 14714
rect 27890 14662 27900 14714
rect 27900 14662 27946 14714
rect 27650 14660 27706 14662
rect 27730 14660 27786 14662
rect 27810 14660 27866 14662
rect 27890 14660 27946 14662
rect 26990 14170 27046 14172
rect 27070 14170 27126 14172
rect 27150 14170 27206 14172
rect 27230 14170 27286 14172
rect 26990 14118 27036 14170
rect 27036 14118 27046 14170
rect 27070 14118 27100 14170
rect 27100 14118 27112 14170
rect 27112 14118 27126 14170
rect 27150 14118 27164 14170
rect 27164 14118 27176 14170
rect 27176 14118 27206 14170
rect 27230 14118 27240 14170
rect 27240 14118 27286 14170
rect 26990 14116 27046 14118
rect 27070 14116 27126 14118
rect 27150 14116 27206 14118
rect 27230 14116 27286 14118
rect 27650 13626 27706 13628
rect 27730 13626 27786 13628
rect 27810 13626 27866 13628
rect 27890 13626 27946 13628
rect 27650 13574 27696 13626
rect 27696 13574 27706 13626
rect 27730 13574 27760 13626
rect 27760 13574 27772 13626
rect 27772 13574 27786 13626
rect 27810 13574 27824 13626
rect 27824 13574 27836 13626
rect 27836 13574 27866 13626
rect 27890 13574 27900 13626
rect 27900 13574 27946 13626
rect 27650 13572 27706 13574
rect 27730 13572 27786 13574
rect 27810 13572 27866 13574
rect 27890 13572 27946 13574
rect 26990 13082 27046 13084
rect 27070 13082 27126 13084
rect 27150 13082 27206 13084
rect 27230 13082 27286 13084
rect 26990 13030 27036 13082
rect 27036 13030 27046 13082
rect 27070 13030 27100 13082
rect 27100 13030 27112 13082
rect 27112 13030 27126 13082
rect 27150 13030 27164 13082
rect 27164 13030 27176 13082
rect 27176 13030 27206 13082
rect 27230 13030 27240 13082
rect 27240 13030 27286 13082
rect 26990 13028 27046 13030
rect 27070 13028 27126 13030
rect 27150 13028 27206 13030
rect 27230 13028 27286 13030
rect 19876 12538 19932 12540
rect 19956 12538 20012 12540
rect 20036 12538 20092 12540
rect 20116 12538 20172 12540
rect 19876 12486 19922 12538
rect 19922 12486 19932 12538
rect 19956 12486 19986 12538
rect 19986 12486 19998 12538
rect 19998 12486 20012 12538
rect 20036 12486 20050 12538
rect 20050 12486 20062 12538
rect 20062 12486 20092 12538
rect 20116 12486 20126 12538
rect 20126 12486 20172 12538
rect 19876 12484 19932 12486
rect 19956 12484 20012 12486
rect 20036 12484 20092 12486
rect 20116 12484 20172 12486
rect 27650 12538 27706 12540
rect 27730 12538 27786 12540
rect 27810 12538 27866 12540
rect 27890 12538 27946 12540
rect 27650 12486 27696 12538
rect 27696 12486 27706 12538
rect 27730 12486 27760 12538
rect 27760 12486 27772 12538
rect 27772 12486 27786 12538
rect 27810 12486 27824 12538
rect 27824 12486 27836 12538
rect 27836 12486 27866 12538
rect 27890 12486 27900 12538
rect 27900 12486 27946 12538
rect 27650 12484 27706 12486
rect 27730 12484 27786 12486
rect 27810 12484 27866 12486
rect 27890 12484 27946 12486
rect 19216 11994 19272 11996
rect 19296 11994 19352 11996
rect 19376 11994 19432 11996
rect 19456 11994 19512 11996
rect 19216 11942 19262 11994
rect 19262 11942 19272 11994
rect 19296 11942 19326 11994
rect 19326 11942 19338 11994
rect 19338 11942 19352 11994
rect 19376 11942 19390 11994
rect 19390 11942 19402 11994
rect 19402 11942 19432 11994
rect 19456 11942 19466 11994
rect 19466 11942 19512 11994
rect 19216 11940 19272 11942
rect 19296 11940 19352 11942
rect 19376 11940 19432 11942
rect 19456 11940 19512 11942
rect 26990 11994 27046 11996
rect 27070 11994 27126 11996
rect 27150 11994 27206 11996
rect 27230 11994 27286 11996
rect 26990 11942 27036 11994
rect 27036 11942 27046 11994
rect 27070 11942 27100 11994
rect 27100 11942 27112 11994
rect 27112 11942 27126 11994
rect 27150 11942 27164 11994
rect 27164 11942 27176 11994
rect 27176 11942 27206 11994
rect 27230 11942 27240 11994
rect 27240 11942 27286 11994
rect 26990 11940 27046 11942
rect 27070 11940 27126 11942
rect 27150 11940 27206 11942
rect 27230 11940 27286 11942
rect 19876 11450 19932 11452
rect 19956 11450 20012 11452
rect 20036 11450 20092 11452
rect 20116 11450 20172 11452
rect 19876 11398 19922 11450
rect 19922 11398 19932 11450
rect 19956 11398 19986 11450
rect 19986 11398 19998 11450
rect 19998 11398 20012 11450
rect 20036 11398 20050 11450
rect 20050 11398 20062 11450
rect 20062 11398 20092 11450
rect 20116 11398 20126 11450
rect 20126 11398 20172 11450
rect 19876 11396 19932 11398
rect 19956 11396 20012 11398
rect 20036 11396 20092 11398
rect 20116 11396 20172 11398
rect 27650 11450 27706 11452
rect 27730 11450 27786 11452
rect 27810 11450 27866 11452
rect 27890 11450 27946 11452
rect 27650 11398 27696 11450
rect 27696 11398 27706 11450
rect 27730 11398 27760 11450
rect 27760 11398 27772 11450
rect 27772 11398 27786 11450
rect 27810 11398 27824 11450
rect 27824 11398 27836 11450
rect 27836 11398 27866 11450
rect 27890 11398 27900 11450
rect 27900 11398 27946 11450
rect 27650 11396 27706 11398
rect 27730 11396 27786 11398
rect 27810 11396 27866 11398
rect 27890 11396 27946 11398
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 11442 10906 11498 10908
rect 11522 10906 11578 10908
rect 11602 10906 11658 10908
rect 11682 10906 11738 10908
rect 11442 10854 11488 10906
rect 11488 10854 11498 10906
rect 11522 10854 11552 10906
rect 11552 10854 11564 10906
rect 11564 10854 11578 10906
rect 11602 10854 11616 10906
rect 11616 10854 11628 10906
rect 11628 10854 11658 10906
rect 11682 10854 11692 10906
rect 11692 10854 11738 10906
rect 11442 10852 11498 10854
rect 11522 10852 11578 10854
rect 11602 10852 11658 10854
rect 11682 10852 11738 10854
rect 19216 10906 19272 10908
rect 19296 10906 19352 10908
rect 19376 10906 19432 10908
rect 19456 10906 19512 10908
rect 19216 10854 19262 10906
rect 19262 10854 19272 10906
rect 19296 10854 19326 10906
rect 19326 10854 19338 10906
rect 19338 10854 19352 10906
rect 19376 10854 19390 10906
rect 19390 10854 19402 10906
rect 19402 10854 19432 10906
rect 19456 10854 19466 10906
rect 19466 10854 19512 10906
rect 19216 10852 19272 10854
rect 19296 10852 19352 10854
rect 19376 10852 19432 10854
rect 19456 10852 19512 10854
rect 26990 10906 27046 10908
rect 27070 10906 27126 10908
rect 27150 10906 27206 10908
rect 27230 10906 27286 10908
rect 26990 10854 27036 10906
rect 27036 10854 27046 10906
rect 27070 10854 27100 10906
rect 27100 10854 27112 10906
rect 27112 10854 27126 10906
rect 27150 10854 27164 10906
rect 27164 10854 27176 10906
rect 27176 10854 27206 10906
rect 27230 10854 27240 10906
rect 27240 10854 27286 10906
rect 26990 10852 27046 10854
rect 27070 10852 27126 10854
rect 27150 10852 27206 10854
rect 27230 10852 27286 10854
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 12102 10362 12158 10364
rect 12182 10362 12238 10364
rect 12262 10362 12318 10364
rect 12342 10362 12398 10364
rect 12102 10310 12148 10362
rect 12148 10310 12158 10362
rect 12182 10310 12212 10362
rect 12212 10310 12224 10362
rect 12224 10310 12238 10362
rect 12262 10310 12276 10362
rect 12276 10310 12288 10362
rect 12288 10310 12318 10362
rect 12342 10310 12352 10362
rect 12352 10310 12398 10362
rect 12102 10308 12158 10310
rect 12182 10308 12238 10310
rect 12262 10308 12318 10310
rect 12342 10308 12398 10310
rect 19876 10362 19932 10364
rect 19956 10362 20012 10364
rect 20036 10362 20092 10364
rect 20116 10362 20172 10364
rect 19876 10310 19922 10362
rect 19922 10310 19932 10362
rect 19956 10310 19986 10362
rect 19986 10310 19998 10362
rect 19998 10310 20012 10362
rect 20036 10310 20050 10362
rect 20050 10310 20062 10362
rect 20062 10310 20092 10362
rect 20116 10310 20126 10362
rect 20126 10310 20172 10362
rect 19876 10308 19932 10310
rect 19956 10308 20012 10310
rect 20036 10308 20092 10310
rect 20116 10308 20172 10310
rect 27650 10362 27706 10364
rect 27730 10362 27786 10364
rect 27810 10362 27866 10364
rect 27890 10362 27946 10364
rect 27650 10310 27696 10362
rect 27696 10310 27706 10362
rect 27730 10310 27760 10362
rect 27760 10310 27772 10362
rect 27772 10310 27786 10362
rect 27810 10310 27824 10362
rect 27824 10310 27836 10362
rect 27836 10310 27866 10362
rect 27890 10310 27900 10362
rect 27900 10310 27946 10362
rect 27650 10308 27706 10310
rect 27730 10308 27786 10310
rect 27810 10308 27866 10310
rect 27890 10308 27946 10310
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 11442 9818 11498 9820
rect 11522 9818 11578 9820
rect 11602 9818 11658 9820
rect 11682 9818 11738 9820
rect 11442 9766 11488 9818
rect 11488 9766 11498 9818
rect 11522 9766 11552 9818
rect 11552 9766 11564 9818
rect 11564 9766 11578 9818
rect 11602 9766 11616 9818
rect 11616 9766 11628 9818
rect 11628 9766 11658 9818
rect 11682 9766 11692 9818
rect 11692 9766 11738 9818
rect 11442 9764 11498 9766
rect 11522 9764 11578 9766
rect 11602 9764 11658 9766
rect 11682 9764 11738 9766
rect 19216 9818 19272 9820
rect 19296 9818 19352 9820
rect 19376 9818 19432 9820
rect 19456 9818 19512 9820
rect 19216 9766 19262 9818
rect 19262 9766 19272 9818
rect 19296 9766 19326 9818
rect 19326 9766 19338 9818
rect 19338 9766 19352 9818
rect 19376 9766 19390 9818
rect 19390 9766 19402 9818
rect 19402 9766 19432 9818
rect 19456 9766 19466 9818
rect 19466 9766 19512 9818
rect 19216 9764 19272 9766
rect 19296 9764 19352 9766
rect 19376 9764 19432 9766
rect 19456 9764 19512 9766
rect 26990 9818 27046 9820
rect 27070 9818 27126 9820
rect 27150 9818 27206 9820
rect 27230 9818 27286 9820
rect 26990 9766 27036 9818
rect 27036 9766 27046 9818
rect 27070 9766 27100 9818
rect 27100 9766 27112 9818
rect 27112 9766 27126 9818
rect 27150 9766 27164 9818
rect 27164 9766 27176 9818
rect 27176 9766 27206 9818
rect 27230 9766 27240 9818
rect 27240 9766 27286 9818
rect 26990 9764 27046 9766
rect 27070 9764 27126 9766
rect 27150 9764 27206 9766
rect 27230 9764 27286 9766
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 12102 9274 12158 9276
rect 12182 9274 12238 9276
rect 12262 9274 12318 9276
rect 12342 9274 12398 9276
rect 12102 9222 12148 9274
rect 12148 9222 12158 9274
rect 12182 9222 12212 9274
rect 12212 9222 12224 9274
rect 12224 9222 12238 9274
rect 12262 9222 12276 9274
rect 12276 9222 12288 9274
rect 12288 9222 12318 9274
rect 12342 9222 12352 9274
rect 12352 9222 12398 9274
rect 12102 9220 12158 9222
rect 12182 9220 12238 9222
rect 12262 9220 12318 9222
rect 12342 9220 12398 9222
rect 19876 9274 19932 9276
rect 19956 9274 20012 9276
rect 20036 9274 20092 9276
rect 20116 9274 20172 9276
rect 19876 9222 19922 9274
rect 19922 9222 19932 9274
rect 19956 9222 19986 9274
rect 19986 9222 19998 9274
rect 19998 9222 20012 9274
rect 20036 9222 20050 9274
rect 20050 9222 20062 9274
rect 20062 9222 20092 9274
rect 20116 9222 20126 9274
rect 20126 9222 20172 9274
rect 19876 9220 19932 9222
rect 19956 9220 20012 9222
rect 20036 9220 20092 9222
rect 20116 9220 20172 9222
rect 27650 9274 27706 9276
rect 27730 9274 27786 9276
rect 27810 9274 27866 9276
rect 27890 9274 27946 9276
rect 27650 9222 27696 9274
rect 27696 9222 27706 9274
rect 27730 9222 27760 9274
rect 27760 9222 27772 9274
rect 27772 9222 27786 9274
rect 27810 9222 27824 9274
rect 27824 9222 27836 9274
rect 27836 9222 27866 9274
rect 27890 9222 27900 9274
rect 27900 9222 27946 9274
rect 27650 9220 27706 9222
rect 27730 9220 27786 9222
rect 27810 9220 27866 9222
rect 27890 9220 27946 9222
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 11442 8730 11498 8732
rect 11522 8730 11578 8732
rect 11602 8730 11658 8732
rect 11682 8730 11738 8732
rect 11442 8678 11488 8730
rect 11488 8678 11498 8730
rect 11522 8678 11552 8730
rect 11552 8678 11564 8730
rect 11564 8678 11578 8730
rect 11602 8678 11616 8730
rect 11616 8678 11628 8730
rect 11628 8678 11658 8730
rect 11682 8678 11692 8730
rect 11692 8678 11738 8730
rect 11442 8676 11498 8678
rect 11522 8676 11578 8678
rect 11602 8676 11658 8678
rect 11682 8676 11738 8678
rect 19216 8730 19272 8732
rect 19296 8730 19352 8732
rect 19376 8730 19432 8732
rect 19456 8730 19512 8732
rect 19216 8678 19262 8730
rect 19262 8678 19272 8730
rect 19296 8678 19326 8730
rect 19326 8678 19338 8730
rect 19338 8678 19352 8730
rect 19376 8678 19390 8730
rect 19390 8678 19402 8730
rect 19402 8678 19432 8730
rect 19456 8678 19466 8730
rect 19466 8678 19512 8730
rect 19216 8676 19272 8678
rect 19296 8676 19352 8678
rect 19376 8676 19432 8678
rect 19456 8676 19512 8678
rect 26990 8730 27046 8732
rect 27070 8730 27126 8732
rect 27150 8730 27206 8732
rect 27230 8730 27286 8732
rect 26990 8678 27036 8730
rect 27036 8678 27046 8730
rect 27070 8678 27100 8730
rect 27100 8678 27112 8730
rect 27112 8678 27126 8730
rect 27150 8678 27164 8730
rect 27164 8678 27176 8730
rect 27176 8678 27206 8730
rect 27230 8678 27240 8730
rect 27240 8678 27286 8730
rect 26990 8676 27046 8678
rect 27070 8676 27126 8678
rect 27150 8676 27206 8678
rect 27230 8676 27286 8678
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 12102 8186 12158 8188
rect 12182 8186 12238 8188
rect 12262 8186 12318 8188
rect 12342 8186 12398 8188
rect 12102 8134 12148 8186
rect 12148 8134 12158 8186
rect 12182 8134 12212 8186
rect 12212 8134 12224 8186
rect 12224 8134 12238 8186
rect 12262 8134 12276 8186
rect 12276 8134 12288 8186
rect 12288 8134 12318 8186
rect 12342 8134 12352 8186
rect 12352 8134 12398 8186
rect 12102 8132 12158 8134
rect 12182 8132 12238 8134
rect 12262 8132 12318 8134
rect 12342 8132 12398 8134
rect 19876 8186 19932 8188
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 19876 8134 19922 8186
rect 19922 8134 19932 8186
rect 19956 8134 19986 8186
rect 19986 8134 19998 8186
rect 19998 8134 20012 8186
rect 20036 8134 20050 8186
rect 20050 8134 20062 8186
rect 20062 8134 20092 8186
rect 20116 8134 20126 8186
rect 20126 8134 20172 8186
rect 19876 8132 19932 8134
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 27650 8186 27706 8188
rect 27730 8186 27786 8188
rect 27810 8186 27866 8188
rect 27890 8186 27946 8188
rect 27650 8134 27696 8186
rect 27696 8134 27706 8186
rect 27730 8134 27760 8186
rect 27760 8134 27772 8186
rect 27772 8134 27786 8186
rect 27810 8134 27824 8186
rect 27824 8134 27836 8186
rect 27836 8134 27866 8186
rect 27890 8134 27900 8186
rect 27900 8134 27946 8186
rect 27650 8132 27706 8134
rect 27730 8132 27786 8134
rect 27810 8132 27866 8134
rect 27890 8132 27946 8134
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 11442 7642 11498 7644
rect 11522 7642 11578 7644
rect 11602 7642 11658 7644
rect 11682 7642 11738 7644
rect 11442 7590 11488 7642
rect 11488 7590 11498 7642
rect 11522 7590 11552 7642
rect 11552 7590 11564 7642
rect 11564 7590 11578 7642
rect 11602 7590 11616 7642
rect 11616 7590 11628 7642
rect 11628 7590 11658 7642
rect 11682 7590 11692 7642
rect 11692 7590 11738 7642
rect 11442 7588 11498 7590
rect 11522 7588 11578 7590
rect 11602 7588 11658 7590
rect 11682 7588 11738 7590
rect 19216 7642 19272 7644
rect 19296 7642 19352 7644
rect 19376 7642 19432 7644
rect 19456 7642 19512 7644
rect 19216 7590 19262 7642
rect 19262 7590 19272 7642
rect 19296 7590 19326 7642
rect 19326 7590 19338 7642
rect 19338 7590 19352 7642
rect 19376 7590 19390 7642
rect 19390 7590 19402 7642
rect 19402 7590 19432 7642
rect 19456 7590 19466 7642
rect 19466 7590 19512 7642
rect 19216 7588 19272 7590
rect 19296 7588 19352 7590
rect 19376 7588 19432 7590
rect 19456 7588 19512 7590
rect 26990 7642 27046 7644
rect 27070 7642 27126 7644
rect 27150 7642 27206 7644
rect 27230 7642 27286 7644
rect 26990 7590 27036 7642
rect 27036 7590 27046 7642
rect 27070 7590 27100 7642
rect 27100 7590 27112 7642
rect 27112 7590 27126 7642
rect 27150 7590 27164 7642
rect 27164 7590 27176 7642
rect 27176 7590 27206 7642
rect 27230 7590 27240 7642
rect 27240 7590 27286 7642
rect 26990 7588 27046 7590
rect 27070 7588 27126 7590
rect 27150 7588 27206 7590
rect 27230 7588 27286 7590
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 12102 7098 12158 7100
rect 12182 7098 12238 7100
rect 12262 7098 12318 7100
rect 12342 7098 12398 7100
rect 12102 7046 12148 7098
rect 12148 7046 12158 7098
rect 12182 7046 12212 7098
rect 12212 7046 12224 7098
rect 12224 7046 12238 7098
rect 12262 7046 12276 7098
rect 12276 7046 12288 7098
rect 12288 7046 12318 7098
rect 12342 7046 12352 7098
rect 12352 7046 12398 7098
rect 12102 7044 12158 7046
rect 12182 7044 12238 7046
rect 12262 7044 12318 7046
rect 12342 7044 12398 7046
rect 19876 7098 19932 7100
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 19876 7046 19922 7098
rect 19922 7046 19932 7098
rect 19956 7046 19986 7098
rect 19986 7046 19998 7098
rect 19998 7046 20012 7098
rect 20036 7046 20050 7098
rect 20050 7046 20062 7098
rect 20062 7046 20092 7098
rect 20116 7046 20126 7098
rect 20126 7046 20172 7098
rect 19876 7044 19932 7046
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 27650 7098 27706 7100
rect 27730 7098 27786 7100
rect 27810 7098 27866 7100
rect 27890 7098 27946 7100
rect 27650 7046 27696 7098
rect 27696 7046 27706 7098
rect 27730 7046 27760 7098
rect 27760 7046 27772 7098
rect 27772 7046 27786 7098
rect 27810 7046 27824 7098
rect 27824 7046 27836 7098
rect 27836 7046 27866 7098
rect 27890 7046 27900 7098
rect 27900 7046 27946 7098
rect 27650 7044 27706 7046
rect 27730 7044 27786 7046
rect 27810 7044 27866 7046
rect 27890 7044 27946 7046
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 11442 6554 11498 6556
rect 11522 6554 11578 6556
rect 11602 6554 11658 6556
rect 11682 6554 11738 6556
rect 11442 6502 11488 6554
rect 11488 6502 11498 6554
rect 11522 6502 11552 6554
rect 11552 6502 11564 6554
rect 11564 6502 11578 6554
rect 11602 6502 11616 6554
rect 11616 6502 11628 6554
rect 11628 6502 11658 6554
rect 11682 6502 11692 6554
rect 11692 6502 11738 6554
rect 11442 6500 11498 6502
rect 11522 6500 11578 6502
rect 11602 6500 11658 6502
rect 11682 6500 11738 6502
rect 19216 6554 19272 6556
rect 19296 6554 19352 6556
rect 19376 6554 19432 6556
rect 19456 6554 19512 6556
rect 19216 6502 19262 6554
rect 19262 6502 19272 6554
rect 19296 6502 19326 6554
rect 19326 6502 19338 6554
rect 19338 6502 19352 6554
rect 19376 6502 19390 6554
rect 19390 6502 19402 6554
rect 19402 6502 19432 6554
rect 19456 6502 19466 6554
rect 19466 6502 19512 6554
rect 19216 6500 19272 6502
rect 19296 6500 19352 6502
rect 19376 6500 19432 6502
rect 19456 6500 19512 6502
rect 26990 6554 27046 6556
rect 27070 6554 27126 6556
rect 27150 6554 27206 6556
rect 27230 6554 27286 6556
rect 26990 6502 27036 6554
rect 27036 6502 27046 6554
rect 27070 6502 27100 6554
rect 27100 6502 27112 6554
rect 27112 6502 27126 6554
rect 27150 6502 27164 6554
rect 27164 6502 27176 6554
rect 27176 6502 27206 6554
rect 27230 6502 27240 6554
rect 27240 6502 27286 6554
rect 26990 6500 27046 6502
rect 27070 6500 27126 6502
rect 27150 6500 27206 6502
rect 27230 6500 27286 6502
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 12102 6010 12158 6012
rect 12182 6010 12238 6012
rect 12262 6010 12318 6012
rect 12342 6010 12398 6012
rect 12102 5958 12148 6010
rect 12148 5958 12158 6010
rect 12182 5958 12212 6010
rect 12212 5958 12224 6010
rect 12224 5958 12238 6010
rect 12262 5958 12276 6010
rect 12276 5958 12288 6010
rect 12288 5958 12318 6010
rect 12342 5958 12352 6010
rect 12352 5958 12398 6010
rect 12102 5956 12158 5958
rect 12182 5956 12238 5958
rect 12262 5956 12318 5958
rect 12342 5956 12398 5958
rect 19876 6010 19932 6012
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 19876 5958 19922 6010
rect 19922 5958 19932 6010
rect 19956 5958 19986 6010
rect 19986 5958 19998 6010
rect 19998 5958 20012 6010
rect 20036 5958 20050 6010
rect 20050 5958 20062 6010
rect 20062 5958 20092 6010
rect 20116 5958 20126 6010
rect 20126 5958 20172 6010
rect 19876 5956 19932 5958
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 27650 6010 27706 6012
rect 27730 6010 27786 6012
rect 27810 6010 27866 6012
rect 27890 6010 27946 6012
rect 27650 5958 27696 6010
rect 27696 5958 27706 6010
rect 27730 5958 27760 6010
rect 27760 5958 27772 6010
rect 27772 5958 27786 6010
rect 27810 5958 27824 6010
rect 27824 5958 27836 6010
rect 27836 5958 27866 6010
rect 27890 5958 27900 6010
rect 27900 5958 27946 6010
rect 27650 5956 27706 5958
rect 27730 5956 27786 5958
rect 27810 5956 27866 5958
rect 27890 5956 27946 5958
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 11442 5466 11498 5468
rect 11522 5466 11578 5468
rect 11602 5466 11658 5468
rect 11682 5466 11738 5468
rect 11442 5414 11488 5466
rect 11488 5414 11498 5466
rect 11522 5414 11552 5466
rect 11552 5414 11564 5466
rect 11564 5414 11578 5466
rect 11602 5414 11616 5466
rect 11616 5414 11628 5466
rect 11628 5414 11658 5466
rect 11682 5414 11692 5466
rect 11692 5414 11738 5466
rect 11442 5412 11498 5414
rect 11522 5412 11578 5414
rect 11602 5412 11658 5414
rect 11682 5412 11738 5414
rect 19216 5466 19272 5468
rect 19296 5466 19352 5468
rect 19376 5466 19432 5468
rect 19456 5466 19512 5468
rect 19216 5414 19262 5466
rect 19262 5414 19272 5466
rect 19296 5414 19326 5466
rect 19326 5414 19338 5466
rect 19338 5414 19352 5466
rect 19376 5414 19390 5466
rect 19390 5414 19402 5466
rect 19402 5414 19432 5466
rect 19456 5414 19466 5466
rect 19466 5414 19512 5466
rect 19216 5412 19272 5414
rect 19296 5412 19352 5414
rect 19376 5412 19432 5414
rect 19456 5412 19512 5414
rect 26990 5466 27046 5468
rect 27070 5466 27126 5468
rect 27150 5466 27206 5468
rect 27230 5466 27286 5468
rect 26990 5414 27036 5466
rect 27036 5414 27046 5466
rect 27070 5414 27100 5466
rect 27100 5414 27112 5466
rect 27112 5414 27126 5466
rect 27150 5414 27164 5466
rect 27164 5414 27176 5466
rect 27176 5414 27206 5466
rect 27230 5414 27240 5466
rect 27240 5414 27286 5466
rect 26990 5412 27046 5414
rect 27070 5412 27126 5414
rect 27150 5412 27206 5414
rect 27230 5412 27286 5414
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 12102 4922 12158 4924
rect 12182 4922 12238 4924
rect 12262 4922 12318 4924
rect 12342 4922 12398 4924
rect 12102 4870 12148 4922
rect 12148 4870 12158 4922
rect 12182 4870 12212 4922
rect 12212 4870 12224 4922
rect 12224 4870 12238 4922
rect 12262 4870 12276 4922
rect 12276 4870 12288 4922
rect 12288 4870 12318 4922
rect 12342 4870 12352 4922
rect 12352 4870 12398 4922
rect 12102 4868 12158 4870
rect 12182 4868 12238 4870
rect 12262 4868 12318 4870
rect 12342 4868 12398 4870
rect 19876 4922 19932 4924
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 19876 4870 19922 4922
rect 19922 4870 19932 4922
rect 19956 4870 19986 4922
rect 19986 4870 19998 4922
rect 19998 4870 20012 4922
rect 20036 4870 20050 4922
rect 20050 4870 20062 4922
rect 20062 4870 20092 4922
rect 20116 4870 20126 4922
rect 20126 4870 20172 4922
rect 19876 4868 19932 4870
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 27650 4922 27706 4924
rect 27730 4922 27786 4924
rect 27810 4922 27866 4924
rect 27890 4922 27946 4924
rect 27650 4870 27696 4922
rect 27696 4870 27706 4922
rect 27730 4870 27760 4922
rect 27760 4870 27772 4922
rect 27772 4870 27786 4922
rect 27810 4870 27824 4922
rect 27824 4870 27836 4922
rect 27836 4870 27866 4922
rect 27890 4870 27900 4922
rect 27900 4870 27946 4922
rect 27650 4868 27706 4870
rect 27730 4868 27786 4870
rect 27810 4868 27866 4870
rect 27890 4868 27946 4870
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 11442 4378 11498 4380
rect 11522 4378 11578 4380
rect 11602 4378 11658 4380
rect 11682 4378 11738 4380
rect 11442 4326 11488 4378
rect 11488 4326 11498 4378
rect 11522 4326 11552 4378
rect 11552 4326 11564 4378
rect 11564 4326 11578 4378
rect 11602 4326 11616 4378
rect 11616 4326 11628 4378
rect 11628 4326 11658 4378
rect 11682 4326 11692 4378
rect 11692 4326 11738 4378
rect 11442 4324 11498 4326
rect 11522 4324 11578 4326
rect 11602 4324 11658 4326
rect 11682 4324 11738 4326
rect 19216 4378 19272 4380
rect 19296 4378 19352 4380
rect 19376 4378 19432 4380
rect 19456 4378 19512 4380
rect 19216 4326 19262 4378
rect 19262 4326 19272 4378
rect 19296 4326 19326 4378
rect 19326 4326 19338 4378
rect 19338 4326 19352 4378
rect 19376 4326 19390 4378
rect 19390 4326 19402 4378
rect 19402 4326 19432 4378
rect 19456 4326 19466 4378
rect 19466 4326 19512 4378
rect 19216 4324 19272 4326
rect 19296 4324 19352 4326
rect 19376 4324 19432 4326
rect 19456 4324 19512 4326
rect 26990 4378 27046 4380
rect 27070 4378 27126 4380
rect 27150 4378 27206 4380
rect 27230 4378 27286 4380
rect 26990 4326 27036 4378
rect 27036 4326 27046 4378
rect 27070 4326 27100 4378
rect 27100 4326 27112 4378
rect 27112 4326 27126 4378
rect 27150 4326 27164 4378
rect 27164 4326 27176 4378
rect 27176 4326 27206 4378
rect 27230 4326 27240 4378
rect 27240 4326 27286 4378
rect 26990 4324 27046 4326
rect 27070 4324 27126 4326
rect 27150 4324 27206 4326
rect 27230 4324 27286 4326
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 12102 3834 12158 3836
rect 12182 3834 12238 3836
rect 12262 3834 12318 3836
rect 12342 3834 12398 3836
rect 12102 3782 12148 3834
rect 12148 3782 12158 3834
rect 12182 3782 12212 3834
rect 12212 3782 12224 3834
rect 12224 3782 12238 3834
rect 12262 3782 12276 3834
rect 12276 3782 12288 3834
rect 12288 3782 12318 3834
rect 12342 3782 12352 3834
rect 12352 3782 12398 3834
rect 12102 3780 12158 3782
rect 12182 3780 12238 3782
rect 12262 3780 12318 3782
rect 12342 3780 12398 3782
rect 19876 3834 19932 3836
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 19876 3782 19922 3834
rect 19922 3782 19932 3834
rect 19956 3782 19986 3834
rect 19986 3782 19998 3834
rect 19998 3782 20012 3834
rect 20036 3782 20050 3834
rect 20050 3782 20062 3834
rect 20062 3782 20092 3834
rect 20116 3782 20126 3834
rect 20126 3782 20172 3834
rect 19876 3780 19932 3782
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 27650 3834 27706 3836
rect 27730 3834 27786 3836
rect 27810 3834 27866 3836
rect 27890 3834 27946 3836
rect 27650 3782 27696 3834
rect 27696 3782 27706 3834
rect 27730 3782 27760 3834
rect 27760 3782 27772 3834
rect 27772 3782 27786 3834
rect 27810 3782 27824 3834
rect 27824 3782 27836 3834
rect 27836 3782 27866 3834
rect 27890 3782 27900 3834
rect 27900 3782 27946 3834
rect 27650 3780 27706 3782
rect 27730 3780 27786 3782
rect 27810 3780 27866 3782
rect 27890 3780 27946 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 11442 3290 11498 3292
rect 11522 3290 11578 3292
rect 11602 3290 11658 3292
rect 11682 3290 11738 3292
rect 11442 3238 11488 3290
rect 11488 3238 11498 3290
rect 11522 3238 11552 3290
rect 11552 3238 11564 3290
rect 11564 3238 11578 3290
rect 11602 3238 11616 3290
rect 11616 3238 11628 3290
rect 11628 3238 11658 3290
rect 11682 3238 11692 3290
rect 11692 3238 11738 3290
rect 11442 3236 11498 3238
rect 11522 3236 11578 3238
rect 11602 3236 11658 3238
rect 11682 3236 11738 3238
rect 19216 3290 19272 3292
rect 19296 3290 19352 3292
rect 19376 3290 19432 3292
rect 19456 3290 19512 3292
rect 19216 3238 19262 3290
rect 19262 3238 19272 3290
rect 19296 3238 19326 3290
rect 19326 3238 19338 3290
rect 19338 3238 19352 3290
rect 19376 3238 19390 3290
rect 19390 3238 19402 3290
rect 19402 3238 19432 3290
rect 19456 3238 19466 3290
rect 19466 3238 19512 3290
rect 19216 3236 19272 3238
rect 19296 3236 19352 3238
rect 19376 3236 19432 3238
rect 19456 3236 19512 3238
rect 26990 3290 27046 3292
rect 27070 3290 27126 3292
rect 27150 3290 27206 3292
rect 27230 3290 27286 3292
rect 26990 3238 27036 3290
rect 27036 3238 27046 3290
rect 27070 3238 27100 3290
rect 27100 3238 27112 3290
rect 27112 3238 27126 3290
rect 27150 3238 27164 3290
rect 27164 3238 27176 3290
rect 27176 3238 27206 3290
rect 27230 3238 27240 3290
rect 27240 3238 27286 3290
rect 26990 3236 27046 3238
rect 27070 3236 27126 3238
rect 27150 3236 27206 3238
rect 27230 3236 27286 3238
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 12102 2746 12158 2748
rect 12182 2746 12238 2748
rect 12262 2746 12318 2748
rect 12342 2746 12398 2748
rect 12102 2694 12148 2746
rect 12148 2694 12158 2746
rect 12182 2694 12212 2746
rect 12212 2694 12224 2746
rect 12224 2694 12238 2746
rect 12262 2694 12276 2746
rect 12276 2694 12288 2746
rect 12288 2694 12318 2746
rect 12342 2694 12352 2746
rect 12352 2694 12398 2746
rect 12102 2692 12158 2694
rect 12182 2692 12238 2694
rect 12262 2692 12318 2694
rect 12342 2692 12398 2694
rect 19876 2746 19932 2748
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 19876 2694 19922 2746
rect 19922 2694 19932 2746
rect 19956 2694 19986 2746
rect 19986 2694 19998 2746
rect 19998 2694 20012 2746
rect 20036 2694 20050 2746
rect 20050 2694 20062 2746
rect 20062 2694 20092 2746
rect 20116 2694 20126 2746
rect 20126 2694 20172 2746
rect 19876 2692 19932 2694
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 27650 2746 27706 2748
rect 27730 2746 27786 2748
rect 27810 2746 27866 2748
rect 27890 2746 27946 2748
rect 27650 2694 27696 2746
rect 27696 2694 27706 2746
rect 27730 2694 27760 2746
rect 27760 2694 27772 2746
rect 27772 2694 27786 2746
rect 27810 2694 27824 2746
rect 27824 2694 27836 2746
rect 27836 2694 27866 2746
rect 27890 2694 27900 2746
rect 27900 2694 27946 2746
rect 27650 2692 27706 2694
rect 27730 2692 27786 2694
rect 27810 2692 27866 2694
rect 27890 2692 27946 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 11442 2202 11498 2204
rect 11522 2202 11578 2204
rect 11602 2202 11658 2204
rect 11682 2202 11738 2204
rect 11442 2150 11488 2202
rect 11488 2150 11498 2202
rect 11522 2150 11552 2202
rect 11552 2150 11564 2202
rect 11564 2150 11578 2202
rect 11602 2150 11616 2202
rect 11616 2150 11628 2202
rect 11628 2150 11658 2202
rect 11682 2150 11692 2202
rect 11692 2150 11738 2202
rect 11442 2148 11498 2150
rect 11522 2148 11578 2150
rect 11602 2148 11658 2150
rect 11682 2148 11738 2150
rect 19216 2202 19272 2204
rect 19296 2202 19352 2204
rect 19376 2202 19432 2204
rect 19456 2202 19512 2204
rect 19216 2150 19262 2202
rect 19262 2150 19272 2202
rect 19296 2150 19326 2202
rect 19326 2150 19338 2202
rect 19338 2150 19352 2202
rect 19376 2150 19390 2202
rect 19390 2150 19402 2202
rect 19402 2150 19432 2202
rect 19456 2150 19466 2202
rect 19466 2150 19512 2202
rect 19216 2148 19272 2150
rect 19296 2148 19352 2150
rect 19376 2148 19432 2150
rect 19456 2148 19512 2150
rect 26990 2202 27046 2204
rect 27070 2202 27126 2204
rect 27150 2202 27206 2204
rect 27230 2202 27286 2204
rect 26990 2150 27036 2202
rect 27036 2150 27046 2202
rect 27070 2150 27100 2202
rect 27100 2150 27112 2202
rect 27112 2150 27126 2202
rect 27150 2150 27164 2202
rect 27164 2150 27176 2202
rect 27176 2150 27206 2202
rect 27230 2150 27240 2202
rect 27240 2150 27286 2202
rect 26990 2148 27046 2150
rect 27070 2148 27126 2150
rect 27150 2148 27206 2150
rect 27230 2148 27286 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 12102 1658 12158 1660
rect 12182 1658 12238 1660
rect 12262 1658 12318 1660
rect 12342 1658 12398 1660
rect 12102 1606 12148 1658
rect 12148 1606 12158 1658
rect 12182 1606 12212 1658
rect 12212 1606 12224 1658
rect 12224 1606 12238 1658
rect 12262 1606 12276 1658
rect 12276 1606 12288 1658
rect 12288 1606 12318 1658
rect 12342 1606 12352 1658
rect 12352 1606 12398 1658
rect 12102 1604 12158 1606
rect 12182 1604 12238 1606
rect 12262 1604 12318 1606
rect 12342 1604 12398 1606
rect 19876 1658 19932 1660
rect 19956 1658 20012 1660
rect 20036 1658 20092 1660
rect 20116 1658 20172 1660
rect 19876 1606 19922 1658
rect 19922 1606 19932 1658
rect 19956 1606 19986 1658
rect 19986 1606 19998 1658
rect 19998 1606 20012 1658
rect 20036 1606 20050 1658
rect 20050 1606 20062 1658
rect 20062 1606 20092 1658
rect 20116 1606 20126 1658
rect 20126 1606 20172 1658
rect 19876 1604 19932 1606
rect 19956 1604 20012 1606
rect 20036 1604 20092 1606
rect 20116 1604 20172 1606
rect 27650 1658 27706 1660
rect 27730 1658 27786 1660
rect 27810 1658 27866 1660
rect 27890 1658 27946 1660
rect 27650 1606 27696 1658
rect 27696 1606 27706 1658
rect 27730 1606 27760 1658
rect 27760 1606 27772 1658
rect 27772 1606 27786 1658
rect 27810 1606 27824 1658
rect 27824 1606 27836 1658
rect 27836 1606 27866 1658
rect 27890 1606 27900 1658
rect 27900 1606 27946 1658
rect 27650 1604 27706 1606
rect 27730 1604 27786 1606
rect 27810 1604 27866 1606
rect 27890 1604 27946 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 11442 1114 11498 1116
rect 11522 1114 11578 1116
rect 11602 1114 11658 1116
rect 11682 1114 11738 1116
rect 11442 1062 11488 1114
rect 11488 1062 11498 1114
rect 11522 1062 11552 1114
rect 11552 1062 11564 1114
rect 11564 1062 11578 1114
rect 11602 1062 11616 1114
rect 11616 1062 11628 1114
rect 11628 1062 11658 1114
rect 11682 1062 11692 1114
rect 11692 1062 11738 1114
rect 11442 1060 11498 1062
rect 11522 1060 11578 1062
rect 11602 1060 11658 1062
rect 11682 1060 11738 1062
rect 19216 1114 19272 1116
rect 19296 1114 19352 1116
rect 19376 1114 19432 1116
rect 19456 1114 19512 1116
rect 19216 1062 19262 1114
rect 19262 1062 19272 1114
rect 19296 1062 19326 1114
rect 19326 1062 19338 1114
rect 19338 1062 19352 1114
rect 19376 1062 19390 1114
rect 19390 1062 19402 1114
rect 19402 1062 19432 1114
rect 19456 1062 19466 1114
rect 19466 1062 19512 1114
rect 19216 1060 19272 1062
rect 19296 1060 19352 1062
rect 19376 1060 19432 1062
rect 19456 1060 19512 1062
rect 26990 1114 27046 1116
rect 27070 1114 27126 1116
rect 27150 1114 27206 1116
rect 27230 1114 27286 1116
rect 26990 1062 27036 1114
rect 27036 1062 27046 1114
rect 27070 1062 27100 1114
rect 27100 1062 27112 1114
rect 27112 1062 27126 1114
rect 27150 1062 27164 1114
rect 27164 1062 27176 1114
rect 27176 1062 27206 1114
rect 27230 1062 27240 1114
rect 27240 1062 27286 1114
rect 26990 1060 27046 1062
rect 27070 1060 27126 1062
rect 27150 1060 27206 1062
rect 27230 1060 27286 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 12102 570 12158 572
rect 12182 570 12238 572
rect 12262 570 12318 572
rect 12342 570 12398 572
rect 12102 518 12148 570
rect 12148 518 12158 570
rect 12182 518 12212 570
rect 12212 518 12224 570
rect 12224 518 12238 570
rect 12262 518 12276 570
rect 12276 518 12288 570
rect 12288 518 12318 570
rect 12342 518 12352 570
rect 12352 518 12398 570
rect 12102 516 12158 518
rect 12182 516 12238 518
rect 12262 516 12318 518
rect 12342 516 12398 518
rect 19876 570 19932 572
rect 19956 570 20012 572
rect 20036 570 20092 572
rect 20116 570 20172 572
rect 19876 518 19922 570
rect 19922 518 19932 570
rect 19956 518 19986 570
rect 19986 518 19998 570
rect 19998 518 20012 570
rect 20036 518 20050 570
rect 20050 518 20062 570
rect 20062 518 20092 570
rect 20116 518 20126 570
rect 20126 518 20172 570
rect 19876 516 19932 518
rect 19956 516 20012 518
rect 20036 516 20092 518
rect 20116 516 20172 518
rect 27650 570 27706 572
rect 27730 570 27786 572
rect 27810 570 27866 572
rect 27890 570 27946 572
rect 27650 518 27696 570
rect 27696 518 27706 570
rect 27730 518 27760 570
rect 27760 518 27772 570
rect 27772 518 27786 570
rect 27810 518 27824 570
rect 27824 518 27836 570
rect 27836 518 27866 570
rect 27890 518 27900 570
rect 27900 518 27946 570
rect 27650 516 27706 518
rect 27730 516 27786 518
rect 27810 516 27866 518
rect 27890 516 27946 518
<< metal3 >>
rect 11646 44780 11652 44844
rect 11716 44842 11722 44844
rect 11789 44842 11855 44845
rect 11716 44840 11855 44842
rect 11716 44784 11794 44840
rect 11850 44784 11855 44840
rect 11716 44782 11855 44784
rect 11716 44780 11722 44782
rect 11789 44779 11855 44782
rect 12198 44780 12204 44844
rect 12268 44842 12274 44844
rect 13077 44842 13143 44845
rect 21633 44844 21699 44845
rect 21582 44842 21588 44844
rect 12268 44840 13143 44842
rect 12268 44784 13082 44840
rect 13138 44784 13143 44840
rect 12268 44782 13143 44784
rect 21542 44782 21588 44842
rect 21652 44840 21699 44844
rect 21694 44784 21699 44840
rect 12268 44780 12274 44782
rect 13077 44779 13143 44782
rect 21582 44780 21588 44782
rect 21652 44780 21699 44784
rect 27102 44780 27108 44844
rect 27172 44842 27178 44844
rect 27429 44842 27495 44845
rect 27172 44840 27495 44842
rect 27172 44784 27434 44840
rect 27490 44784 27495 44840
rect 27172 44782 27495 44784
rect 27172 44780 27178 44782
rect 21633 44779 21699 44780
rect 27429 44779 27495 44782
rect 27654 44780 27660 44844
rect 27724 44842 27730 44844
rect 28165 44842 28231 44845
rect 27724 44840 28231 44842
rect 27724 44784 28170 44840
rect 28226 44784 28231 44840
rect 27724 44782 28231 44784
rect 27724 44780 27730 44782
rect 28165 44779 28231 44782
rect 23790 44644 23796 44708
rect 23860 44706 23866 44708
rect 24025 44706 24091 44709
rect 24393 44708 24459 44709
rect 24945 44708 25011 44709
rect 25497 44708 25563 44709
rect 26049 44708 26115 44709
rect 24342 44706 24348 44708
rect 23860 44704 24091 44706
rect 23860 44648 24030 44704
rect 24086 44648 24091 44704
rect 23860 44646 24091 44648
rect 24302 44646 24348 44706
rect 24412 44704 24459 44708
rect 24894 44706 24900 44708
rect 24454 44648 24459 44704
rect 23860 44644 23866 44646
rect 24025 44643 24091 44646
rect 24342 44644 24348 44646
rect 24412 44644 24459 44648
rect 24854 44646 24900 44706
rect 24964 44704 25011 44708
rect 25446 44706 25452 44708
rect 25006 44648 25011 44704
rect 24894 44644 24900 44646
rect 24964 44644 25011 44648
rect 25406 44646 25452 44706
rect 25516 44704 25563 44708
rect 25998 44706 26004 44708
rect 25558 44648 25563 44704
rect 25446 44644 25452 44646
rect 25516 44644 25563 44648
rect 25958 44646 26004 44706
rect 26068 44704 26115 44708
rect 26110 44648 26115 44704
rect 25998 44644 26004 44646
rect 26068 44644 26115 44648
rect 24393 44643 24459 44644
rect 24945 44643 25011 44644
rect 25497 44643 25563 44644
rect 26049 44643 26115 44644
rect 26509 44708 26575 44709
rect 26509 44704 26556 44708
rect 26620 44706 26626 44708
rect 26509 44648 26514 44704
rect 26509 44644 26556 44648
rect 26620 44646 26666 44706
rect 26620 44644 26626 44646
rect 28206 44644 28212 44708
rect 28276 44706 28282 44708
rect 28993 44706 29059 44709
rect 28276 44704 29059 44706
rect 28276 44648 28998 44704
rect 29054 44648 29059 44704
rect 28276 44646 29059 44648
rect 28276 44644 28282 44646
rect 26509 44643 26575 44644
rect 28993 44643 29059 44646
rect 3658 44640 3974 44641
rect 3658 44576 3664 44640
rect 3728 44576 3744 44640
rect 3808 44576 3824 44640
rect 3888 44576 3904 44640
rect 3968 44576 3974 44640
rect 3658 44575 3974 44576
rect 11432 44640 11748 44641
rect 11432 44576 11438 44640
rect 11502 44576 11518 44640
rect 11582 44576 11598 44640
rect 11662 44576 11678 44640
rect 11742 44576 11748 44640
rect 11432 44575 11748 44576
rect 19206 44640 19522 44641
rect 19206 44576 19212 44640
rect 19276 44576 19292 44640
rect 19356 44576 19372 44640
rect 19436 44576 19452 44640
rect 19516 44576 19522 44640
rect 19206 44575 19522 44576
rect 26980 44640 27296 44641
rect 26980 44576 26986 44640
rect 27050 44576 27066 44640
rect 27130 44576 27146 44640
rect 27210 44576 27226 44640
rect 27290 44576 27296 44640
rect 26980 44575 27296 44576
rect 7189 44572 7255 44573
rect 7189 44570 7236 44572
rect 7144 44568 7236 44570
rect 7144 44512 7194 44568
rect 7144 44510 7236 44512
rect 7189 44508 7236 44510
rect 7300 44508 7306 44572
rect 7649 44570 7715 44573
rect 8293 44572 8359 44573
rect 7782 44570 7788 44572
rect 7649 44568 7788 44570
rect 7649 44512 7654 44568
rect 7710 44512 7788 44568
rect 7649 44510 7788 44512
rect 7189 44507 7255 44508
rect 7649 44507 7715 44510
rect 7782 44508 7788 44510
rect 7852 44508 7858 44572
rect 8293 44570 8340 44572
rect 8248 44568 8340 44570
rect 8248 44512 8298 44568
rect 8248 44510 8340 44512
rect 8293 44508 8340 44510
rect 8404 44508 8410 44572
rect 8753 44570 8819 44573
rect 8886 44570 8892 44572
rect 8753 44568 8892 44570
rect 8753 44512 8758 44568
rect 8814 44512 8892 44568
rect 8753 44510 8892 44512
rect 8293 44507 8359 44508
rect 8753 44507 8819 44510
rect 8886 44508 8892 44510
rect 8956 44508 8962 44572
rect 9305 44570 9371 44573
rect 12801 44572 12867 44573
rect 9438 44570 9444 44572
rect 9305 44568 9444 44570
rect 9305 44512 9310 44568
rect 9366 44512 9444 44568
rect 9305 44510 9444 44512
rect 9305 44507 9371 44510
rect 9438 44508 9444 44510
rect 9508 44508 9514 44572
rect 12750 44508 12756 44572
rect 12820 44570 12867 44572
rect 12820 44568 12912 44570
rect 12862 44512 12912 44568
rect 12820 44510 12912 44512
rect 12820 44508 12867 44510
rect 12801 44507 12867 44508
rect 4318 44096 4634 44097
rect 4318 44032 4324 44096
rect 4388 44032 4404 44096
rect 4468 44032 4484 44096
rect 4548 44032 4564 44096
rect 4628 44032 4634 44096
rect 4318 44031 4634 44032
rect 12092 44096 12408 44097
rect 12092 44032 12098 44096
rect 12162 44032 12178 44096
rect 12242 44032 12258 44096
rect 12322 44032 12338 44096
rect 12402 44032 12408 44096
rect 12092 44031 12408 44032
rect 19866 44096 20182 44097
rect 19866 44032 19872 44096
rect 19936 44032 19952 44096
rect 20016 44032 20032 44096
rect 20096 44032 20112 44096
rect 20176 44032 20182 44096
rect 19866 44031 20182 44032
rect 27640 44096 27956 44097
rect 27640 44032 27646 44096
rect 27710 44032 27726 44096
rect 27790 44032 27806 44096
rect 27870 44032 27886 44096
rect 27950 44032 27956 44096
rect 27640 44031 27956 44032
rect 6126 43964 6132 44028
rect 6196 44026 6202 44028
rect 6545 44026 6611 44029
rect 6196 44024 6611 44026
rect 6196 43968 6550 44024
rect 6606 43968 6611 44024
rect 6196 43966 6611 43968
rect 6196 43964 6202 43966
rect 6545 43963 6611 43966
rect 6678 43964 6684 44028
rect 6748 44026 6754 44028
rect 6913 44026 6979 44029
rect 6748 44024 6979 44026
rect 6748 43968 6918 44024
rect 6974 43968 6979 44024
rect 6748 43966 6979 43968
rect 6748 43964 6754 43966
rect 6913 43963 6979 43966
rect 9990 43964 9996 44028
rect 10060 44026 10066 44028
rect 10685 44026 10751 44029
rect 13261 44028 13327 44029
rect 16573 44028 16639 44029
rect 13261 44026 13308 44028
rect 10060 44024 10751 44026
rect 10060 43968 10690 44024
rect 10746 43968 10751 44024
rect 10060 43966 10751 43968
rect 13216 44024 13308 44026
rect 13216 43968 13266 44024
rect 13216 43966 13308 43968
rect 10060 43964 10066 43966
rect 10685 43963 10751 43966
rect 13261 43964 13308 43966
rect 13372 43964 13378 44028
rect 16573 44026 16620 44028
rect 16528 44024 16620 44026
rect 16528 43968 16578 44024
rect 16528 43966 16620 43968
rect 16573 43964 16620 43966
rect 16684 43964 16690 44028
rect 17166 43964 17172 44028
rect 17236 44026 17242 44028
rect 17401 44026 17467 44029
rect 18137 44026 18203 44029
rect 17236 44024 18203 44026
rect 17236 43968 17406 44024
rect 17462 43968 18142 44024
rect 18198 43968 18203 44024
rect 17236 43966 18203 43968
rect 17236 43964 17242 43966
rect 13261 43963 13327 43964
rect 16573 43963 16639 43964
rect 17401 43963 17467 43966
rect 18137 43963 18203 43966
rect 11094 43828 11100 43892
rect 11164 43890 11170 43892
rect 11329 43890 11395 43893
rect 11164 43888 11395 43890
rect 11164 43832 11334 43888
rect 11390 43832 11395 43888
rect 11164 43830 11395 43832
rect 11164 43828 11170 43830
rect 11329 43827 11395 43830
rect 13813 43756 13879 43757
rect 13813 43754 13860 43756
rect 13768 43752 13860 43754
rect 13768 43696 13818 43752
rect 13768 43694 13860 43696
rect 13813 43692 13860 43694
rect 13924 43692 13930 43756
rect 13813 43691 13879 43692
rect 3658 43552 3974 43553
rect 3658 43488 3664 43552
rect 3728 43488 3744 43552
rect 3808 43488 3824 43552
rect 3888 43488 3904 43552
rect 3968 43488 3974 43552
rect 3658 43487 3974 43488
rect 11432 43552 11748 43553
rect 11432 43488 11438 43552
rect 11502 43488 11518 43552
rect 11582 43488 11598 43552
rect 11662 43488 11678 43552
rect 11742 43488 11748 43552
rect 11432 43487 11748 43488
rect 19206 43552 19522 43553
rect 19206 43488 19212 43552
rect 19276 43488 19292 43552
rect 19356 43488 19372 43552
rect 19436 43488 19452 43552
rect 19516 43488 19522 43552
rect 19206 43487 19522 43488
rect 26980 43552 27296 43553
rect 26980 43488 26986 43552
rect 27050 43488 27066 43552
rect 27130 43488 27146 43552
rect 27210 43488 27226 43552
rect 27290 43488 27296 43552
rect 26980 43487 27296 43488
rect 14365 43484 14431 43485
rect 14365 43482 14412 43484
rect 14320 43480 14412 43482
rect 14320 43424 14370 43480
rect 14320 43422 14412 43424
rect 14365 43420 14412 43422
rect 14476 43420 14482 43484
rect 14365 43419 14431 43420
rect 18822 43284 18828 43348
rect 18892 43346 18898 43348
rect 19609 43346 19675 43349
rect 18892 43344 19675 43346
rect 18892 43288 19614 43344
rect 19670 43288 19675 43344
rect 18892 43286 19675 43288
rect 18892 43284 18898 43286
rect 19609 43283 19675 43286
rect 14958 43148 14964 43212
rect 15028 43210 15034 43212
rect 15101 43210 15167 43213
rect 15028 43208 15167 43210
rect 15028 43152 15106 43208
rect 15162 43152 15167 43208
rect 15028 43150 15167 43152
rect 15028 43148 15034 43150
rect 15101 43147 15167 43150
rect 18270 43148 18276 43212
rect 18340 43210 18346 43212
rect 19149 43210 19215 43213
rect 18340 43208 19215 43210
rect 18340 43152 19154 43208
rect 19210 43152 19215 43208
rect 18340 43150 19215 43152
rect 18340 43148 18346 43150
rect 19149 43147 19215 43150
rect 4318 43008 4634 43009
rect 4318 42944 4324 43008
rect 4388 42944 4404 43008
rect 4468 42944 4484 43008
rect 4548 42944 4564 43008
rect 4628 42944 4634 43008
rect 4318 42943 4634 42944
rect 12092 43008 12408 43009
rect 12092 42944 12098 43008
rect 12162 42944 12178 43008
rect 12242 42944 12258 43008
rect 12322 42944 12338 43008
rect 12402 42944 12408 43008
rect 12092 42943 12408 42944
rect 19866 43008 20182 43009
rect 19866 42944 19872 43008
rect 19936 42944 19952 43008
rect 20016 42944 20032 43008
rect 20096 42944 20112 43008
rect 20176 42944 20182 43008
rect 19866 42943 20182 42944
rect 27640 43008 27956 43009
rect 27640 42944 27646 43008
rect 27710 42944 27726 43008
rect 27790 42944 27806 43008
rect 27870 42944 27886 43008
rect 27950 42944 27956 43008
rect 27640 42943 27956 42944
rect 15469 42940 15535 42941
rect 15469 42938 15516 42940
rect 15424 42936 15516 42938
rect 15424 42880 15474 42936
rect 15424 42878 15516 42880
rect 15469 42876 15516 42878
rect 15580 42876 15586 42940
rect 17718 42876 17724 42940
rect 17788 42938 17794 42940
rect 17953 42938 18019 42941
rect 17788 42936 18019 42938
rect 17788 42880 17958 42936
rect 18014 42880 18019 42936
rect 17788 42878 18019 42880
rect 17788 42876 17794 42878
rect 15469 42875 15535 42876
rect 17953 42875 18019 42878
rect 3658 42464 3974 42465
rect 3658 42400 3664 42464
rect 3728 42400 3744 42464
rect 3808 42400 3824 42464
rect 3888 42400 3904 42464
rect 3968 42400 3974 42464
rect 3658 42399 3974 42400
rect 11432 42464 11748 42465
rect 11432 42400 11438 42464
rect 11502 42400 11518 42464
rect 11582 42400 11598 42464
rect 11662 42400 11678 42464
rect 11742 42400 11748 42464
rect 11432 42399 11748 42400
rect 19206 42464 19522 42465
rect 19206 42400 19212 42464
rect 19276 42400 19292 42464
rect 19356 42400 19372 42464
rect 19436 42400 19452 42464
rect 19516 42400 19522 42464
rect 19206 42399 19522 42400
rect 26980 42464 27296 42465
rect 26980 42400 26986 42464
rect 27050 42400 27066 42464
rect 27130 42400 27146 42464
rect 27210 42400 27226 42464
rect 27290 42400 27296 42464
rect 26980 42399 27296 42400
rect 17401 42258 17467 42261
rect 18321 42258 18387 42261
rect 19149 42258 19215 42261
rect 23657 42260 23723 42261
rect 17401 42256 19215 42258
rect 17401 42200 17406 42256
rect 17462 42200 18326 42256
rect 18382 42200 19154 42256
rect 19210 42200 19215 42256
rect 17401 42198 19215 42200
rect 17401 42195 17467 42198
rect 18321 42195 18387 42198
rect 19149 42195 19215 42198
rect 23606 42196 23612 42260
rect 23676 42258 23723 42260
rect 23676 42256 23768 42258
rect 23718 42200 23768 42256
rect 23676 42198 23768 42200
rect 23676 42196 23723 42198
rect 23657 42195 23723 42196
rect 4318 41920 4634 41921
rect 4318 41856 4324 41920
rect 4388 41856 4404 41920
rect 4468 41856 4484 41920
rect 4548 41856 4564 41920
rect 4628 41856 4634 41920
rect 4318 41855 4634 41856
rect 12092 41920 12408 41921
rect 12092 41856 12098 41920
rect 12162 41856 12178 41920
rect 12242 41856 12258 41920
rect 12322 41856 12338 41920
rect 12402 41856 12408 41920
rect 12092 41855 12408 41856
rect 19866 41920 20182 41921
rect 19866 41856 19872 41920
rect 19936 41856 19952 41920
rect 20016 41856 20032 41920
rect 20096 41856 20112 41920
rect 20176 41856 20182 41920
rect 19866 41855 20182 41856
rect 27640 41920 27956 41921
rect 27640 41856 27646 41920
rect 27710 41856 27726 41920
rect 27790 41856 27806 41920
rect 27870 41856 27886 41920
rect 27950 41856 27956 41920
rect 27640 41855 27956 41856
rect 13721 41852 13787 41853
rect 13670 41850 13676 41852
rect 13630 41790 13676 41850
rect 13740 41848 13787 41852
rect 13782 41792 13787 41848
rect 13670 41788 13676 41790
rect 13740 41788 13787 41792
rect 13721 41787 13787 41788
rect 23933 41578 23999 41581
rect 24526 41578 24532 41580
rect 23933 41576 24532 41578
rect 23933 41520 23938 41576
rect 23994 41520 24532 41576
rect 23933 41518 24532 41520
rect 23933 41515 23999 41518
rect 24526 41516 24532 41518
rect 24596 41516 24602 41580
rect 3658 41376 3974 41377
rect 3658 41312 3664 41376
rect 3728 41312 3744 41376
rect 3808 41312 3824 41376
rect 3888 41312 3904 41376
rect 3968 41312 3974 41376
rect 3658 41311 3974 41312
rect 11432 41376 11748 41377
rect 11432 41312 11438 41376
rect 11502 41312 11518 41376
rect 11582 41312 11598 41376
rect 11662 41312 11678 41376
rect 11742 41312 11748 41376
rect 11432 41311 11748 41312
rect 19206 41376 19522 41377
rect 19206 41312 19212 41376
rect 19276 41312 19292 41376
rect 19356 41312 19372 41376
rect 19436 41312 19452 41376
rect 19516 41312 19522 41376
rect 19206 41311 19522 41312
rect 26980 41376 27296 41377
rect 26980 41312 26986 41376
rect 27050 41312 27066 41376
rect 27130 41312 27146 41376
rect 27210 41312 27226 41376
rect 27290 41312 27296 41376
rect 26980 41311 27296 41312
rect 16062 41108 16068 41172
rect 16132 41170 16138 41172
rect 16297 41170 16363 41173
rect 16132 41168 16363 41170
rect 16132 41112 16302 41168
rect 16358 41112 16363 41168
rect 16132 41110 16363 41112
rect 16132 41108 16138 41110
rect 16297 41107 16363 41110
rect 4318 40832 4634 40833
rect 4318 40768 4324 40832
rect 4388 40768 4404 40832
rect 4468 40768 4484 40832
rect 4548 40768 4564 40832
rect 4628 40768 4634 40832
rect 4318 40767 4634 40768
rect 12092 40832 12408 40833
rect 12092 40768 12098 40832
rect 12162 40768 12178 40832
rect 12242 40768 12258 40832
rect 12322 40768 12338 40832
rect 12402 40768 12408 40832
rect 12092 40767 12408 40768
rect 19866 40832 20182 40833
rect 19866 40768 19872 40832
rect 19936 40768 19952 40832
rect 20016 40768 20032 40832
rect 20096 40768 20112 40832
rect 20176 40768 20182 40832
rect 19866 40767 20182 40768
rect 27640 40832 27956 40833
rect 27640 40768 27646 40832
rect 27710 40768 27726 40832
rect 27790 40768 27806 40832
rect 27870 40768 27886 40832
rect 27950 40768 27956 40832
rect 27640 40767 27956 40768
rect 3658 40288 3974 40289
rect 3658 40224 3664 40288
rect 3728 40224 3744 40288
rect 3808 40224 3824 40288
rect 3888 40224 3904 40288
rect 3968 40224 3974 40288
rect 3658 40223 3974 40224
rect 11432 40288 11748 40289
rect 11432 40224 11438 40288
rect 11502 40224 11518 40288
rect 11582 40224 11598 40288
rect 11662 40224 11678 40288
rect 11742 40224 11748 40288
rect 11432 40223 11748 40224
rect 19206 40288 19522 40289
rect 19206 40224 19212 40288
rect 19276 40224 19292 40288
rect 19356 40224 19372 40288
rect 19436 40224 19452 40288
rect 19516 40224 19522 40288
rect 19206 40223 19522 40224
rect 26980 40288 27296 40289
rect 26980 40224 26986 40288
rect 27050 40224 27066 40288
rect 27130 40224 27146 40288
rect 27210 40224 27226 40288
rect 27290 40224 27296 40288
rect 26980 40223 27296 40224
rect 10961 39946 11027 39949
rect 12985 39946 13051 39949
rect 10961 39944 13051 39946
rect 10961 39888 10966 39944
rect 11022 39888 12990 39944
rect 13046 39888 13051 39944
rect 10961 39886 13051 39888
rect 10961 39883 11027 39886
rect 12985 39883 13051 39886
rect 4318 39744 4634 39745
rect 4318 39680 4324 39744
rect 4388 39680 4404 39744
rect 4468 39680 4484 39744
rect 4548 39680 4564 39744
rect 4628 39680 4634 39744
rect 4318 39679 4634 39680
rect 12092 39744 12408 39745
rect 12092 39680 12098 39744
rect 12162 39680 12178 39744
rect 12242 39680 12258 39744
rect 12322 39680 12338 39744
rect 12402 39680 12408 39744
rect 12092 39679 12408 39680
rect 19866 39744 20182 39745
rect 19866 39680 19872 39744
rect 19936 39680 19952 39744
rect 20016 39680 20032 39744
rect 20096 39680 20112 39744
rect 20176 39680 20182 39744
rect 19866 39679 20182 39680
rect 27640 39744 27956 39745
rect 27640 39680 27646 39744
rect 27710 39680 27726 39744
rect 27790 39680 27806 39744
rect 27870 39680 27886 39744
rect 27950 39680 27956 39744
rect 27640 39679 27956 39680
rect 20345 39402 20411 39405
rect 20478 39402 20484 39404
rect 20345 39400 20484 39402
rect 20345 39344 20350 39400
rect 20406 39344 20484 39400
rect 20345 39342 20484 39344
rect 20345 39339 20411 39342
rect 20478 39340 20484 39342
rect 20548 39340 20554 39404
rect 3658 39200 3974 39201
rect 3658 39136 3664 39200
rect 3728 39136 3744 39200
rect 3808 39136 3824 39200
rect 3888 39136 3904 39200
rect 3968 39136 3974 39200
rect 3658 39135 3974 39136
rect 11432 39200 11748 39201
rect 11432 39136 11438 39200
rect 11502 39136 11518 39200
rect 11582 39136 11598 39200
rect 11662 39136 11678 39200
rect 11742 39136 11748 39200
rect 11432 39135 11748 39136
rect 19206 39200 19522 39201
rect 19206 39136 19212 39200
rect 19276 39136 19292 39200
rect 19356 39136 19372 39200
rect 19436 39136 19452 39200
rect 19516 39136 19522 39200
rect 19206 39135 19522 39136
rect 26980 39200 27296 39201
rect 26980 39136 26986 39200
rect 27050 39136 27066 39200
rect 27130 39136 27146 39200
rect 27210 39136 27226 39200
rect 27290 39136 27296 39200
rect 26980 39135 27296 39136
rect 25865 38994 25931 38997
rect 27705 38994 27771 38997
rect 25865 38992 27771 38994
rect 25865 38936 25870 38992
rect 25926 38936 27710 38992
rect 27766 38936 27771 38992
rect 25865 38934 27771 38936
rect 25865 38931 25931 38934
rect 27705 38931 27771 38934
rect 20161 38858 20227 38861
rect 20294 38858 20300 38860
rect 20161 38856 20300 38858
rect 20161 38800 20166 38856
rect 20222 38800 20300 38856
rect 20161 38798 20300 38800
rect 20161 38795 20227 38798
rect 20294 38796 20300 38798
rect 20364 38796 20370 38860
rect 4318 38656 4634 38657
rect 4318 38592 4324 38656
rect 4388 38592 4404 38656
rect 4468 38592 4484 38656
rect 4548 38592 4564 38656
rect 4628 38592 4634 38656
rect 4318 38591 4634 38592
rect 12092 38656 12408 38657
rect 12092 38592 12098 38656
rect 12162 38592 12178 38656
rect 12242 38592 12258 38656
rect 12322 38592 12338 38656
rect 12402 38592 12408 38656
rect 12092 38591 12408 38592
rect 19866 38656 20182 38657
rect 19866 38592 19872 38656
rect 19936 38592 19952 38656
rect 20016 38592 20032 38656
rect 20096 38592 20112 38656
rect 20176 38592 20182 38656
rect 19866 38591 20182 38592
rect 27640 38656 27956 38657
rect 27640 38592 27646 38656
rect 27710 38592 27726 38656
rect 27790 38592 27806 38656
rect 27870 38592 27886 38656
rect 27950 38592 27956 38656
rect 27640 38591 27956 38592
rect 19609 38450 19675 38453
rect 20161 38450 20227 38453
rect 19609 38448 20227 38450
rect 19609 38392 19614 38448
rect 19670 38392 20166 38448
rect 20222 38392 20227 38448
rect 19609 38390 20227 38392
rect 19609 38387 19675 38390
rect 20161 38387 20227 38390
rect 19425 38314 19491 38317
rect 20529 38314 20595 38317
rect 19425 38312 20595 38314
rect 19425 38256 19430 38312
rect 19486 38256 20534 38312
rect 20590 38256 20595 38312
rect 19425 38254 20595 38256
rect 19425 38251 19491 38254
rect 20529 38251 20595 38254
rect 19885 38178 19951 38181
rect 19750 38176 19951 38178
rect 19750 38120 19890 38176
rect 19946 38120 19951 38176
rect 19750 38118 19951 38120
rect 3658 38112 3974 38113
rect 3658 38048 3664 38112
rect 3728 38048 3744 38112
rect 3808 38048 3824 38112
rect 3888 38048 3904 38112
rect 3968 38048 3974 38112
rect 3658 38047 3974 38048
rect 11432 38112 11748 38113
rect 11432 38048 11438 38112
rect 11502 38048 11518 38112
rect 11582 38048 11598 38112
rect 11662 38048 11678 38112
rect 11742 38048 11748 38112
rect 11432 38047 11748 38048
rect 19206 38112 19522 38113
rect 19206 38048 19212 38112
rect 19276 38048 19292 38112
rect 19356 38048 19372 38112
rect 19436 38048 19452 38112
rect 19516 38048 19522 38112
rect 19206 38047 19522 38048
rect 19750 38045 19810 38118
rect 19885 38115 19951 38118
rect 26980 38112 27296 38113
rect 26980 38048 26986 38112
rect 27050 38048 27066 38112
rect 27130 38048 27146 38112
rect 27210 38048 27226 38112
rect 27290 38048 27296 38112
rect 26980 38047 27296 38048
rect 19750 38040 19859 38045
rect 19750 37984 19798 38040
rect 19854 37984 19859 38040
rect 19750 37982 19859 37984
rect 19793 37979 19859 37982
rect 20161 38040 20227 38045
rect 20161 37984 20166 38040
rect 20222 37984 20227 38040
rect 20161 37979 20227 37984
rect 19333 37906 19399 37909
rect 20164 37906 20224 37979
rect 19333 37904 20224 37906
rect 19333 37848 19338 37904
rect 19394 37848 20224 37904
rect 19333 37846 20224 37848
rect 19333 37843 19399 37846
rect 20069 37770 20135 37773
rect 20294 37770 20300 37772
rect 20069 37768 20300 37770
rect 20069 37712 20074 37768
rect 20130 37712 20300 37768
rect 20069 37710 20300 37712
rect 20069 37707 20135 37710
rect 20294 37708 20300 37710
rect 20364 37708 20370 37772
rect 4318 37568 4634 37569
rect 4318 37504 4324 37568
rect 4388 37504 4404 37568
rect 4468 37504 4484 37568
rect 4548 37504 4564 37568
rect 4628 37504 4634 37568
rect 4318 37503 4634 37504
rect 12092 37568 12408 37569
rect 12092 37504 12098 37568
rect 12162 37504 12178 37568
rect 12242 37504 12258 37568
rect 12322 37504 12338 37568
rect 12402 37504 12408 37568
rect 12092 37503 12408 37504
rect 19866 37568 20182 37569
rect 19866 37504 19872 37568
rect 19936 37504 19952 37568
rect 20016 37504 20032 37568
rect 20096 37504 20112 37568
rect 20176 37504 20182 37568
rect 19866 37503 20182 37504
rect 27640 37568 27956 37569
rect 27640 37504 27646 37568
rect 27710 37504 27726 37568
rect 27790 37504 27806 37568
rect 27870 37504 27886 37568
rect 27950 37504 27956 37568
rect 27640 37503 27956 37504
rect 19333 37362 19399 37365
rect 20161 37362 20227 37365
rect 21817 37362 21883 37365
rect 19333 37360 21883 37362
rect 19333 37304 19338 37360
rect 19394 37304 20166 37360
rect 20222 37304 21822 37360
rect 21878 37304 21883 37360
rect 19333 37302 21883 37304
rect 19333 37299 19399 37302
rect 20161 37299 20227 37302
rect 21817 37299 21883 37302
rect 19517 37226 19583 37229
rect 20662 37226 20668 37228
rect 19517 37224 20668 37226
rect 19517 37168 19522 37224
rect 19578 37168 20668 37224
rect 19517 37166 20668 37168
rect 19517 37163 19583 37166
rect 20662 37164 20668 37166
rect 20732 37226 20738 37228
rect 20805 37226 20871 37229
rect 20732 37224 20871 37226
rect 20732 37168 20810 37224
rect 20866 37168 20871 37224
rect 20732 37166 20871 37168
rect 20732 37164 20738 37166
rect 20805 37163 20871 37166
rect 3658 37024 3974 37025
rect 3658 36960 3664 37024
rect 3728 36960 3744 37024
rect 3808 36960 3824 37024
rect 3888 36960 3904 37024
rect 3968 36960 3974 37024
rect 3658 36959 3974 36960
rect 11432 37024 11748 37025
rect 11432 36960 11438 37024
rect 11502 36960 11518 37024
rect 11582 36960 11598 37024
rect 11662 36960 11678 37024
rect 11742 36960 11748 37024
rect 11432 36959 11748 36960
rect 19206 37024 19522 37025
rect 19206 36960 19212 37024
rect 19276 36960 19292 37024
rect 19356 36960 19372 37024
rect 19436 36960 19452 37024
rect 19516 36960 19522 37024
rect 19206 36959 19522 36960
rect 26980 37024 27296 37025
rect 26980 36960 26986 37024
rect 27050 36960 27066 37024
rect 27130 36960 27146 37024
rect 27210 36960 27226 37024
rect 27290 36960 27296 37024
rect 26980 36959 27296 36960
rect 19517 36818 19583 36821
rect 20294 36818 20300 36820
rect 19517 36816 20300 36818
rect 19517 36760 19522 36816
rect 19578 36760 20300 36816
rect 19517 36758 20300 36760
rect 19517 36755 19583 36758
rect 20294 36756 20300 36758
rect 20364 36756 20370 36820
rect 21909 36684 21975 36685
rect 21909 36682 21956 36684
rect 21864 36680 21956 36682
rect 21864 36624 21914 36680
rect 21864 36622 21956 36624
rect 21909 36620 21956 36622
rect 22020 36620 22026 36684
rect 21909 36619 21975 36620
rect 4318 36480 4634 36481
rect 4318 36416 4324 36480
rect 4388 36416 4404 36480
rect 4468 36416 4484 36480
rect 4548 36416 4564 36480
rect 4628 36416 4634 36480
rect 4318 36415 4634 36416
rect 12092 36480 12408 36481
rect 12092 36416 12098 36480
rect 12162 36416 12178 36480
rect 12242 36416 12258 36480
rect 12322 36416 12338 36480
rect 12402 36416 12408 36480
rect 12092 36415 12408 36416
rect 19866 36480 20182 36481
rect 19866 36416 19872 36480
rect 19936 36416 19952 36480
rect 20016 36416 20032 36480
rect 20096 36416 20112 36480
rect 20176 36416 20182 36480
rect 19866 36415 20182 36416
rect 27640 36480 27956 36481
rect 27640 36416 27646 36480
rect 27710 36416 27726 36480
rect 27790 36416 27806 36480
rect 27870 36416 27886 36480
rect 27950 36416 27956 36480
rect 27640 36415 27956 36416
rect 19057 36274 19123 36277
rect 22093 36274 22159 36277
rect 19057 36272 22159 36274
rect 19057 36216 19062 36272
rect 19118 36216 22098 36272
rect 22154 36216 22159 36272
rect 19057 36214 22159 36216
rect 19057 36211 19123 36214
rect 22093 36211 22159 36214
rect 10542 36076 10548 36140
rect 10612 36138 10618 36140
rect 22277 36138 22343 36141
rect 10612 36136 22343 36138
rect 10612 36080 22282 36136
rect 22338 36080 22343 36136
rect 10612 36078 22343 36080
rect 10612 36076 10618 36078
rect 22277 36075 22343 36078
rect 14273 36002 14339 36005
rect 18454 36002 18460 36004
rect 14273 36000 18460 36002
rect 14273 35944 14278 36000
rect 14334 35944 18460 36000
rect 14273 35942 18460 35944
rect 14273 35939 14339 35942
rect 18454 35940 18460 35942
rect 18524 35940 18530 36004
rect 3658 35936 3974 35937
rect 3658 35872 3664 35936
rect 3728 35872 3744 35936
rect 3808 35872 3824 35936
rect 3888 35872 3904 35936
rect 3968 35872 3974 35936
rect 3658 35871 3974 35872
rect 11432 35936 11748 35937
rect 11432 35872 11438 35936
rect 11502 35872 11518 35936
rect 11582 35872 11598 35936
rect 11662 35872 11678 35936
rect 11742 35872 11748 35936
rect 11432 35871 11748 35872
rect 19206 35936 19522 35937
rect 19206 35872 19212 35936
rect 19276 35872 19292 35936
rect 19356 35872 19372 35936
rect 19436 35872 19452 35936
rect 19516 35872 19522 35936
rect 19206 35871 19522 35872
rect 26980 35936 27296 35937
rect 26980 35872 26986 35936
rect 27050 35872 27066 35936
rect 27130 35872 27146 35936
rect 27210 35872 27226 35936
rect 27290 35872 27296 35936
rect 26980 35871 27296 35872
rect 4318 35392 4634 35393
rect 4318 35328 4324 35392
rect 4388 35328 4404 35392
rect 4468 35328 4484 35392
rect 4548 35328 4564 35392
rect 4628 35328 4634 35392
rect 4318 35327 4634 35328
rect 12092 35392 12408 35393
rect 12092 35328 12098 35392
rect 12162 35328 12178 35392
rect 12242 35328 12258 35392
rect 12322 35328 12338 35392
rect 12402 35328 12408 35392
rect 12092 35327 12408 35328
rect 19866 35392 20182 35393
rect 19866 35328 19872 35392
rect 19936 35328 19952 35392
rect 20016 35328 20032 35392
rect 20096 35328 20112 35392
rect 20176 35328 20182 35392
rect 19866 35327 20182 35328
rect 27640 35392 27956 35393
rect 27640 35328 27646 35392
rect 27710 35328 27726 35392
rect 27790 35328 27806 35392
rect 27870 35328 27886 35392
rect 27950 35328 27956 35392
rect 27640 35327 27956 35328
rect 12709 35050 12775 35053
rect 13721 35050 13787 35053
rect 12709 35048 13787 35050
rect 12709 34992 12714 35048
rect 12770 34992 13726 35048
rect 13782 34992 13787 35048
rect 12709 34990 13787 34992
rect 12709 34987 12775 34990
rect 13721 34987 13787 34990
rect 3658 34848 3974 34849
rect 3658 34784 3664 34848
rect 3728 34784 3744 34848
rect 3808 34784 3824 34848
rect 3888 34784 3904 34848
rect 3968 34784 3974 34848
rect 3658 34783 3974 34784
rect 11432 34848 11748 34849
rect 11432 34784 11438 34848
rect 11502 34784 11518 34848
rect 11582 34784 11598 34848
rect 11662 34784 11678 34848
rect 11742 34784 11748 34848
rect 11432 34783 11748 34784
rect 19206 34848 19522 34849
rect 19206 34784 19212 34848
rect 19276 34784 19292 34848
rect 19356 34784 19372 34848
rect 19436 34784 19452 34848
rect 19516 34784 19522 34848
rect 19206 34783 19522 34784
rect 26980 34848 27296 34849
rect 26980 34784 26986 34848
rect 27050 34784 27066 34848
rect 27130 34784 27146 34848
rect 27210 34784 27226 34848
rect 27290 34784 27296 34848
rect 26980 34783 27296 34784
rect 4318 34304 4634 34305
rect 4318 34240 4324 34304
rect 4388 34240 4404 34304
rect 4468 34240 4484 34304
rect 4548 34240 4564 34304
rect 4628 34240 4634 34304
rect 4318 34239 4634 34240
rect 12092 34304 12408 34305
rect 12092 34240 12098 34304
rect 12162 34240 12178 34304
rect 12242 34240 12258 34304
rect 12322 34240 12338 34304
rect 12402 34240 12408 34304
rect 12092 34239 12408 34240
rect 19866 34304 20182 34305
rect 19866 34240 19872 34304
rect 19936 34240 19952 34304
rect 20016 34240 20032 34304
rect 20096 34240 20112 34304
rect 20176 34240 20182 34304
rect 19866 34239 20182 34240
rect 27640 34304 27956 34305
rect 27640 34240 27646 34304
rect 27710 34240 27726 34304
rect 27790 34240 27806 34304
rect 27870 34240 27886 34304
rect 27950 34240 27956 34304
rect 27640 34239 27956 34240
rect 18505 34100 18571 34101
rect 18454 34036 18460 34100
rect 18524 34098 18571 34100
rect 18524 34096 18616 34098
rect 18566 34040 18616 34096
rect 18524 34038 18616 34040
rect 18524 34036 18571 34038
rect 18505 34035 18571 34036
rect 18597 33962 18663 33965
rect 19149 33962 19215 33965
rect 18597 33960 19215 33962
rect 18597 33904 18602 33960
rect 18658 33904 19154 33960
rect 19210 33904 19215 33960
rect 18597 33902 19215 33904
rect 18597 33899 18663 33902
rect 19149 33899 19215 33902
rect 3658 33760 3974 33761
rect 3658 33696 3664 33760
rect 3728 33696 3744 33760
rect 3808 33696 3824 33760
rect 3888 33696 3904 33760
rect 3968 33696 3974 33760
rect 3658 33695 3974 33696
rect 11432 33760 11748 33761
rect 11432 33696 11438 33760
rect 11502 33696 11518 33760
rect 11582 33696 11598 33760
rect 11662 33696 11678 33760
rect 11742 33696 11748 33760
rect 11432 33695 11748 33696
rect 19206 33760 19522 33761
rect 19206 33696 19212 33760
rect 19276 33696 19292 33760
rect 19356 33696 19372 33760
rect 19436 33696 19452 33760
rect 19516 33696 19522 33760
rect 19206 33695 19522 33696
rect 26980 33760 27296 33761
rect 26980 33696 26986 33760
rect 27050 33696 27066 33760
rect 27130 33696 27146 33760
rect 27210 33696 27226 33760
rect 27290 33696 27296 33760
rect 26980 33695 27296 33696
rect 11605 33418 11671 33421
rect 12525 33418 12591 33421
rect 11605 33416 12591 33418
rect 11605 33360 11610 33416
rect 11666 33360 12530 33416
rect 12586 33360 12591 33416
rect 11605 33358 12591 33360
rect 11605 33355 11671 33358
rect 12525 33355 12591 33358
rect 4318 33216 4634 33217
rect 4318 33152 4324 33216
rect 4388 33152 4404 33216
rect 4468 33152 4484 33216
rect 4548 33152 4564 33216
rect 4628 33152 4634 33216
rect 4318 33151 4634 33152
rect 12092 33216 12408 33217
rect 12092 33152 12098 33216
rect 12162 33152 12178 33216
rect 12242 33152 12258 33216
rect 12322 33152 12338 33216
rect 12402 33152 12408 33216
rect 12092 33151 12408 33152
rect 19866 33216 20182 33217
rect 19866 33152 19872 33216
rect 19936 33152 19952 33216
rect 20016 33152 20032 33216
rect 20096 33152 20112 33216
rect 20176 33152 20182 33216
rect 19866 33151 20182 33152
rect 27640 33216 27956 33217
rect 27640 33152 27646 33216
rect 27710 33152 27726 33216
rect 27790 33152 27806 33216
rect 27870 33152 27886 33216
rect 27950 33152 27956 33216
rect 27640 33151 27956 33152
rect 3658 32672 3974 32673
rect 3658 32608 3664 32672
rect 3728 32608 3744 32672
rect 3808 32608 3824 32672
rect 3888 32608 3904 32672
rect 3968 32608 3974 32672
rect 3658 32607 3974 32608
rect 11432 32672 11748 32673
rect 11432 32608 11438 32672
rect 11502 32608 11518 32672
rect 11582 32608 11598 32672
rect 11662 32608 11678 32672
rect 11742 32608 11748 32672
rect 11432 32607 11748 32608
rect 19206 32672 19522 32673
rect 19206 32608 19212 32672
rect 19276 32608 19292 32672
rect 19356 32608 19372 32672
rect 19436 32608 19452 32672
rect 19516 32608 19522 32672
rect 19206 32607 19522 32608
rect 26980 32672 27296 32673
rect 26980 32608 26986 32672
rect 27050 32608 27066 32672
rect 27130 32608 27146 32672
rect 27210 32608 27226 32672
rect 27290 32608 27296 32672
rect 26980 32607 27296 32608
rect 20069 32466 20135 32469
rect 20897 32466 20963 32469
rect 20069 32464 20963 32466
rect 20069 32408 20074 32464
rect 20130 32408 20902 32464
rect 20958 32408 20963 32464
rect 20069 32406 20963 32408
rect 20069 32403 20135 32406
rect 20897 32403 20963 32406
rect 20161 32330 20227 32333
rect 22553 32330 22619 32333
rect 20161 32328 22619 32330
rect 20161 32272 20166 32328
rect 20222 32272 22558 32328
rect 22614 32272 22619 32328
rect 20161 32270 22619 32272
rect 20161 32267 20227 32270
rect 22553 32267 22619 32270
rect 4318 32128 4634 32129
rect 4318 32064 4324 32128
rect 4388 32064 4404 32128
rect 4468 32064 4484 32128
rect 4548 32064 4564 32128
rect 4628 32064 4634 32128
rect 4318 32063 4634 32064
rect 12092 32128 12408 32129
rect 12092 32064 12098 32128
rect 12162 32064 12178 32128
rect 12242 32064 12258 32128
rect 12322 32064 12338 32128
rect 12402 32064 12408 32128
rect 12092 32063 12408 32064
rect 19866 32128 20182 32129
rect 19866 32064 19872 32128
rect 19936 32064 19952 32128
rect 20016 32064 20032 32128
rect 20096 32064 20112 32128
rect 20176 32064 20182 32128
rect 19866 32063 20182 32064
rect 27640 32128 27956 32129
rect 27640 32064 27646 32128
rect 27710 32064 27726 32128
rect 27790 32064 27806 32128
rect 27870 32064 27886 32128
rect 27950 32064 27956 32128
rect 27640 32063 27956 32064
rect 16665 31922 16731 31925
rect 20345 31924 20411 31925
rect 16982 31922 16988 31924
rect 16665 31920 16988 31922
rect 16665 31864 16670 31920
rect 16726 31864 16988 31920
rect 16665 31862 16988 31864
rect 16665 31859 16731 31862
rect 16982 31860 16988 31862
rect 17052 31860 17058 31924
rect 20294 31922 20300 31924
rect 20254 31862 20300 31922
rect 20364 31920 20411 31924
rect 20406 31864 20411 31920
rect 20294 31860 20300 31862
rect 20364 31860 20411 31864
rect 20345 31859 20411 31860
rect 20345 31652 20411 31653
rect 20294 31588 20300 31652
rect 20364 31650 20411 31652
rect 20364 31648 20456 31650
rect 20406 31592 20456 31648
rect 20364 31590 20456 31592
rect 20364 31588 20411 31590
rect 20345 31587 20411 31588
rect 3658 31584 3974 31585
rect 3658 31520 3664 31584
rect 3728 31520 3744 31584
rect 3808 31520 3824 31584
rect 3888 31520 3904 31584
rect 3968 31520 3974 31584
rect 3658 31519 3974 31520
rect 11432 31584 11748 31585
rect 11432 31520 11438 31584
rect 11502 31520 11518 31584
rect 11582 31520 11598 31584
rect 11662 31520 11678 31584
rect 11742 31520 11748 31584
rect 11432 31519 11748 31520
rect 19206 31584 19522 31585
rect 19206 31520 19212 31584
rect 19276 31520 19292 31584
rect 19356 31520 19372 31584
rect 19436 31520 19452 31584
rect 19516 31520 19522 31584
rect 19206 31519 19522 31520
rect 26980 31584 27296 31585
rect 26980 31520 26986 31584
rect 27050 31520 27066 31584
rect 27130 31520 27146 31584
rect 27210 31520 27226 31584
rect 27290 31520 27296 31584
rect 26980 31519 27296 31520
rect 4318 31040 4634 31041
rect 4318 30976 4324 31040
rect 4388 30976 4404 31040
rect 4468 30976 4484 31040
rect 4548 30976 4564 31040
rect 4628 30976 4634 31040
rect 4318 30975 4634 30976
rect 12092 31040 12408 31041
rect 12092 30976 12098 31040
rect 12162 30976 12178 31040
rect 12242 30976 12258 31040
rect 12322 30976 12338 31040
rect 12402 30976 12408 31040
rect 12092 30975 12408 30976
rect 19866 31040 20182 31041
rect 19866 30976 19872 31040
rect 19936 30976 19952 31040
rect 20016 30976 20032 31040
rect 20096 30976 20112 31040
rect 20176 30976 20182 31040
rect 19866 30975 20182 30976
rect 27640 31040 27956 31041
rect 27640 30976 27646 31040
rect 27710 30976 27726 31040
rect 27790 30976 27806 31040
rect 27870 30976 27886 31040
rect 27950 30976 27956 31040
rect 27640 30975 27956 30976
rect 26693 30700 26759 30701
rect 26693 30698 26740 30700
rect 26648 30696 26740 30698
rect 26648 30640 26698 30696
rect 26648 30638 26740 30640
rect 26693 30636 26740 30638
rect 26804 30636 26810 30700
rect 26693 30635 26759 30636
rect 3658 30496 3974 30497
rect 3658 30432 3664 30496
rect 3728 30432 3744 30496
rect 3808 30432 3824 30496
rect 3888 30432 3904 30496
rect 3968 30432 3974 30496
rect 3658 30431 3974 30432
rect 11432 30496 11748 30497
rect 11432 30432 11438 30496
rect 11502 30432 11518 30496
rect 11582 30432 11598 30496
rect 11662 30432 11678 30496
rect 11742 30432 11748 30496
rect 11432 30431 11748 30432
rect 19206 30496 19522 30497
rect 19206 30432 19212 30496
rect 19276 30432 19292 30496
rect 19356 30432 19372 30496
rect 19436 30432 19452 30496
rect 19516 30432 19522 30496
rect 19206 30431 19522 30432
rect 26980 30496 27296 30497
rect 26980 30432 26986 30496
rect 27050 30432 27066 30496
rect 27130 30432 27146 30496
rect 27210 30432 27226 30496
rect 27290 30432 27296 30496
rect 26980 30431 27296 30432
rect 23565 30292 23631 30293
rect 23565 30288 23612 30292
rect 23676 30290 23682 30292
rect 23565 30232 23570 30288
rect 23565 30228 23612 30232
rect 23676 30230 23722 30290
rect 23676 30228 23682 30230
rect 23565 30227 23631 30228
rect 4318 29952 4634 29953
rect 4318 29888 4324 29952
rect 4388 29888 4404 29952
rect 4468 29888 4484 29952
rect 4548 29888 4564 29952
rect 4628 29888 4634 29952
rect 4318 29887 4634 29888
rect 12092 29952 12408 29953
rect 12092 29888 12098 29952
rect 12162 29888 12178 29952
rect 12242 29888 12258 29952
rect 12322 29888 12338 29952
rect 12402 29888 12408 29952
rect 12092 29887 12408 29888
rect 19866 29952 20182 29953
rect 19866 29888 19872 29952
rect 19936 29888 19952 29952
rect 20016 29888 20032 29952
rect 20096 29888 20112 29952
rect 20176 29888 20182 29952
rect 19866 29887 20182 29888
rect 27640 29952 27956 29953
rect 27640 29888 27646 29952
rect 27710 29888 27726 29952
rect 27790 29888 27806 29952
rect 27870 29888 27886 29952
rect 27950 29888 27956 29952
rect 27640 29887 27956 29888
rect 3658 29408 3974 29409
rect 3658 29344 3664 29408
rect 3728 29344 3744 29408
rect 3808 29344 3824 29408
rect 3888 29344 3904 29408
rect 3968 29344 3974 29408
rect 3658 29343 3974 29344
rect 11432 29408 11748 29409
rect 11432 29344 11438 29408
rect 11502 29344 11518 29408
rect 11582 29344 11598 29408
rect 11662 29344 11678 29408
rect 11742 29344 11748 29408
rect 11432 29343 11748 29344
rect 19206 29408 19522 29409
rect 19206 29344 19212 29408
rect 19276 29344 19292 29408
rect 19356 29344 19372 29408
rect 19436 29344 19452 29408
rect 19516 29344 19522 29408
rect 19206 29343 19522 29344
rect 26980 29408 27296 29409
rect 26980 29344 26986 29408
rect 27050 29344 27066 29408
rect 27130 29344 27146 29408
rect 27210 29344 27226 29408
rect 27290 29344 27296 29408
rect 26980 29343 27296 29344
rect 19517 29202 19583 29205
rect 20662 29202 20668 29204
rect 19517 29200 20668 29202
rect 19517 29144 19522 29200
rect 19578 29144 20668 29200
rect 19517 29142 20668 29144
rect 19517 29139 19583 29142
rect 20662 29140 20668 29142
rect 20732 29140 20738 29204
rect 4318 28864 4634 28865
rect 4318 28800 4324 28864
rect 4388 28800 4404 28864
rect 4468 28800 4484 28864
rect 4548 28800 4564 28864
rect 4628 28800 4634 28864
rect 4318 28799 4634 28800
rect 12092 28864 12408 28865
rect 12092 28800 12098 28864
rect 12162 28800 12178 28864
rect 12242 28800 12258 28864
rect 12322 28800 12338 28864
rect 12402 28800 12408 28864
rect 12092 28799 12408 28800
rect 19866 28864 20182 28865
rect 19866 28800 19872 28864
rect 19936 28800 19952 28864
rect 20016 28800 20032 28864
rect 20096 28800 20112 28864
rect 20176 28800 20182 28864
rect 19866 28799 20182 28800
rect 27640 28864 27956 28865
rect 27640 28800 27646 28864
rect 27710 28800 27726 28864
rect 27790 28800 27806 28864
rect 27870 28800 27886 28864
rect 27950 28800 27956 28864
rect 27640 28799 27956 28800
rect 13670 28732 13676 28796
rect 13740 28794 13746 28796
rect 14273 28794 14339 28797
rect 13740 28792 14339 28794
rect 13740 28736 14278 28792
rect 14334 28736 14339 28792
rect 13740 28734 14339 28736
rect 13740 28732 13746 28734
rect 14273 28731 14339 28734
rect 21909 28660 21975 28661
rect 21909 28656 21956 28660
rect 22020 28658 22026 28660
rect 21909 28600 21914 28656
rect 21909 28596 21956 28600
rect 22020 28598 22066 28658
rect 22020 28596 22026 28598
rect 21909 28595 21975 28596
rect 20897 28522 20963 28525
rect 28758 28522 28764 28524
rect 20897 28520 28764 28522
rect 20897 28464 20902 28520
rect 20958 28464 28764 28520
rect 20897 28462 28764 28464
rect 20897 28459 20963 28462
rect 28758 28460 28764 28462
rect 28828 28460 28834 28524
rect 3658 28320 3974 28321
rect 3658 28256 3664 28320
rect 3728 28256 3744 28320
rect 3808 28256 3824 28320
rect 3888 28256 3904 28320
rect 3968 28256 3974 28320
rect 3658 28255 3974 28256
rect 11432 28320 11748 28321
rect 11432 28256 11438 28320
rect 11502 28256 11518 28320
rect 11582 28256 11598 28320
rect 11662 28256 11678 28320
rect 11742 28256 11748 28320
rect 11432 28255 11748 28256
rect 19206 28320 19522 28321
rect 19206 28256 19212 28320
rect 19276 28256 19292 28320
rect 19356 28256 19372 28320
rect 19436 28256 19452 28320
rect 19516 28256 19522 28320
rect 19206 28255 19522 28256
rect 26980 28320 27296 28321
rect 26980 28256 26986 28320
rect 27050 28256 27066 28320
rect 27130 28256 27146 28320
rect 27210 28256 27226 28320
rect 27290 28256 27296 28320
rect 26980 28255 27296 28256
rect 24485 28116 24551 28117
rect 24485 28112 24532 28116
rect 24596 28114 24602 28116
rect 24485 28056 24490 28112
rect 24485 28052 24532 28056
rect 24596 28054 24642 28114
rect 24596 28052 24602 28054
rect 24485 28051 24551 28052
rect 4318 27776 4634 27777
rect 4318 27712 4324 27776
rect 4388 27712 4404 27776
rect 4468 27712 4484 27776
rect 4548 27712 4564 27776
rect 4628 27712 4634 27776
rect 4318 27711 4634 27712
rect 12092 27776 12408 27777
rect 12092 27712 12098 27776
rect 12162 27712 12178 27776
rect 12242 27712 12258 27776
rect 12322 27712 12338 27776
rect 12402 27712 12408 27776
rect 12092 27711 12408 27712
rect 19866 27776 20182 27777
rect 19866 27712 19872 27776
rect 19936 27712 19952 27776
rect 20016 27712 20032 27776
rect 20096 27712 20112 27776
rect 20176 27712 20182 27776
rect 19866 27711 20182 27712
rect 27640 27776 27956 27777
rect 27640 27712 27646 27776
rect 27710 27712 27726 27776
rect 27790 27712 27806 27776
rect 27870 27712 27886 27776
rect 27950 27712 27956 27776
rect 27640 27711 27956 27712
rect 20529 27434 20595 27437
rect 23657 27434 23723 27437
rect 20529 27432 23723 27434
rect 20529 27376 20534 27432
rect 20590 27376 23662 27432
rect 23718 27376 23723 27432
rect 20529 27374 23723 27376
rect 20529 27371 20595 27374
rect 23657 27371 23723 27374
rect 3658 27232 3974 27233
rect 3658 27168 3664 27232
rect 3728 27168 3744 27232
rect 3808 27168 3824 27232
rect 3888 27168 3904 27232
rect 3968 27168 3974 27232
rect 3658 27167 3974 27168
rect 11432 27232 11748 27233
rect 11432 27168 11438 27232
rect 11502 27168 11518 27232
rect 11582 27168 11598 27232
rect 11662 27168 11678 27232
rect 11742 27168 11748 27232
rect 11432 27167 11748 27168
rect 19206 27232 19522 27233
rect 19206 27168 19212 27232
rect 19276 27168 19292 27232
rect 19356 27168 19372 27232
rect 19436 27168 19452 27232
rect 19516 27168 19522 27232
rect 19206 27167 19522 27168
rect 26980 27232 27296 27233
rect 26980 27168 26986 27232
rect 27050 27168 27066 27232
rect 27130 27168 27146 27232
rect 27210 27168 27226 27232
rect 27290 27168 27296 27232
rect 26980 27167 27296 27168
rect 4318 26688 4634 26689
rect 4318 26624 4324 26688
rect 4388 26624 4404 26688
rect 4468 26624 4484 26688
rect 4548 26624 4564 26688
rect 4628 26624 4634 26688
rect 4318 26623 4634 26624
rect 12092 26688 12408 26689
rect 12092 26624 12098 26688
rect 12162 26624 12178 26688
rect 12242 26624 12258 26688
rect 12322 26624 12338 26688
rect 12402 26624 12408 26688
rect 12092 26623 12408 26624
rect 19866 26688 20182 26689
rect 19866 26624 19872 26688
rect 19936 26624 19952 26688
rect 20016 26624 20032 26688
rect 20096 26624 20112 26688
rect 20176 26624 20182 26688
rect 19866 26623 20182 26624
rect 27640 26688 27956 26689
rect 27640 26624 27646 26688
rect 27710 26624 27726 26688
rect 27790 26624 27806 26688
rect 27870 26624 27886 26688
rect 27950 26624 27956 26688
rect 27640 26623 27956 26624
rect 3658 26144 3974 26145
rect 3658 26080 3664 26144
rect 3728 26080 3744 26144
rect 3808 26080 3824 26144
rect 3888 26080 3904 26144
rect 3968 26080 3974 26144
rect 3658 26079 3974 26080
rect 11432 26144 11748 26145
rect 11432 26080 11438 26144
rect 11502 26080 11518 26144
rect 11582 26080 11598 26144
rect 11662 26080 11678 26144
rect 11742 26080 11748 26144
rect 11432 26079 11748 26080
rect 19206 26144 19522 26145
rect 19206 26080 19212 26144
rect 19276 26080 19292 26144
rect 19356 26080 19372 26144
rect 19436 26080 19452 26144
rect 19516 26080 19522 26144
rect 19206 26079 19522 26080
rect 26980 26144 27296 26145
rect 26980 26080 26986 26144
rect 27050 26080 27066 26144
rect 27130 26080 27146 26144
rect 27210 26080 27226 26144
rect 27290 26080 27296 26144
rect 26980 26079 27296 26080
rect 27705 25802 27771 25805
rect 28533 25802 28599 25805
rect 27705 25800 28599 25802
rect 27705 25744 27710 25800
rect 27766 25744 28538 25800
rect 28594 25744 28599 25800
rect 27705 25742 28599 25744
rect 27705 25739 27771 25742
rect 28030 25669 28090 25742
rect 28533 25739 28599 25742
rect 28030 25664 28139 25669
rect 28030 25608 28078 25664
rect 28134 25608 28139 25664
rect 28030 25606 28139 25608
rect 28073 25603 28139 25606
rect 4318 25600 4634 25601
rect 4318 25536 4324 25600
rect 4388 25536 4404 25600
rect 4468 25536 4484 25600
rect 4548 25536 4564 25600
rect 4628 25536 4634 25600
rect 4318 25535 4634 25536
rect 12092 25600 12408 25601
rect 12092 25536 12098 25600
rect 12162 25536 12178 25600
rect 12242 25536 12258 25600
rect 12322 25536 12338 25600
rect 12402 25536 12408 25600
rect 12092 25535 12408 25536
rect 19866 25600 20182 25601
rect 19866 25536 19872 25600
rect 19936 25536 19952 25600
rect 20016 25536 20032 25600
rect 20096 25536 20112 25600
rect 20176 25536 20182 25600
rect 19866 25535 20182 25536
rect 27640 25600 27956 25601
rect 27640 25536 27646 25600
rect 27710 25536 27726 25600
rect 27790 25536 27806 25600
rect 27870 25536 27886 25600
rect 27950 25536 27956 25600
rect 27640 25535 27956 25536
rect 3658 25056 3974 25057
rect 3658 24992 3664 25056
rect 3728 24992 3744 25056
rect 3808 24992 3824 25056
rect 3888 24992 3904 25056
rect 3968 24992 3974 25056
rect 3658 24991 3974 24992
rect 11432 25056 11748 25057
rect 11432 24992 11438 25056
rect 11502 24992 11518 25056
rect 11582 24992 11598 25056
rect 11662 24992 11678 25056
rect 11742 24992 11748 25056
rect 11432 24991 11748 24992
rect 19206 25056 19522 25057
rect 19206 24992 19212 25056
rect 19276 24992 19292 25056
rect 19356 24992 19372 25056
rect 19436 24992 19452 25056
rect 19516 24992 19522 25056
rect 19206 24991 19522 24992
rect 26980 25056 27296 25057
rect 26980 24992 26986 25056
rect 27050 24992 27066 25056
rect 27130 24992 27146 25056
rect 27210 24992 27226 25056
rect 27290 24992 27296 25056
rect 26980 24991 27296 24992
rect 21633 24578 21699 24581
rect 24117 24578 24183 24581
rect 21633 24576 24183 24578
rect 21633 24520 21638 24576
rect 21694 24520 24122 24576
rect 24178 24520 24183 24576
rect 21633 24518 24183 24520
rect 21633 24515 21699 24518
rect 24117 24515 24183 24518
rect 4318 24512 4634 24513
rect 4318 24448 4324 24512
rect 4388 24448 4404 24512
rect 4468 24448 4484 24512
rect 4548 24448 4564 24512
rect 4628 24448 4634 24512
rect 4318 24447 4634 24448
rect 12092 24512 12408 24513
rect 12092 24448 12098 24512
rect 12162 24448 12178 24512
rect 12242 24448 12258 24512
rect 12322 24448 12338 24512
rect 12402 24448 12408 24512
rect 12092 24447 12408 24448
rect 19866 24512 20182 24513
rect 19866 24448 19872 24512
rect 19936 24448 19952 24512
rect 20016 24448 20032 24512
rect 20096 24448 20112 24512
rect 20176 24448 20182 24512
rect 19866 24447 20182 24448
rect 27640 24512 27956 24513
rect 27640 24448 27646 24512
rect 27710 24448 27726 24512
rect 27790 24448 27806 24512
rect 27870 24448 27886 24512
rect 27950 24448 27956 24512
rect 27640 24447 27956 24448
rect 20253 24442 20319 24445
rect 21909 24442 21975 24445
rect 22461 24442 22527 24445
rect 20253 24440 22527 24442
rect 20253 24384 20258 24440
rect 20314 24384 21914 24440
rect 21970 24384 22466 24440
rect 22522 24384 22527 24440
rect 20253 24382 22527 24384
rect 20253 24379 20319 24382
rect 21909 24379 21975 24382
rect 22461 24379 22527 24382
rect 3658 23968 3974 23969
rect 3658 23904 3664 23968
rect 3728 23904 3744 23968
rect 3808 23904 3824 23968
rect 3888 23904 3904 23968
rect 3968 23904 3974 23968
rect 3658 23903 3974 23904
rect 11432 23968 11748 23969
rect 11432 23904 11438 23968
rect 11502 23904 11518 23968
rect 11582 23904 11598 23968
rect 11662 23904 11678 23968
rect 11742 23904 11748 23968
rect 11432 23903 11748 23904
rect 19206 23968 19522 23969
rect 19206 23904 19212 23968
rect 19276 23904 19292 23968
rect 19356 23904 19372 23968
rect 19436 23904 19452 23968
rect 19516 23904 19522 23968
rect 19206 23903 19522 23904
rect 26980 23968 27296 23969
rect 26980 23904 26986 23968
rect 27050 23904 27066 23968
rect 27130 23904 27146 23968
rect 27210 23904 27226 23968
rect 27290 23904 27296 23968
rect 26980 23903 27296 23904
rect 20345 23898 20411 23901
rect 20478 23898 20484 23900
rect 20345 23896 20484 23898
rect 20345 23840 20350 23896
rect 20406 23840 20484 23896
rect 20345 23838 20484 23840
rect 20345 23835 20411 23838
rect 20478 23836 20484 23838
rect 20548 23836 20554 23900
rect 18781 23626 18847 23629
rect 19241 23626 19307 23629
rect 18781 23624 19307 23626
rect 18781 23568 18786 23624
rect 18842 23568 19246 23624
rect 19302 23568 19307 23624
rect 18781 23566 19307 23568
rect 18781 23563 18847 23566
rect 19241 23563 19307 23566
rect 4318 23424 4634 23425
rect 4318 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4634 23424
rect 4318 23359 4634 23360
rect 12092 23424 12408 23425
rect 12092 23360 12098 23424
rect 12162 23360 12178 23424
rect 12242 23360 12258 23424
rect 12322 23360 12338 23424
rect 12402 23360 12408 23424
rect 12092 23359 12408 23360
rect 19866 23424 20182 23425
rect 19866 23360 19872 23424
rect 19936 23360 19952 23424
rect 20016 23360 20032 23424
rect 20096 23360 20112 23424
rect 20176 23360 20182 23424
rect 19866 23359 20182 23360
rect 27640 23424 27956 23425
rect 27640 23360 27646 23424
rect 27710 23360 27726 23424
rect 27790 23360 27806 23424
rect 27870 23360 27886 23424
rect 27950 23360 27956 23424
rect 27640 23359 27956 23360
rect 3658 22880 3974 22881
rect 3658 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3974 22880
rect 3658 22815 3974 22816
rect 11432 22880 11748 22881
rect 11432 22816 11438 22880
rect 11502 22816 11518 22880
rect 11582 22816 11598 22880
rect 11662 22816 11678 22880
rect 11742 22816 11748 22880
rect 11432 22815 11748 22816
rect 19206 22880 19522 22881
rect 19206 22816 19212 22880
rect 19276 22816 19292 22880
rect 19356 22816 19372 22880
rect 19436 22816 19452 22880
rect 19516 22816 19522 22880
rect 19206 22815 19522 22816
rect 26980 22880 27296 22881
rect 26980 22816 26986 22880
rect 27050 22816 27066 22880
rect 27130 22816 27146 22880
rect 27210 22816 27226 22880
rect 27290 22816 27296 22880
rect 26980 22815 27296 22816
rect 27153 22674 27219 22677
rect 28625 22674 28691 22677
rect 27153 22672 28691 22674
rect 27153 22616 27158 22672
rect 27214 22616 28630 22672
rect 28686 22616 28691 22672
rect 27153 22614 28691 22616
rect 27153 22611 27219 22614
rect 28625 22611 28691 22614
rect 27613 22538 27679 22541
rect 26558 22536 27679 22538
rect 26558 22480 27618 22536
rect 27674 22480 27679 22536
rect 26558 22478 27679 22480
rect 4318 22336 4634 22337
rect 4318 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4634 22336
rect 4318 22271 4634 22272
rect 12092 22336 12408 22337
rect 12092 22272 12098 22336
rect 12162 22272 12178 22336
rect 12242 22272 12258 22336
rect 12322 22272 12338 22336
rect 12402 22272 12408 22336
rect 12092 22271 12408 22272
rect 19866 22336 20182 22337
rect 19866 22272 19872 22336
rect 19936 22272 19952 22336
rect 20016 22272 20032 22336
rect 20096 22272 20112 22336
rect 20176 22272 20182 22336
rect 19866 22271 20182 22272
rect 23197 22266 23263 22269
rect 23565 22266 23631 22269
rect 26417 22266 26483 22269
rect 23197 22264 23631 22266
rect 23197 22208 23202 22264
rect 23258 22208 23570 22264
rect 23626 22208 23631 22264
rect 23197 22206 23631 22208
rect 23197 22203 23263 22206
rect 23565 22203 23631 22206
rect 26190 22264 26483 22266
rect 26190 22208 26422 22264
rect 26478 22208 26483 22264
rect 26190 22206 26483 22208
rect 26190 22133 26250 22206
rect 26417 22203 26483 22206
rect 26190 22128 26299 22133
rect 26190 22072 26238 22128
rect 26294 22072 26299 22128
rect 26190 22070 26299 22072
rect 26233 22067 26299 22070
rect 26417 22130 26483 22133
rect 26558 22130 26618 22478
rect 27613 22475 27679 22478
rect 27640 22336 27956 22337
rect 27640 22272 27646 22336
rect 27710 22272 27726 22336
rect 27790 22272 27806 22336
rect 27870 22272 27886 22336
rect 27950 22272 27956 22336
rect 27640 22271 27956 22272
rect 26417 22128 26618 22130
rect 26417 22072 26422 22128
rect 26478 22072 26618 22128
rect 26417 22070 26618 22072
rect 26417 22067 26483 22070
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 11432 21792 11748 21793
rect 11432 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11748 21792
rect 11432 21727 11748 21728
rect 19206 21792 19522 21793
rect 19206 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19522 21792
rect 19206 21727 19522 21728
rect 26980 21792 27296 21793
rect 26980 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27296 21792
rect 26980 21727 27296 21728
rect 23197 21450 23263 21453
rect 23749 21450 23815 21453
rect 23197 21448 23815 21450
rect 23197 21392 23202 21448
rect 23258 21392 23754 21448
rect 23810 21392 23815 21448
rect 23197 21390 23815 21392
rect 23197 21387 23263 21390
rect 23749 21387 23815 21390
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 12092 21248 12408 21249
rect 12092 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12408 21248
rect 12092 21183 12408 21184
rect 19866 21248 20182 21249
rect 19866 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20182 21248
rect 19866 21183 20182 21184
rect 27640 21248 27956 21249
rect 27640 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27956 21248
rect 27640 21183 27956 21184
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 11432 20704 11748 20705
rect 11432 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11748 20704
rect 11432 20639 11748 20640
rect 19206 20704 19522 20705
rect 19206 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19522 20704
rect 19206 20639 19522 20640
rect 26980 20704 27296 20705
rect 26980 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27296 20704
rect 26980 20639 27296 20640
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 12092 20160 12408 20161
rect 12092 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12408 20160
rect 12092 20095 12408 20096
rect 19866 20160 20182 20161
rect 19866 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20182 20160
rect 19866 20095 20182 20096
rect 27640 20160 27956 20161
rect 27640 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27956 20160
rect 27640 20095 27956 20096
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 3658 19551 3974 19552
rect 11432 19616 11748 19617
rect 11432 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11748 19616
rect 11432 19551 11748 19552
rect 19206 19616 19522 19617
rect 19206 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19522 19616
rect 19206 19551 19522 19552
rect 26980 19616 27296 19617
rect 26980 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27296 19616
rect 26980 19551 27296 19552
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 12092 19072 12408 19073
rect 12092 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12408 19072
rect 12092 19007 12408 19008
rect 19866 19072 20182 19073
rect 19866 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20182 19072
rect 19866 19007 20182 19008
rect 27640 19072 27956 19073
rect 27640 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27956 19072
rect 27640 19007 27956 19008
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 11432 18528 11748 18529
rect 11432 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11748 18528
rect 11432 18463 11748 18464
rect 19206 18528 19522 18529
rect 19206 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19522 18528
rect 19206 18463 19522 18464
rect 26980 18528 27296 18529
rect 26980 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27296 18528
rect 26980 18463 27296 18464
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 12092 17984 12408 17985
rect 12092 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12408 17984
rect 12092 17919 12408 17920
rect 19866 17984 20182 17985
rect 19866 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20182 17984
rect 19866 17919 20182 17920
rect 27640 17984 27956 17985
rect 27640 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27956 17984
rect 27640 17919 27956 17920
rect 20805 17914 20871 17917
rect 25681 17914 25747 17917
rect 20805 17912 25747 17914
rect 20805 17856 20810 17912
rect 20866 17856 25686 17912
rect 25742 17856 25747 17912
rect 20805 17854 25747 17856
rect 20805 17851 20871 17854
rect 25681 17851 25747 17854
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 11432 17440 11748 17441
rect 11432 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11748 17440
rect 11432 17375 11748 17376
rect 19206 17440 19522 17441
rect 19206 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19522 17440
rect 19206 17375 19522 17376
rect 26980 17440 27296 17441
rect 26980 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27296 17440
rect 26980 17375 27296 17376
rect 22093 17370 22159 17373
rect 24301 17370 24367 17373
rect 22093 17368 24367 17370
rect 22093 17312 22098 17368
rect 22154 17312 24306 17368
rect 24362 17312 24367 17368
rect 22093 17310 24367 17312
rect 22093 17307 22159 17310
rect 24301 17307 24367 17310
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 12092 16896 12408 16897
rect 12092 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12408 16896
rect 12092 16831 12408 16832
rect 19866 16896 20182 16897
rect 19866 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20182 16896
rect 19866 16831 20182 16832
rect 27640 16896 27956 16897
rect 27640 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27956 16896
rect 27640 16831 27956 16832
rect 17217 16690 17283 16693
rect 19609 16690 19675 16693
rect 17217 16688 19675 16690
rect 17217 16632 17222 16688
rect 17278 16632 19614 16688
rect 19670 16632 19675 16688
rect 17217 16630 19675 16632
rect 17217 16627 17283 16630
rect 19609 16627 19675 16630
rect 26734 16628 26740 16692
rect 26804 16690 26810 16692
rect 26877 16690 26943 16693
rect 26804 16688 26943 16690
rect 26804 16632 26882 16688
rect 26938 16632 26943 16688
rect 26804 16630 26943 16632
rect 26804 16628 26810 16630
rect 26877 16627 26943 16630
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 11432 16352 11748 16353
rect 11432 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11748 16352
rect 11432 16287 11748 16288
rect 19206 16352 19522 16353
rect 19206 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19522 16352
rect 19206 16287 19522 16288
rect 26980 16352 27296 16353
rect 26980 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27296 16352
rect 26980 16287 27296 16288
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 12092 15808 12408 15809
rect 12092 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12408 15808
rect 12092 15743 12408 15744
rect 19866 15808 20182 15809
rect 19866 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20182 15808
rect 19866 15743 20182 15744
rect 27640 15808 27956 15809
rect 27640 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27956 15808
rect 27640 15743 27956 15744
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 11432 15264 11748 15265
rect 11432 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11748 15264
rect 11432 15199 11748 15200
rect 19206 15264 19522 15265
rect 19206 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19522 15264
rect 19206 15199 19522 15200
rect 26980 15264 27296 15265
rect 26980 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27296 15264
rect 26980 15199 27296 15200
rect 16941 15196 17007 15197
rect 16941 15194 16988 15196
rect 16896 15192 16988 15194
rect 16896 15136 16946 15192
rect 16896 15134 16988 15136
rect 16941 15132 16988 15134
rect 17052 15132 17058 15196
rect 16941 15131 17007 15132
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 12092 14720 12408 14721
rect 12092 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12408 14720
rect 12092 14655 12408 14656
rect 19866 14720 20182 14721
rect 19866 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20182 14720
rect 19866 14655 20182 14656
rect 27640 14720 27956 14721
rect 27640 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27956 14720
rect 27640 14655 27956 14656
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 11432 14176 11748 14177
rect 11432 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11748 14176
rect 11432 14111 11748 14112
rect 19206 14176 19522 14177
rect 19206 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19522 14176
rect 19206 14111 19522 14112
rect 26980 14176 27296 14177
rect 26980 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27296 14176
rect 26980 14111 27296 14112
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 12092 13632 12408 13633
rect 12092 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12408 13632
rect 12092 13567 12408 13568
rect 19866 13632 20182 13633
rect 19866 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20182 13632
rect 19866 13567 20182 13568
rect 27640 13632 27956 13633
rect 27640 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27956 13632
rect 27640 13567 27956 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 11432 13088 11748 13089
rect 11432 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11748 13088
rect 11432 13023 11748 13024
rect 19206 13088 19522 13089
rect 19206 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19522 13088
rect 19206 13023 19522 13024
rect 26980 13088 27296 13089
rect 26980 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27296 13088
rect 26980 13023 27296 13024
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 12092 12544 12408 12545
rect 12092 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12408 12544
rect 12092 12479 12408 12480
rect 19866 12544 20182 12545
rect 19866 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20182 12544
rect 19866 12479 20182 12480
rect 27640 12544 27956 12545
rect 27640 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27956 12544
rect 27640 12479 27956 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 11432 12000 11748 12001
rect 11432 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11748 12000
rect 11432 11935 11748 11936
rect 19206 12000 19522 12001
rect 19206 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19522 12000
rect 19206 11935 19522 11936
rect 26980 12000 27296 12001
rect 26980 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27296 12000
rect 26980 11935 27296 11936
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 12092 11456 12408 11457
rect 12092 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12408 11456
rect 12092 11391 12408 11392
rect 19866 11456 20182 11457
rect 19866 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20182 11456
rect 19866 11391 20182 11392
rect 27640 11456 27956 11457
rect 27640 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27956 11456
rect 27640 11391 27956 11392
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 11432 10912 11748 10913
rect 11432 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11748 10912
rect 11432 10847 11748 10848
rect 19206 10912 19522 10913
rect 19206 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19522 10912
rect 19206 10847 19522 10848
rect 26980 10912 27296 10913
rect 26980 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27296 10912
rect 26980 10847 27296 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 12092 10368 12408 10369
rect 12092 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12408 10368
rect 12092 10303 12408 10304
rect 19866 10368 20182 10369
rect 19866 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20182 10368
rect 19866 10303 20182 10304
rect 27640 10368 27956 10369
rect 27640 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27956 10368
rect 27640 10303 27956 10304
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 11432 9824 11748 9825
rect 11432 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11748 9824
rect 11432 9759 11748 9760
rect 19206 9824 19522 9825
rect 19206 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19522 9824
rect 19206 9759 19522 9760
rect 26980 9824 27296 9825
rect 26980 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27296 9824
rect 26980 9759 27296 9760
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 12092 9280 12408 9281
rect 12092 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12408 9280
rect 12092 9215 12408 9216
rect 19866 9280 20182 9281
rect 19866 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20182 9280
rect 19866 9215 20182 9216
rect 27640 9280 27956 9281
rect 27640 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27956 9280
rect 27640 9215 27956 9216
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 11432 8736 11748 8737
rect 11432 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11748 8736
rect 11432 8671 11748 8672
rect 19206 8736 19522 8737
rect 19206 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19522 8736
rect 19206 8671 19522 8672
rect 26980 8736 27296 8737
rect 26980 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27296 8736
rect 26980 8671 27296 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 12092 8192 12408 8193
rect 12092 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12408 8192
rect 12092 8127 12408 8128
rect 19866 8192 20182 8193
rect 19866 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20182 8192
rect 19866 8127 20182 8128
rect 27640 8192 27956 8193
rect 27640 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27956 8192
rect 27640 8127 27956 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 11432 7648 11748 7649
rect 11432 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11748 7648
rect 11432 7583 11748 7584
rect 19206 7648 19522 7649
rect 19206 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19522 7648
rect 19206 7583 19522 7584
rect 26980 7648 27296 7649
rect 26980 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27296 7648
rect 26980 7583 27296 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 12092 7104 12408 7105
rect 12092 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12408 7104
rect 12092 7039 12408 7040
rect 19866 7104 20182 7105
rect 19866 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20182 7104
rect 19866 7039 20182 7040
rect 27640 7104 27956 7105
rect 27640 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27956 7104
rect 27640 7039 27956 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 11432 6560 11748 6561
rect 11432 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11748 6560
rect 11432 6495 11748 6496
rect 19206 6560 19522 6561
rect 19206 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19522 6560
rect 19206 6495 19522 6496
rect 26980 6560 27296 6561
rect 26980 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27296 6560
rect 26980 6495 27296 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 12092 6016 12408 6017
rect 12092 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12408 6016
rect 12092 5951 12408 5952
rect 19866 6016 20182 6017
rect 19866 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20182 6016
rect 19866 5951 20182 5952
rect 27640 6016 27956 6017
rect 27640 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27956 6016
rect 27640 5951 27956 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 11432 5472 11748 5473
rect 11432 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11748 5472
rect 11432 5407 11748 5408
rect 19206 5472 19522 5473
rect 19206 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19522 5472
rect 19206 5407 19522 5408
rect 26980 5472 27296 5473
rect 26980 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27296 5472
rect 26980 5407 27296 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 12092 4928 12408 4929
rect 12092 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12408 4928
rect 12092 4863 12408 4864
rect 19866 4928 20182 4929
rect 19866 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20182 4928
rect 19866 4863 20182 4864
rect 27640 4928 27956 4929
rect 27640 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27956 4928
rect 27640 4863 27956 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 11432 4384 11748 4385
rect 11432 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11748 4384
rect 11432 4319 11748 4320
rect 19206 4384 19522 4385
rect 19206 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19522 4384
rect 19206 4319 19522 4320
rect 26980 4384 27296 4385
rect 26980 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27296 4384
rect 26980 4319 27296 4320
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 12092 3840 12408 3841
rect 12092 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12408 3840
rect 12092 3775 12408 3776
rect 19866 3840 20182 3841
rect 19866 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20182 3840
rect 19866 3775 20182 3776
rect 27640 3840 27956 3841
rect 27640 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27956 3840
rect 27640 3775 27956 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 11432 3296 11748 3297
rect 11432 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11748 3296
rect 11432 3231 11748 3232
rect 19206 3296 19522 3297
rect 19206 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19522 3296
rect 19206 3231 19522 3232
rect 26980 3296 27296 3297
rect 26980 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27296 3296
rect 26980 3231 27296 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 12092 2752 12408 2753
rect 12092 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12408 2752
rect 12092 2687 12408 2688
rect 19866 2752 20182 2753
rect 19866 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20182 2752
rect 19866 2687 20182 2688
rect 27640 2752 27956 2753
rect 27640 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27956 2752
rect 27640 2687 27956 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 11432 2208 11748 2209
rect 11432 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11748 2208
rect 11432 2143 11748 2144
rect 19206 2208 19522 2209
rect 19206 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19522 2208
rect 19206 2143 19522 2144
rect 26980 2208 27296 2209
rect 26980 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27296 2208
rect 26980 2143 27296 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 12092 1664 12408 1665
rect 12092 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12408 1664
rect 12092 1599 12408 1600
rect 19866 1664 20182 1665
rect 19866 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20182 1664
rect 19866 1599 20182 1600
rect 27640 1664 27956 1665
rect 27640 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27956 1664
rect 27640 1599 27956 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 11432 1120 11748 1121
rect 11432 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11748 1120
rect 11432 1055 11748 1056
rect 19206 1120 19522 1121
rect 19206 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19522 1120
rect 19206 1055 19522 1056
rect 26980 1120 27296 1121
rect 26980 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27296 1120
rect 26980 1055 27296 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 12092 576 12408 577
rect 12092 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12408 576
rect 12092 511 12408 512
rect 19866 576 20182 577
rect 19866 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20182 576
rect 19866 511 20182 512
rect 27640 576 27956 577
rect 27640 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27956 576
rect 27640 511 27956 512
<< via3 >>
rect 11652 44780 11716 44844
rect 12204 44780 12268 44844
rect 21588 44840 21652 44844
rect 21588 44784 21638 44840
rect 21638 44784 21652 44840
rect 21588 44780 21652 44784
rect 27108 44780 27172 44844
rect 27660 44780 27724 44844
rect 23796 44644 23860 44708
rect 24348 44704 24412 44708
rect 24348 44648 24398 44704
rect 24398 44648 24412 44704
rect 24348 44644 24412 44648
rect 24900 44704 24964 44708
rect 24900 44648 24950 44704
rect 24950 44648 24964 44704
rect 24900 44644 24964 44648
rect 25452 44704 25516 44708
rect 25452 44648 25502 44704
rect 25502 44648 25516 44704
rect 25452 44644 25516 44648
rect 26004 44704 26068 44708
rect 26004 44648 26054 44704
rect 26054 44648 26068 44704
rect 26004 44644 26068 44648
rect 26556 44704 26620 44708
rect 26556 44648 26570 44704
rect 26570 44648 26620 44704
rect 26556 44644 26620 44648
rect 28212 44644 28276 44708
rect 3664 44636 3728 44640
rect 3664 44580 3668 44636
rect 3668 44580 3724 44636
rect 3724 44580 3728 44636
rect 3664 44576 3728 44580
rect 3744 44636 3808 44640
rect 3744 44580 3748 44636
rect 3748 44580 3804 44636
rect 3804 44580 3808 44636
rect 3744 44576 3808 44580
rect 3824 44636 3888 44640
rect 3824 44580 3828 44636
rect 3828 44580 3884 44636
rect 3884 44580 3888 44636
rect 3824 44576 3888 44580
rect 3904 44636 3968 44640
rect 3904 44580 3908 44636
rect 3908 44580 3964 44636
rect 3964 44580 3968 44636
rect 3904 44576 3968 44580
rect 11438 44636 11502 44640
rect 11438 44580 11442 44636
rect 11442 44580 11498 44636
rect 11498 44580 11502 44636
rect 11438 44576 11502 44580
rect 11518 44636 11582 44640
rect 11518 44580 11522 44636
rect 11522 44580 11578 44636
rect 11578 44580 11582 44636
rect 11518 44576 11582 44580
rect 11598 44636 11662 44640
rect 11598 44580 11602 44636
rect 11602 44580 11658 44636
rect 11658 44580 11662 44636
rect 11598 44576 11662 44580
rect 11678 44636 11742 44640
rect 11678 44580 11682 44636
rect 11682 44580 11738 44636
rect 11738 44580 11742 44636
rect 11678 44576 11742 44580
rect 19212 44636 19276 44640
rect 19212 44580 19216 44636
rect 19216 44580 19272 44636
rect 19272 44580 19276 44636
rect 19212 44576 19276 44580
rect 19292 44636 19356 44640
rect 19292 44580 19296 44636
rect 19296 44580 19352 44636
rect 19352 44580 19356 44636
rect 19292 44576 19356 44580
rect 19372 44636 19436 44640
rect 19372 44580 19376 44636
rect 19376 44580 19432 44636
rect 19432 44580 19436 44636
rect 19372 44576 19436 44580
rect 19452 44636 19516 44640
rect 19452 44580 19456 44636
rect 19456 44580 19512 44636
rect 19512 44580 19516 44636
rect 19452 44576 19516 44580
rect 26986 44636 27050 44640
rect 26986 44580 26990 44636
rect 26990 44580 27046 44636
rect 27046 44580 27050 44636
rect 26986 44576 27050 44580
rect 27066 44636 27130 44640
rect 27066 44580 27070 44636
rect 27070 44580 27126 44636
rect 27126 44580 27130 44636
rect 27066 44576 27130 44580
rect 27146 44636 27210 44640
rect 27146 44580 27150 44636
rect 27150 44580 27206 44636
rect 27206 44580 27210 44636
rect 27146 44576 27210 44580
rect 27226 44636 27290 44640
rect 27226 44580 27230 44636
rect 27230 44580 27286 44636
rect 27286 44580 27290 44636
rect 27226 44576 27290 44580
rect 7236 44568 7300 44572
rect 7236 44512 7250 44568
rect 7250 44512 7300 44568
rect 7236 44508 7300 44512
rect 7788 44508 7852 44572
rect 8340 44568 8404 44572
rect 8340 44512 8354 44568
rect 8354 44512 8404 44568
rect 8340 44508 8404 44512
rect 8892 44508 8956 44572
rect 9444 44508 9508 44572
rect 12756 44568 12820 44572
rect 12756 44512 12806 44568
rect 12806 44512 12820 44568
rect 12756 44508 12820 44512
rect 4324 44092 4388 44096
rect 4324 44036 4328 44092
rect 4328 44036 4384 44092
rect 4384 44036 4388 44092
rect 4324 44032 4388 44036
rect 4404 44092 4468 44096
rect 4404 44036 4408 44092
rect 4408 44036 4464 44092
rect 4464 44036 4468 44092
rect 4404 44032 4468 44036
rect 4484 44092 4548 44096
rect 4484 44036 4488 44092
rect 4488 44036 4544 44092
rect 4544 44036 4548 44092
rect 4484 44032 4548 44036
rect 4564 44092 4628 44096
rect 4564 44036 4568 44092
rect 4568 44036 4624 44092
rect 4624 44036 4628 44092
rect 4564 44032 4628 44036
rect 12098 44092 12162 44096
rect 12098 44036 12102 44092
rect 12102 44036 12158 44092
rect 12158 44036 12162 44092
rect 12098 44032 12162 44036
rect 12178 44092 12242 44096
rect 12178 44036 12182 44092
rect 12182 44036 12238 44092
rect 12238 44036 12242 44092
rect 12178 44032 12242 44036
rect 12258 44092 12322 44096
rect 12258 44036 12262 44092
rect 12262 44036 12318 44092
rect 12318 44036 12322 44092
rect 12258 44032 12322 44036
rect 12338 44092 12402 44096
rect 12338 44036 12342 44092
rect 12342 44036 12398 44092
rect 12398 44036 12402 44092
rect 12338 44032 12402 44036
rect 19872 44092 19936 44096
rect 19872 44036 19876 44092
rect 19876 44036 19932 44092
rect 19932 44036 19936 44092
rect 19872 44032 19936 44036
rect 19952 44092 20016 44096
rect 19952 44036 19956 44092
rect 19956 44036 20012 44092
rect 20012 44036 20016 44092
rect 19952 44032 20016 44036
rect 20032 44092 20096 44096
rect 20032 44036 20036 44092
rect 20036 44036 20092 44092
rect 20092 44036 20096 44092
rect 20032 44032 20096 44036
rect 20112 44092 20176 44096
rect 20112 44036 20116 44092
rect 20116 44036 20172 44092
rect 20172 44036 20176 44092
rect 20112 44032 20176 44036
rect 27646 44092 27710 44096
rect 27646 44036 27650 44092
rect 27650 44036 27706 44092
rect 27706 44036 27710 44092
rect 27646 44032 27710 44036
rect 27726 44092 27790 44096
rect 27726 44036 27730 44092
rect 27730 44036 27786 44092
rect 27786 44036 27790 44092
rect 27726 44032 27790 44036
rect 27806 44092 27870 44096
rect 27806 44036 27810 44092
rect 27810 44036 27866 44092
rect 27866 44036 27870 44092
rect 27806 44032 27870 44036
rect 27886 44092 27950 44096
rect 27886 44036 27890 44092
rect 27890 44036 27946 44092
rect 27946 44036 27950 44092
rect 27886 44032 27950 44036
rect 6132 43964 6196 44028
rect 6684 43964 6748 44028
rect 9996 43964 10060 44028
rect 13308 44024 13372 44028
rect 13308 43968 13322 44024
rect 13322 43968 13372 44024
rect 13308 43964 13372 43968
rect 16620 44024 16684 44028
rect 16620 43968 16634 44024
rect 16634 43968 16684 44024
rect 16620 43964 16684 43968
rect 17172 43964 17236 44028
rect 11100 43828 11164 43892
rect 13860 43752 13924 43756
rect 13860 43696 13874 43752
rect 13874 43696 13924 43752
rect 13860 43692 13924 43696
rect 3664 43548 3728 43552
rect 3664 43492 3668 43548
rect 3668 43492 3724 43548
rect 3724 43492 3728 43548
rect 3664 43488 3728 43492
rect 3744 43548 3808 43552
rect 3744 43492 3748 43548
rect 3748 43492 3804 43548
rect 3804 43492 3808 43548
rect 3744 43488 3808 43492
rect 3824 43548 3888 43552
rect 3824 43492 3828 43548
rect 3828 43492 3884 43548
rect 3884 43492 3888 43548
rect 3824 43488 3888 43492
rect 3904 43548 3968 43552
rect 3904 43492 3908 43548
rect 3908 43492 3964 43548
rect 3964 43492 3968 43548
rect 3904 43488 3968 43492
rect 11438 43548 11502 43552
rect 11438 43492 11442 43548
rect 11442 43492 11498 43548
rect 11498 43492 11502 43548
rect 11438 43488 11502 43492
rect 11518 43548 11582 43552
rect 11518 43492 11522 43548
rect 11522 43492 11578 43548
rect 11578 43492 11582 43548
rect 11518 43488 11582 43492
rect 11598 43548 11662 43552
rect 11598 43492 11602 43548
rect 11602 43492 11658 43548
rect 11658 43492 11662 43548
rect 11598 43488 11662 43492
rect 11678 43548 11742 43552
rect 11678 43492 11682 43548
rect 11682 43492 11738 43548
rect 11738 43492 11742 43548
rect 11678 43488 11742 43492
rect 19212 43548 19276 43552
rect 19212 43492 19216 43548
rect 19216 43492 19272 43548
rect 19272 43492 19276 43548
rect 19212 43488 19276 43492
rect 19292 43548 19356 43552
rect 19292 43492 19296 43548
rect 19296 43492 19352 43548
rect 19352 43492 19356 43548
rect 19292 43488 19356 43492
rect 19372 43548 19436 43552
rect 19372 43492 19376 43548
rect 19376 43492 19432 43548
rect 19432 43492 19436 43548
rect 19372 43488 19436 43492
rect 19452 43548 19516 43552
rect 19452 43492 19456 43548
rect 19456 43492 19512 43548
rect 19512 43492 19516 43548
rect 19452 43488 19516 43492
rect 26986 43548 27050 43552
rect 26986 43492 26990 43548
rect 26990 43492 27046 43548
rect 27046 43492 27050 43548
rect 26986 43488 27050 43492
rect 27066 43548 27130 43552
rect 27066 43492 27070 43548
rect 27070 43492 27126 43548
rect 27126 43492 27130 43548
rect 27066 43488 27130 43492
rect 27146 43548 27210 43552
rect 27146 43492 27150 43548
rect 27150 43492 27206 43548
rect 27206 43492 27210 43548
rect 27146 43488 27210 43492
rect 27226 43548 27290 43552
rect 27226 43492 27230 43548
rect 27230 43492 27286 43548
rect 27286 43492 27290 43548
rect 27226 43488 27290 43492
rect 14412 43480 14476 43484
rect 14412 43424 14426 43480
rect 14426 43424 14476 43480
rect 14412 43420 14476 43424
rect 18828 43284 18892 43348
rect 14964 43148 15028 43212
rect 18276 43148 18340 43212
rect 4324 43004 4388 43008
rect 4324 42948 4328 43004
rect 4328 42948 4384 43004
rect 4384 42948 4388 43004
rect 4324 42944 4388 42948
rect 4404 43004 4468 43008
rect 4404 42948 4408 43004
rect 4408 42948 4464 43004
rect 4464 42948 4468 43004
rect 4404 42944 4468 42948
rect 4484 43004 4548 43008
rect 4484 42948 4488 43004
rect 4488 42948 4544 43004
rect 4544 42948 4548 43004
rect 4484 42944 4548 42948
rect 4564 43004 4628 43008
rect 4564 42948 4568 43004
rect 4568 42948 4624 43004
rect 4624 42948 4628 43004
rect 4564 42944 4628 42948
rect 12098 43004 12162 43008
rect 12098 42948 12102 43004
rect 12102 42948 12158 43004
rect 12158 42948 12162 43004
rect 12098 42944 12162 42948
rect 12178 43004 12242 43008
rect 12178 42948 12182 43004
rect 12182 42948 12238 43004
rect 12238 42948 12242 43004
rect 12178 42944 12242 42948
rect 12258 43004 12322 43008
rect 12258 42948 12262 43004
rect 12262 42948 12318 43004
rect 12318 42948 12322 43004
rect 12258 42944 12322 42948
rect 12338 43004 12402 43008
rect 12338 42948 12342 43004
rect 12342 42948 12398 43004
rect 12398 42948 12402 43004
rect 12338 42944 12402 42948
rect 19872 43004 19936 43008
rect 19872 42948 19876 43004
rect 19876 42948 19932 43004
rect 19932 42948 19936 43004
rect 19872 42944 19936 42948
rect 19952 43004 20016 43008
rect 19952 42948 19956 43004
rect 19956 42948 20012 43004
rect 20012 42948 20016 43004
rect 19952 42944 20016 42948
rect 20032 43004 20096 43008
rect 20032 42948 20036 43004
rect 20036 42948 20092 43004
rect 20092 42948 20096 43004
rect 20032 42944 20096 42948
rect 20112 43004 20176 43008
rect 20112 42948 20116 43004
rect 20116 42948 20172 43004
rect 20172 42948 20176 43004
rect 20112 42944 20176 42948
rect 27646 43004 27710 43008
rect 27646 42948 27650 43004
rect 27650 42948 27706 43004
rect 27706 42948 27710 43004
rect 27646 42944 27710 42948
rect 27726 43004 27790 43008
rect 27726 42948 27730 43004
rect 27730 42948 27786 43004
rect 27786 42948 27790 43004
rect 27726 42944 27790 42948
rect 27806 43004 27870 43008
rect 27806 42948 27810 43004
rect 27810 42948 27866 43004
rect 27866 42948 27870 43004
rect 27806 42944 27870 42948
rect 27886 43004 27950 43008
rect 27886 42948 27890 43004
rect 27890 42948 27946 43004
rect 27946 42948 27950 43004
rect 27886 42944 27950 42948
rect 15516 42936 15580 42940
rect 15516 42880 15530 42936
rect 15530 42880 15580 42936
rect 15516 42876 15580 42880
rect 17724 42876 17788 42940
rect 3664 42460 3728 42464
rect 3664 42404 3668 42460
rect 3668 42404 3724 42460
rect 3724 42404 3728 42460
rect 3664 42400 3728 42404
rect 3744 42460 3808 42464
rect 3744 42404 3748 42460
rect 3748 42404 3804 42460
rect 3804 42404 3808 42460
rect 3744 42400 3808 42404
rect 3824 42460 3888 42464
rect 3824 42404 3828 42460
rect 3828 42404 3884 42460
rect 3884 42404 3888 42460
rect 3824 42400 3888 42404
rect 3904 42460 3968 42464
rect 3904 42404 3908 42460
rect 3908 42404 3964 42460
rect 3964 42404 3968 42460
rect 3904 42400 3968 42404
rect 11438 42460 11502 42464
rect 11438 42404 11442 42460
rect 11442 42404 11498 42460
rect 11498 42404 11502 42460
rect 11438 42400 11502 42404
rect 11518 42460 11582 42464
rect 11518 42404 11522 42460
rect 11522 42404 11578 42460
rect 11578 42404 11582 42460
rect 11518 42400 11582 42404
rect 11598 42460 11662 42464
rect 11598 42404 11602 42460
rect 11602 42404 11658 42460
rect 11658 42404 11662 42460
rect 11598 42400 11662 42404
rect 11678 42460 11742 42464
rect 11678 42404 11682 42460
rect 11682 42404 11738 42460
rect 11738 42404 11742 42460
rect 11678 42400 11742 42404
rect 19212 42460 19276 42464
rect 19212 42404 19216 42460
rect 19216 42404 19272 42460
rect 19272 42404 19276 42460
rect 19212 42400 19276 42404
rect 19292 42460 19356 42464
rect 19292 42404 19296 42460
rect 19296 42404 19352 42460
rect 19352 42404 19356 42460
rect 19292 42400 19356 42404
rect 19372 42460 19436 42464
rect 19372 42404 19376 42460
rect 19376 42404 19432 42460
rect 19432 42404 19436 42460
rect 19372 42400 19436 42404
rect 19452 42460 19516 42464
rect 19452 42404 19456 42460
rect 19456 42404 19512 42460
rect 19512 42404 19516 42460
rect 19452 42400 19516 42404
rect 26986 42460 27050 42464
rect 26986 42404 26990 42460
rect 26990 42404 27046 42460
rect 27046 42404 27050 42460
rect 26986 42400 27050 42404
rect 27066 42460 27130 42464
rect 27066 42404 27070 42460
rect 27070 42404 27126 42460
rect 27126 42404 27130 42460
rect 27066 42400 27130 42404
rect 27146 42460 27210 42464
rect 27146 42404 27150 42460
rect 27150 42404 27206 42460
rect 27206 42404 27210 42460
rect 27146 42400 27210 42404
rect 27226 42460 27290 42464
rect 27226 42404 27230 42460
rect 27230 42404 27286 42460
rect 27286 42404 27290 42460
rect 27226 42400 27290 42404
rect 23612 42256 23676 42260
rect 23612 42200 23662 42256
rect 23662 42200 23676 42256
rect 23612 42196 23676 42200
rect 4324 41916 4388 41920
rect 4324 41860 4328 41916
rect 4328 41860 4384 41916
rect 4384 41860 4388 41916
rect 4324 41856 4388 41860
rect 4404 41916 4468 41920
rect 4404 41860 4408 41916
rect 4408 41860 4464 41916
rect 4464 41860 4468 41916
rect 4404 41856 4468 41860
rect 4484 41916 4548 41920
rect 4484 41860 4488 41916
rect 4488 41860 4544 41916
rect 4544 41860 4548 41916
rect 4484 41856 4548 41860
rect 4564 41916 4628 41920
rect 4564 41860 4568 41916
rect 4568 41860 4624 41916
rect 4624 41860 4628 41916
rect 4564 41856 4628 41860
rect 12098 41916 12162 41920
rect 12098 41860 12102 41916
rect 12102 41860 12158 41916
rect 12158 41860 12162 41916
rect 12098 41856 12162 41860
rect 12178 41916 12242 41920
rect 12178 41860 12182 41916
rect 12182 41860 12238 41916
rect 12238 41860 12242 41916
rect 12178 41856 12242 41860
rect 12258 41916 12322 41920
rect 12258 41860 12262 41916
rect 12262 41860 12318 41916
rect 12318 41860 12322 41916
rect 12258 41856 12322 41860
rect 12338 41916 12402 41920
rect 12338 41860 12342 41916
rect 12342 41860 12398 41916
rect 12398 41860 12402 41916
rect 12338 41856 12402 41860
rect 19872 41916 19936 41920
rect 19872 41860 19876 41916
rect 19876 41860 19932 41916
rect 19932 41860 19936 41916
rect 19872 41856 19936 41860
rect 19952 41916 20016 41920
rect 19952 41860 19956 41916
rect 19956 41860 20012 41916
rect 20012 41860 20016 41916
rect 19952 41856 20016 41860
rect 20032 41916 20096 41920
rect 20032 41860 20036 41916
rect 20036 41860 20092 41916
rect 20092 41860 20096 41916
rect 20032 41856 20096 41860
rect 20112 41916 20176 41920
rect 20112 41860 20116 41916
rect 20116 41860 20172 41916
rect 20172 41860 20176 41916
rect 20112 41856 20176 41860
rect 27646 41916 27710 41920
rect 27646 41860 27650 41916
rect 27650 41860 27706 41916
rect 27706 41860 27710 41916
rect 27646 41856 27710 41860
rect 27726 41916 27790 41920
rect 27726 41860 27730 41916
rect 27730 41860 27786 41916
rect 27786 41860 27790 41916
rect 27726 41856 27790 41860
rect 27806 41916 27870 41920
rect 27806 41860 27810 41916
rect 27810 41860 27866 41916
rect 27866 41860 27870 41916
rect 27806 41856 27870 41860
rect 27886 41916 27950 41920
rect 27886 41860 27890 41916
rect 27890 41860 27946 41916
rect 27946 41860 27950 41916
rect 27886 41856 27950 41860
rect 13676 41848 13740 41852
rect 13676 41792 13726 41848
rect 13726 41792 13740 41848
rect 13676 41788 13740 41792
rect 24532 41516 24596 41580
rect 3664 41372 3728 41376
rect 3664 41316 3668 41372
rect 3668 41316 3724 41372
rect 3724 41316 3728 41372
rect 3664 41312 3728 41316
rect 3744 41372 3808 41376
rect 3744 41316 3748 41372
rect 3748 41316 3804 41372
rect 3804 41316 3808 41372
rect 3744 41312 3808 41316
rect 3824 41372 3888 41376
rect 3824 41316 3828 41372
rect 3828 41316 3884 41372
rect 3884 41316 3888 41372
rect 3824 41312 3888 41316
rect 3904 41372 3968 41376
rect 3904 41316 3908 41372
rect 3908 41316 3964 41372
rect 3964 41316 3968 41372
rect 3904 41312 3968 41316
rect 11438 41372 11502 41376
rect 11438 41316 11442 41372
rect 11442 41316 11498 41372
rect 11498 41316 11502 41372
rect 11438 41312 11502 41316
rect 11518 41372 11582 41376
rect 11518 41316 11522 41372
rect 11522 41316 11578 41372
rect 11578 41316 11582 41372
rect 11518 41312 11582 41316
rect 11598 41372 11662 41376
rect 11598 41316 11602 41372
rect 11602 41316 11658 41372
rect 11658 41316 11662 41372
rect 11598 41312 11662 41316
rect 11678 41372 11742 41376
rect 11678 41316 11682 41372
rect 11682 41316 11738 41372
rect 11738 41316 11742 41372
rect 11678 41312 11742 41316
rect 19212 41372 19276 41376
rect 19212 41316 19216 41372
rect 19216 41316 19272 41372
rect 19272 41316 19276 41372
rect 19212 41312 19276 41316
rect 19292 41372 19356 41376
rect 19292 41316 19296 41372
rect 19296 41316 19352 41372
rect 19352 41316 19356 41372
rect 19292 41312 19356 41316
rect 19372 41372 19436 41376
rect 19372 41316 19376 41372
rect 19376 41316 19432 41372
rect 19432 41316 19436 41372
rect 19372 41312 19436 41316
rect 19452 41372 19516 41376
rect 19452 41316 19456 41372
rect 19456 41316 19512 41372
rect 19512 41316 19516 41372
rect 19452 41312 19516 41316
rect 26986 41372 27050 41376
rect 26986 41316 26990 41372
rect 26990 41316 27046 41372
rect 27046 41316 27050 41372
rect 26986 41312 27050 41316
rect 27066 41372 27130 41376
rect 27066 41316 27070 41372
rect 27070 41316 27126 41372
rect 27126 41316 27130 41372
rect 27066 41312 27130 41316
rect 27146 41372 27210 41376
rect 27146 41316 27150 41372
rect 27150 41316 27206 41372
rect 27206 41316 27210 41372
rect 27146 41312 27210 41316
rect 27226 41372 27290 41376
rect 27226 41316 27230 41372
rect 27230 41316 27286 41372
rect 27286 41316 27290 41372
rect 27226 41312 27290 41316
rect 16068 41108 16132 41172
rect 4324 40828 4388 40832
rect 4324 40772 4328 40828
rect 4328 40772 4384 40828
rect 4384 40772 4388 40828
rect 4324 40768 4388 40772
rect 4404 40828 4468 40832
rect 4404 40772 4408 40828
rect 4408 40772 4464 40828
rect 4464 40772 4468 40828
rect 4404 40768 4468 40772
rect 4484 40828 4548 40832
rect 4484 40772 4488 40828
rect 4488 40772 4544 40828
rect 4544 40772 4548 40828
rect 4484 40768 4548 40772
rect 4564 40828 4628 40832
rect 4564 40772 4568 40828
rect 4568 40772 4624 40828
rect 4624 40772 4628 40828
rect 4564 40768 4628 40772
rect 12098 40828 12162 40832
rect 12098 40772 12102 40828
rect 12102 40772 12158 40828
rect 12158 40772 12162 40828
rect 12098 40768 12162 40772
rect 12178 40828 12242 40832
rect 12178 40772 12182 40828
rect 12182 40772 12238 40828
rect 12238 40772 12242 40828
rect 12178 40768 12242 40772
rect 12258 40828 12322 40832
rect 12258 40772 12262 40828
rect 12262 40772 12318 40828
rect 12318 40772 12322 40828
rect 12258 40768 12322 40772
rect 12338 40828 12402 40832
rect 12338 40772 12342 40828
rect 12342 40772 12398 40828
rect 12398 40772 12402 40828
rect 12338 40768 12402 40772
rect 19872 40828 19936 40832
rect 19872 40772 19876 40828
rect 19876 40772 19932 40828
rect 19932 40772 19936 40828
rect 19872 40768 19936 40772
rect 19952 40828 20016 40832
rect 19952 40772 19956 40828
rect 19956 40772 20012 40828
rect 20012 40772 20016 40828
rect 19952 40768 20016 40772
rect 20032 40828 20096 40832
rect 20032 40772 20036 40828
rect 20036 40772 20092 40828
rect 20092 40772 20096 40828
rect 20032 40768 20096 40772
rect 20112 40828 20176 40832
rect 20112 40772 20116 40828
rect 20116 40772 20172 40828
rect 20172 40772 20176 40828
rect 20112 40768 20176 40772
rect 27646 40828 27710 40832
rect 27646 40772 27650 40828
rect 27650 40772 27706 40828
rect 27706 40772 27710 40828
rect 27646 40768 27710 40772
rect 27726 40828 27790 40832
rect 27726 40772 27730 40828
rect 27730 40772 27786 40828
rect 27786 40772 27790 40828
rect 27726 40768 27790 40772
rect 27806 40828 27870 40832
rect 27806 40772 27810 40828
rect 27810 40772 27866 40828
rect 27866 40772 27870 40828
rect 27806 40768 27870 40772
rect 27886 40828 27950 40832
rect 27886 40772 27890 40828
rect 27890 40772 27946 40828
rect 27946 40772 27950 40828
rect 27886 40768 27950 40772
rect 3664 40284 3728 40288
rect 3664 40228 3668 40284
rect 3668 40228 3724 40284
rect 3724 40228 3728 40284
rect 3664 40224 3728 40228
rect 3744 40284 3808 40288
rect 3744 40228 3748 40284
rect 3748 40228 3804 40284
rect 3804 40228 3808 40284
rect 3744 40224 3808 40228
rect 3824 40284 3888 40288
rect 3824 40228 3828 40284
rect 3828 40228 3884 40284
rect 3884 40228 3888 40284
rect 3824 40224 3888 40228
rect 3904 40284 3968 40288
rect 3904 40228 3908 40284
rect 3908 40228 3964 40284
rect 3964 40228 3968 40284
rect 3904 40224 3968 40228
rect 11438 40284 11502 40288
rect 11438 40228 11442 40284
rect 11442 40228 11498 40284
rect 11498 40228 11502 40284
rect 11438 40224 11502 40228
rect 11518 40284 11582 40288
rect 11518 40228 11522 40284
rect 11522 40228 11578 40284
rect 11578 40228 11582 40284
rect 11518 40224 11582 40228
rect 11598 40284 11662 40288
rect 11598 40228 11602 40284
rect 11602 40228 11658 40284
rect 11658 40228 11662 40284
rect 11598 40224 11662 40228
rect 11678 40284 11742 40288
rect 11678 40228 11682 40284
rect 11682 40228 11738 40284
rect 11738 40228 11742 40284
rect 11678 40224 11742 40228
rect 19212 40284 19276 40288
rect 19212 40228 19216 40284
rect 19216 40228 19272 40284
rect 19272 40228 19276 40284
rect 19212 40224 19276 40228
rect 19292 40284 19356 40288
rect 19292 40228 19296 40284
rect 19296 40228 19352 40284
rect 19352 40228 19356 40284
rect 19292 40224 19356 40228
rect 19372 40284 19436 40288
rect 19372 40228 19376 40284
rect 19376 40228 19432 40284
rect 19432 40228 19436 40284
rect 19372 40224 19436 40228
rect 19452 40284 19516 40288
rect 19452 40228 19456 40284
rect 19456 40228 19512 40284
rect 19512 40228 19516 40284
rect 19452 40224 19516 40228
rect 26986 40284 27050 40288
rect 26986 40228 26990 40284
rect 26990 40228 27046 40284
rect 27046 40228 27050 40284
rect 26986 40224 27050 40228
rect 27066 40284 27130 40288
rect 27066 40228 27070 40284
rect 27070 40228 27126 40284
rect 27126 40228 27130 40284
rect 27066 40224 27130 40228
rect 27146 40284 27210 40288
rect 27146 40228 27150 40284
rect 27150 40228 27206 40284
rect 27206 40228 27210 40284
rect 27146 40224 27210 40228
rect 27226 40284 27290 40288
rect 27226 40228 27230 40284
rect 27230 40228 27286 40284
rect 27286 40228 27290 40284
rect 27226 40224 27290 40228
rect 4324 39740 4388 39744
rect 4324 39684 4328 39740
rect 4328 39684 4384 39740
rect 4384 39684 4388 39740
rect 4324 39680 4388 39684
rect 4404 39740 4468 39744
rect 4404 39684 4408 39740
rect 4408 39684 4464 39740
rect 4464 39684 4468 39740
rect 4404 39680 4468 39684
rect 4484 39740 4548 39744
rect 4484 39684 4488 39740
rect 4488 39684 4544 39740
rect 4544 39684 4548 39740
rect 4484 39680 4548 39684
rect 4564 39740 4628 39744
rect 4564 39684 4568 39740
rect 4568 39684 4624 39740
rect 4624 39684 4628 39740
rect 4564 39680 4628 39684
rect 12098 39740 12162 39744
rect 12098 39684 12102 39740
rect 12102 39684 12158 39740
rect 12158 39684 12162 39740
rect 12098 39680 12162 39684
rect 12178 39740 12242 39744
rect 12178 39684 12182 39740
rect 12182 39684 12238 39740
rect 12238 39684 12242 39740
rect 12178 39680 12242 39684
rect 12258 39740 12322 39744
rect 12258 39684 12262 39740
rect 12262 39684 12318 39740
rect 12318 39684 12322 39740
rect 12258 39680 12322 39684
rect 12338 39740 12402 39744
rect 12338 39684 12342 39740
rect 12342 39684 12398 39740
rect 12398 39684 12402 39740
rect 12338 39680 12402 39684
rect 19872 39740 19936 39744
rect 19872 39684 19876 39740
rect 19876 39684 19932 39740
rect 19932 39684 19936 39740
rect 19872 39680 19936 39684
rect 19952 39740 20016 39744
rect 19952 39684 19956 39740
rect 19956 39684 20012 39740
rect 20012 39684 20016 39740
rect 19952 39680 20016 39684
rect 20032 39740 20096 39744
rect 20032 39684 20036 39740
rect 20036 39684 20092 39740
rect 20092 39684 20096 39740
rect 20032 39680 20096 39684
rect 20112 39740 20176 39744
rect 20112 39684 20116 39740
rect 20116 39684 20172 39740
rect 20172 39684 20176 39740
rect 20112 39680 20176 39684
rect 27646 39740 27710 39744
rect 27646 39684 27650 39740
rect 27650 39684 27706 39740
rect 27706 39684 27710 39740
rect 27646 39680 27710 39684
rect 27726 39740 27790 39744
rect 27726 39684 27730 39740
rect 27730 39684 27786 39740
rect 27786 39684 27790 39740
rect 27726 39680 27790 39684
rect 27806 39740 27870 39744
rect 27806 39684 27810 39740
rect 27810 39684 27866 39740
rect 27866 39684 27870 39740
rect 27806 39680 27870 39684
rect 27886 39740 27950 39744
rect 27886 39684 27890 39740
rect 27890 39684 27946 39740
rect 27946 39684 27950 39740
rect 27886 39680 27950 39684
rect 20484 39340 20548 39404
rect 3664 39196 3728 39200
rect 3664 39140 3668 39196
rect 3668 39140 3724 39196
rect 3724 39140 3728 39196
rect 3664 39136 3728 39140
rect 3744 39196 3808 39200
rect 3744 39140 3748 39196
rect 3748 39140 3804 39196
rect 3804 39140 3808 39196
rect 3744 39136 3808 39140
rect 3824 39196 3888 39200
rect 3824 39140 3828 39196
rect 3828 39140 3884 39196
rect 3884 39140 3888 39196
rect 3824 39136 3888 39140
rect 3904 39196 3968 39200
rect 3904 39140 3908 39196
rect 3908 39140 3964 39196
rect 3964 39140 3968 39196
rect 3904 39136 3968 39140
rect 11438 39196 11502 39200
rect 11438 39140 11442 39196
rect 11442 39140 11498 39196
rect 11498 39140 11502 39196
rect 11438 39136 11502 39140
rect 11518 39196 11582 39200
rect 11518 39140 11522 39196
rect 11522 39140 11578 39196
rect 11578 39140 11582 39196
rect 11518 39136 11582 39140
rect 11598 39196 11662 39200
rect 11598 39140 11602 39196
rect 11602 39140 11658 39196
rect 11658 39140 11662 39196
rect 11598 39136 11662 39140
rect 11678 39196 11742 39200
rect 11678 39140 11682 39196
rect 11682 39140 11738 39196
rect 11738 39140 11742 39196
rect 11678 39136 11742 39140
rect 19212 39196 19276 39200
rect 19212 39140 19216 39196
rect 19216 39140 19272 39196
rect 19272 39140 19276 39196
rect 19212 39136 19276 39140
rect 19292 39196 19356 39200
rect 19292 39140 19296 39196
rect 19296 39140 19352 39196
rect 19352 39140 19356 39196
rect 19292 39136 19356 39140
rect 19372 39196 19436 39200
rect 19372 39140 19376 39196
rect 19376 39140 19432 39196
rect 19432 39140 19436 39196
rect 19372 39136 19436 39140
rect 19452 39196 19516 39200
rect 19452 39140 19456 39196
rect 19456 39140 19512 39196
rect 19512 39140 19516 39196
rect 19452 39136 19516 39140
rect 26986 39196 27050 39200
rect 26986 39140 26990 39196
rect 26990 39140 27046 39196
rect 27046 39140 27050 39196
rect 26986 39136 27050 39140
rect 27066 39196 27130 39200
rect 27066 39140 27070 39196
rect 27070 39140 27126 39196
rect 27126 39140 27130 39196
rect 27066 39136 27130 39140
rect 27146 39196 27210 39200
rect 27146 39140 27150 39196
rect 27150 39140 27206 39196
rect 27206 39140 27210 39196
rect 27146 39136 27210 39140
rect 27226 39196 27290 39200
rect 27226 39140 27230 39196
rect 27230 39140 27286 39196
rect 27286 39140 27290 39196
rect 27226 39136 27290 39140
rect 20300 38796 20364 38860
rect 4324 38652 4388 38656
rect 4324 38596 4328 38652
rect 4328 38596 4384 38652
rect 4384 38596 4388 38652
rect 4324 38592 4388 38596
rect 4404 38652 4468 38656
rect 4404 38596 4408 38652
rect 4408 38596 4464 38652
rect 4464 38596 4468 38652
rect 4404 38592 4468 38596
rect 4484 38652 4548 38656
rect 4484 38596 4488 38652
rect 4488 38596 4544 38652
rect 4544 38596 4548 38652
rect 4484 38592 4548 38596
rect 4564 38652 4628 38656
rect 4564 38596 4568 38652
rect 4568 38596 4624 38652
rect 4624 38596 4628 38652
rect 4564 38592 4628 38596
rect 12098 38652 12162 38656
rect 12098 38596 12102 38652
rect 12102 38596 12158 38652
rect 12158 38596 12162 38652
rect 12098 38592 12162 38596
rect 12178 38652 12242 38656
rect 12178 38596 12182 38652
rect 12182 38596 12238 38652
rect 12238 38596 12242 38652
rect 12178 38592 12242 38596
rect 12258 38652 12322 38656
rect 12258 38596 12262 38652
rect 12262 38596 12318 38652
rect 12318 38596 12322 38652
rect 12258 38592 12322 38596
rect 12338 38652 12402 38656
rect 12338 38596 12342 38652
rect 12342 38596 12398 38652
rect 12398 38596 12402 38652
rect 12338 38592 12402 38596
rect 19872 38652 19936 38656
rect 19872 38596 19876 38652
rect 19876 38596 19932 38652
rect 19932 38596 19936 38652
rect 19872 38592 19936 38596
rect 19952 38652 20016 38656
rect 19952 38596 19956 38652
rect 19956 38596 20012 38652
rect 20012 38596 20016 38652
rect 19952 38592 20016 38596
rect 20032 38652 20096 38656
rect 20032 38596 20036 38652
rect 20036 38596 20092 38652
rect 20092 38596 20096 38652
rect 20032 38592 20096 38596
rect 20112 38652 20176 38656
rect 20112 38596 20116 38652
rect 20116 38596 20172 38652
rect 20172 38596 20176 38652
rect 20112 38592 20176 38596
rect 27646 38652 27710 38656
rect 27646 38596 27650 38652
rect 27650 38596 27706 38652
rect 27706 38596 27710 38652
rect 27646 38592 27710 38596
rect 27726 38652 27790 38656
rect 27726 38596 27730 38652
rect 27730 38596 27786 38652
rect 27786 38596 27790 38652
rect 27726 38592 27790 38596
rect 27806 38652 27870 38656
rect 27806 38596 27810 38652
rect 27810 38596 27866 38652
rect 27866 38596 27870 38652
rect 27806 38592 27870 38596
rect 27886 38652 27950 38656
rect 27886 38596 27890 38652
rect 27890 38596 27946 38652
rect 27946 38596 27950 38652
rect 27886 38592 27950 38596
rect 3664 38108 3728 38112
rect 3664 38052 3668 38108
rect 3668 38052 3724 38108
rect 3724 38052 3728 38108
rect 3664 38048 3728 38052
rect 3744 38108 3808 38112
rect 3744 38052 3748 38108
rect 3748 38052 3804 38108
rect 3804 38052 3808 38108
rect 3744 38048 3808 38052
rect 3824 38108 3888 38112
rect 3824 38052 3828 38108
rect 3828 38052 3884 38108
rect 3884 38052 3888 38108
rect 3824 38048 3888 38052
rect 3904 38108 3968 38112
rect 3904 38052 3908 38108
rect 3908 38052 3964 38108
rect 3964 38052 3968 38108
rect 3904 38048 3968 38052
rect 11438 38108 11502 38112
rect 11438 38052 11442 38108
rect 11442 38052 11498 38108
rect 11498 38052 11502 38108
rect 11438 38048 11502 38052
rect 11518 38108 11582 38112
rect 11518 38052 11522 38108
rect 11522 38052 11578 38108
rect 11578 38052 11582 38108
rect 11518 38048 11582 38052
rect 11598 38108 11662 38112
rect 11598 38052 11602 38108
rect 11602 38052 11658 38108
rect 11658 38052 11662 38108
rect 11598 38048 11662 38052
rect 11678 38108 11742 38112
rect 11678 38052 11682 38108
rect 11682 38052 11738 38108
rect 11738 38052 11742 38108
rect 11678 38048 11742 38052
rect 19212 38108 19276 38112
rect 19212 38052 19216 38108
rect 19216 38052 19272 38108
rect 19272 38052 19276 38108
rect 19212 38048 19276 38052
rect 19292 38108 19356 38112
rect 19292 38052 19296 38108
rect 19296 38052 19352 38108
rect 19352 38052 19356 38108
rect 19292 38048 19356 38052
rect 19372 38108 19436 38112
rect 19372 38052 19376 38108
rect 19376 38052 19432 38108
rect 19432 38052 19436 38108
rect 19372 38048 19436 38052
rect 19452 38108 19516 38112
rect 19452 38052 19456 38108
rect 19456 38052 19512 38108
rect 19512 38052 19516 38108
rect 19452 38048 19516 38052
rect 26986 38108 27050 38112
rect 26986 38052 26990 38108
rect 26990 38052 27046 38108
rect 27046 38052 27050 38108
rect 26986 38048 27050 38052
rect 27066 38108 27130 38112
rect 27066 38052 27070 38108
rect 27070 38052 27126 38108
rect 27126 38052 27130 38108
rect 27066 38048 27130 38052
rect 27146 38108 27210 38112
rect 27146 38052 27150 38108
rect 27150 38052 27206 38108
rect 27206 38052 27210 38108
rect 27146 38048 27210 38052
rect 27226 38108 27290 38112
rect 27226 38052 27230 38108
rect 27230 38052 27286 38108
rect 27286 38052 27290 38108
rect 27226 38048 27290 38052
rect 20300 37708 20364 37772
rect 4324 37564 4388 37568
rect 4324 37508 4328 37564
rect 4328 37508 4384 37564
rect 4384 37508 4388 37564
rect 4324 37504 4388 37508
rect 4404 37564 4468 37568
rect 4404 37508 4408 37564
rect 4408 37508 4464 37564
rect 4464 37508 4468 37564
rect 4404 37504 4468 37508
rect 4484 37564 4548 37568
rect 4484 37508 4488 37564
rect 4488 37508 4544 37564
rect 4544 37508 4548 37564
rect 4484 37504 4548 37508
rect 4564 37564 4628 37568
rect 4564 37508 4568 37564
rect 4568 37508 4624 37564
rect 4624 37508 4628 37564
rect 4564 37504 4628 37508
rect 12098 37564 12162 37568
rect 12098 37508 12102 37564
rect 12102 37508 12158 37564
rect 12158 37508 12162 37564
rect 12098 37504 12162 37508
rect 12178 37564 12242 37568
rect 12178 37508 12182 37564
rect 12182 37508 12238 37564
rect 12238 37508 12242 37564
rect 12178 37504 12242 37508
rect 12258 37564 12322 37568
rect 12258 37508 12262 37564
rect 12262 37508 12318 37564
rect 12318 37508 12322 37564
rect 12258 37504 12322 37508
rect 12338 37564 12402 37568
rect 12338 37508 12342 37564
rect 12342 37508 12398 37564
rect 12398 37508 12402 37564
rect 12338 37504 12402 37508
rect 19872 37564 19936 37568
rect 19872 37508 19876 37564
rect 19876 37508 19932 37564
rect 19932 37508 19936 37564
rect 19872 37504 19936 37508
rect 19952 37564 20016 37568
rect 19952 37508 19956 37564
rect 19956 37508 20012 37564
rect 20012 37508 20016 37564
rect 19952 37504 20016 37508
rect 20032 37564 20096 37568
rect 20032 37508 20036 37564
rect 20036 37508 20092 37564
rect 20092 37508 20096 37564
rect 20032 37504 20096 37508
rect 20112 37564 20176 37568
rect 20112 37508 20116 37564
rect 20116 37508 20172 37564
rect 20172 37508 20176 37564
rect 20112 37504 20176 37508
rect 27646 37564 27710 37568
rect 27646 37508 27650 37564
rect 27650 37508 27706 37564
rect 27706 37508 27710 37564
rect 27646 37504 27710 37508
rect 27726 37564 27790 37568
rect 27726 37508 27730 37564
rect 27730 37508 27786 37564
rect 27786 37508 27790 37564
rect 27726 37504 27790 37508
rect 27806 37564 27870 37568
rect 27806 37508 27810 37564
rect 27810 37508 27866 37564
rect 27866 37508 27870 37564
rect 27806 37504 27870 37508
rect 27886 37564 27950 37568
rect 27886 37508 27890 37564
rect 27890 37508 27946 37564
rect 27946 37508 27950 37564
rect 27886 37504 27950 37508
rect 20668 37164 20732 37228
rect 3664 37020 3728 37024
rect 3664 36964 3668 37020
rect 3668 36964 3724 37020
rect 3724 36964 3728 37020
rect 3664 36960 3728 36964
rect 3744 37020 3808 37024
rect 3744 36964 3748 37020
rect 3748 36964 3804 37020
rect 3804 36964 3808 37020
rect 3744 36960 3808 36964
rect 3824 37020 3888 37024
rect 3824 36964 3828 37020
rect 3828 36964 3884 37020
rect 3884 36964 3888 37020
rect 3824 36960 3888 36964
rect 3904 37020 3968 37024
rect 3904 36964 3908 37020
rect 3908 36964 3964 37020
rect 3964 36964 3968 37020
rect 3904 36960 3968 36964
rect 11438 37020 11502 37024
rect 11438 36964 11442 37020
rect 11442 36964 11498 37020
rect 11498 36964 11502 37020
rect 11438 36960 11502 36964
rect 11518 37020 11582 37024
rect 11518 36964 11522 37020
rect 11522 36964 11578 37020
rect 11578 36964 11582 37020
rect 11518 36960 11582 36964
rect 11598 37020 11662 37024
rect 11598 36964 11602 37020
rect 11602 36964 11658 37020
rect 11658 36964 11662 37020
rect 11598 36960 11662 36964
rect 11678 37020 11742 37024
rect 11678 36964 11682 37020
rect 11682 36964 11738 37020
rect 11738 36964 11742 37020
rect 11678 36960 11742 36964
rect 19212 37020 19276 37024
rect 19212 36964 19216 37020
rect 19216 36964 19272 37020
rect 19272 36964 19276 37020
rect 19212 36960 19276 36964
rect 19292 37020 19356 37024
rect 19292 36964 19296 37020
rect 19296 36964 19352 37020
rect 19352 36964 19356 37020
rect 19292 36960 19356 36964
rect 19372 37020 19436 37024
rect 19372 36964 19376 37020
rect 19376 36964 19432 37020
rect 19432 36964 19436 37020
rect 19372 36960 19436 36964
rect 19452 37020 19516 37024
rect 19452 36964 19456 37020
rect 19456 36964 19512 37020
rect 19512 36964 19516 37020
rect 19452 36960 19516 36964
rect 26986 37020 27050 37024
rect 26986 36964 26990 37020
rect 26990 36964 27046 37020
rect 27046 36964 27050 37020
rect 26986 36960 27050 36964
rect 27066 37020 27130 37024
rect 27066 36964 27070 37020
rect 27070 36964 27126 37020
rect 27126 36964 27130 37020
rect 27066 36960 27130 36964
rect 27146 37020 27210 37024
rect 27146 36964 27150 37020
rect 27150 36964 27206 37020
rect 27206 36964 27210 37020
rect 27146 36960 27210 36964
rect 27226 37020 27290 37024
rect 27226 36964 27230 37020
rect 27230 36964 27286 37020
rect 27286 36964 27290 37020
rect 27226 36960 27290 36964
rect 20300 36756 20364 36820
rect 21956 36680 22020 36684
rect 21956 36624 21970 36680
rect 21970 36624 22020 36680
rect 21956 36620 22020 36624
rect 4324 36476 4388 36480
rect 4324 36420 4328 36476
rect 4328 36420 4384 36476
rect 4384 36420 4388 36476
rect 4324 36416 4388 36420
rect 4404 36476 4468 36480
rect 4404 36420 4408 36476
rect 4408 36420 4464 36476
rect 4464 36420 4468 36476
rect 4404 36416 4468 36420
rect 4484 36476 4548 36480
rect 4484 36420 4488 36476
rect 4488 36420 4544 36476
rect 4544 36420 4548 36476
rect 4484 36416 4548 36420
rect 4564 36476 4628 36480
rect 4564 36420 4568 36476
rect 4568 36420 4624 36476
rect 4624 36420 4628 36476
rect 4564 36416 4628 36420
rect 12098 36476 12162 36480
rect 12098 36420 12102 36476
rect 12102 36420 12158 36476
rect 12158 36420 12162 36476
rect 12098 36416 12162 36420
rect 12178 36476 12242 36480
rect 12178 36420 12182 36476
rect 12182 36420 12238 36476
rect 12238 36420 12242 36476
rect 12178 36416 12242 36420
rect 12258 36476 12322 36480
rect 12258 36420 12262 36476
rect 12262 36420 12318 36476
rect 12318 36420 12322 36476
rect 12258 36416 12322 36420
rect 12338 36476 12402 36480
rect 12338 36420 12342 36476
rect 12342 36420 12398 36476
rect 12398 36420 12402 36476
rect 12338 36416 12402 36420
rect 19872 36476 19936 36480
rect 19872 36420 19876 36476
rect 19876 36420 19932 36476
rect 19932 36420 19936 36476
rect 19872 36416 19936 36420
rect 19952 36476 20016 36480
rect 19952 36420 19956 36476
rect 19956 36420 20012 36476
rect 20012 36420 20016 36476
rect 19952 36416 20016 36420
rect 20032 36476 20096 36480
rect 20032 36420 20036 36476
rect 20036 36420 20092 36476
rect 20092 36420 20096 36476
rect 20032 36416 20096 36420
rect 20112 36476 20176 36480
rect 20112 36420 20116 36476
rect 20116 36420 20172 36476
rect 20172 36420 20176 36476
rect 20112 36416 20176 36420
rect 27646 36476 27710 36480
rect 27646 36420 27650 36476
rect 27650 36420 27706 36476
rect 27706 36420 27710 36476
rect 27646 36416 27710 36420
rect 27726 36476 27790 36480
rect 27726 36420 27730 36476
rect 27730 36420 27786 36476
rect 27786 36420 27790 36476
rect 27726 36416 27790 36420
rect 27806 36476 27870 36480
rect 27806 36420 27810 36476
rect 27810 36420 27866 36476
rect 27866 36420 27870 36476
rect 27806 36416 27870 36420
rect 27886 36476 27950 36480
rect 27886 36420 27890 36476
rect 27890 36420 27946 36476
rect 27946 36420 27950 36476
rect 27886 36416 27950 36420
rect 10548 36076 10612 36140
rect 18460 35940 18524 36004
rect 3664 35932 3728 35936
rect 3664 35876 3668 35932
rect 3668 35876 3724 35932
rect 3724 35876 3728 35932
rect 3664 35872 3728 35876
rect 3744 35932 3808 35936
rect 3744 35876 3748 35932
rect 3748 35876 3804 35932
rect 3804 35876 3808 35932
rect 3744 35872 3808 35876
rect 3824 35932 3888 35936
rect 3824 35876 3828 35932
rect 3828 35876 3884 35932
rect 3884 35876 3888 35932
rect 3824 35872 3888 35876
rect 3904 35932 3968 35936
rect 3904 35876 3908 35932
rect 3908 35876 3964 35932
rect 3964 35876 3968 35932
rect 3904 35872 3968 35876
rect 11438 35932 11502 35936
rect 11438 35876 11442 35932
rect 11442 35876 11498 35932
rect 11498 35876 11502 35932
rect 11438 35872 11502 35876
rect 11518 35932 11582 35936
rect 11518 35876 11522 35932
rect 11522 35876 11578 35932
rect 11578 35876 11582 35932
rect 11518 35872 11582 35876
rect 11598 35932 11662 35936
rect 11598 35876 11602 35932
rect 11602 35876 11658 35932
rect 11658 35876 11662 35932
rect 11598 35872 11662 35876
rect 11678 35932 11742 35936
rect 11678 35876 11682 35932
rect 11682 35876 11738 35932
rect 11738 35876 11742 35932
rect 11678 35872 11742 35876
rect 19212 35932 19276 35936
rect 19212 35876 19216 35932
rect 19216 35876 19272 35932
rect 19272 35876 19276 35932
rect 19212 35872 19276 35876
rect 19292 35932 19356 35936
rect 19292 35876 19296 35932
rect 19296 35876 19352 35932
rect 19352 35876 19356 35932
rect 19292 35872 19356 35876
rect 19372 35932 19436 35936
rect 19372 35876 19376 35932
rect 19376 35876 19432 35932
rect 19432 35876 19436 35932
rect 19372 35872 19436 35876
rect 19452 35932 19516 35936
rect 19452 35876 19456 35932
rect 19456 35876 19512 35932
rect 19512 35876 19516 35932
rect 19452 35872 19516 35876
rect 26986 35932 27050 35936
rect 26986 35876 26990 35932
rect 26990 35876 27046 35932
rect 27046 35876 27050 35932
rect 26986 35872 27050 35876
rect 27066 35932 27130 35936
rect 27066 35876 27070 35932
rect 27070 35876 27126 35932
rect 27126 35876 27130 35932
rect 27066 35872 27130 35876
rect 27146 35932 27210 35936
rect 27146 35876 27150 35932
rect 27150 35876 27206 35932
rect 27206 35876 27210 35932
rect 27146 35872 27210 35876
rect 27226 35932 27290 35936
rect 27226 35876 27230 35932
rect 27230 35876 27286 35932
rect 27286 35876 27290 35932
rect 27226 35872 27290 35876
rect 4324 35388 4388 35392
rect 4324 35332 4328 35388
rect 4328 35332 4384 35388
rect 4384 35332 4388 35388
rect 4324 35328 4388 35332
rect 4404 35388 4468 35392
rect 4404 35332 4408 35388
rect 4408 35332 4464 35388
rect 4464 35332 4468 35388
rect 4404 35328 4468 35332
rect 4484 35388 4548 35392
rect 4484 35332 4488 35388
rect 4488 35332 4544 35388
rect 4544 35332 4548 35388
rect 4484 35328 4548 35332
rect 4564 35388 4628 35392
rect 4564 35332 4568 35388
rect 4568 35332 4624 35388
rect 4624 35332 4628 35388
rect 4564 35328 4628 35332
rect 12098 35388 12162 35392
rect 12098 35332 12102 35388
rect 12102 35332 12158 35388
rect 12158 35332 12162 35388
rect 12098 35328 12162 35332
rect 12178 35388 12242 35392
rect 12178 35332 12182 35388
rect 12182 35332 12238 35388
rect 12238 35332 12242 35388
rect 12178 35328 12242 35332
rect 12258 35388 12322 35392
rect 12258 35332 12262 35388
rect 12262 35332 12318 35388
rect 12318 35332 12322 35388
rect 12258 35328 12322 35332
rect 12338 35388 12402 35392
rect 12338 35332 12342 35388
rect 12342 35332 12398 35388
rect 12398 35332 12402 35388
rect 12338 35328 12402 35332
rect 19872 35388 19936 35392
rect 19872 35332 19876 35388
rect 19876 35332 19932 35388
rect 19932 35332 19936 35388
rect 19872 35328 19936 35332
rect 19952 35388 20016 35392
rect 19952 35332 19956 35388
rect 19956 35332 20012 35388
rect 20012 35332 20016 35388
rect 19952 35328 20016 35332
rect 20032 35388 20096 35392
rect 20032 35332 20036 35388
rect 20036 35332 20092 35388
rect 20092 35332 20096 35388
rect 20032 35328 20096 35332
rect 20112 35388 20176 35392
rect 20112 35332 20116 35388
rect 20116 35332 20172 35388
rect 20172 35332 20176 35388
rect 20112 35328 20176 35332
rect 27646 35388 27710 35392
rect 27646 35332 27650 35388
rect 27650 35332 27706 35388
rect 27706 35332 27710 35388
rect 27646 35328 27710 35332
rect 27726 35388 27790 35392
rect 27726 35332 27730 35388
rect 27730 35332 27786 35388
rect 27786 35332 27790 35388
rect 27726 35328 27790 35332
rect 27806 35388 27870 35392
rect 27806 35332 27810 35388
rect 27810 35332 27866 35388
rect 27866 35332 27870 35388
rect 27806 35328 27870 35332
rect 27886 35388 27950 35392
rect 27886 35332 27890 35388
rect 27890 35332 27946 35388
rect 27946 35332 27950 35388
rect 27886 35328 27950 35332
rect 3664 34844 3728 34848
rect 3664 34788 3668 34844
rect 3668 34788 3724 34844
rect 3724 34788 3728 34844
rect 3664 34784 3728 34788
rect 3744 34844 3808 34848
rect 3744 34788 3748 34844
rect 3748 34788 3804 34844
rect 3804 34788 3808 34844
rect 3744 34784 3808 34788
rect 3824 34844 3888 34848
rect 3824 34788 3828 34844
rect 3828 34788 3884 34844
rect 3884 34788 3888 34844
rect 3824 34784 3888 34788
rect 3904 34844 3968 34848
rect 3904 34788 3908 34844
rect 3908 34788 3964 34844
rect 3964 34788 3968 34844
rect 3904 34784 3968 34788
rect 11438 34844 11502 34848
rect 11438 34788 11442 34844
rect 11442 34788 11498 34844
rect 11498 34788 11502 34844
rect 11438 34784 11502 34788
rect 11518 34844 11582 34848
rect 11518 34788 11522 34844
rect 11522 34788 11578 34844
rect 11578 34788 11582 34844
rect 11518 34784 11582 34788
rect 11598 34844 11662 34848
rect 11598 34788 11602 34844
rect 11602 34788 11658 34844
rect 11658 34788 11662 34844
rect 11598 34784 11662 34788
rect 11678 34844 11742 34848
rect 11678 34788 11682 34844
rect 11682 34788 11738 34844
rect 11738 34788 11742 34844
rect 11678 34784 11742 34788
rect 19212 34844 19276 34848
rect 19212 34788 19216 34844
rect 19216 34788 19272 34844
rect 19272 34788 19276 34844
rect 19212 34784 19276 34788
rect 19292 34844 19356 34848
rect 19292 34788 19296 34844
rect 19296 34788 19352 34844
rect 19352 34788 19356 34844
rect 19292 34784 19356 34788
rect 19372 34844 19436 34848
rect 19372 34788 19376 34844
rect 19376 34788 19432 34844
rect 19432 34788 19436 34844
rect 19372 34784 19436 34788
rect 19452 34844 19516 34848
rect 19452 34788 19456 34844
rect 19456 34788 19512 34844
rect 19512 34788 19516 34844
rect 19452 34784 19516 34788
rect 26986 34844 27050 34848
rect 26986 34788 26990 34844
rect 26990 34788 27046 34844
rect 27046 34788 27050 34844
rect 26986 34784 27050 34788
rect 27066 34844 27130 34848
rect 27066 34788 27070 34844
rect 27070 34788 27126 34844
rect 27126 34788 27130 34844
rect 27066 34784 27130 34788
rect 27146 34844 27210 34848
rect 27146 34788 27150 34844
rect 27150 34788 27206 34844
rect 27206 34788 27210 34844
rect 27146 34784 27210 34788
rect 27226 34844 27290 34848
rect 27226 34788 27230 34844
rect 27230 34788 27286 34844
rect 27286 34788 27290 34844
rect 27226 34784 27290 34788
rect 4324 34300 4388 34304
rect 4324 34244 4328 34300
rect 4328 34244 4384 34300
rect 4384 34244 4388 34300
rect 4324 34240 4388 34244
rect 4404 34300 4468 34304
rect 4404 34244 4408 34300
rect 4408 34244 4464 34300
rect 4464 34244 4468 34300
rect 4404 34240 4468 34244
rect 4484 34300 4548 34304
rect 4484 34244 4488 34300
rect 4488 34244 4544 34300
rect 4544 34244 4548 34300
rect 4484 34240 4548 34244
rect 4564 34300 4628 34304
rect 4564 34244 4568 34300
rect 4568 34244 4624 34300
rect 4624 34244 4628 34300
rect 4564 34240 4628 34244
rect 12098 34300 12162 34304
rect 12098 34244 12102 34300
rect 12102 34244 12158 34300
rect 12158 34244 12162 34300
rect 12098 34240 12162 34244
rect 12178 34300 12242 34304
rect 12178 34244 12182 34300
rect 12182 34244 12238 34300
rect 12238 34244 12242 34300
rect 12178 34240 12242 34244
rect 12258 34300 12322 34304
rect 12258 34244 12262 34300
rect 12262 34244 12318 34300
rect 12318 34244 12322 34300
rect 12258 34240 12322 34244
rect 12338 34300 12402 34304
rect 12338 34244 12342 34300
rect 12342 34244 12398 34300
rect 12398 34244 12402 34300
rect 12338 34240 12402 34244
rect 19872 34300 19936 34304
rect 19872 34244 19876 34300
rect 19876 34244 19932 34300
rect 19932 34244 19936 34300
rect 19872 34240 19936 34244
rect 19952 34300 20016 34304
rect 19952 34244 19956 34300
rect 19956 34244 20012 34300
rect 20012 34244 20016 34300
rect 19952 34240 20016 34244
rect 20032 34300 20096 34304
rect 20032 34244 20036 34300
rect 20036 34244 20092 34300
rect 20092 34244 20096 34300
rect 20032 34240 20096 34244
rect 20112 34300 20176 34304
rect 20112 34244 20116 34300
rect 20116 34244 20172 34300
rect 20172 34244 20176 34300
rect 20112 34240 20176 34244
rect 27646 34300 27710 34304
rect 27646 34244 27650 34300
rect 27650 34244 27706 34300
rect 27706 34244 27710 34300
rect 27646 34240 27710 34244
rect 27726 34300 27790 34304
rect 27726 34244 27730 34300
rect 27730 34244 27786 34300
rect 27786 34244 27790 34300
rect 27726 34240 27790 34244
rect 27806 34300 27870 34304
rect 27806 34244 27810 34300
rect 27810 34244 27866 34300
rect 27866 34244 27870 34300
rect 27806 34240 27870 34244
rect 27886 34300 27950 34304
rect 27886 34244 27890 34300
rect 27890 34244 27946 34300
rect 27946 34244 27950 34300
rect 27886 34240 27950 34244
rect 18460 34096 18524 34100
rect 18460 34040 18510 34096
rect 18510 34040 18524 34096
rect 18460 34036 18524 34040
rect 3664 33756 3728 33760
rect 3664 33700 3668 33756
rect 3668 33700 3724 33756
rect 3724 33700 3728 33756
rect 3664 33696 3728 33700
rect 3744 33756 3808 33760
rect 3744 33700 3748 33756
rect 3748 33700 3804 33756
rect 3804 33700 3808 33756
rect 3744 33696 3808 33700
rect 3824 33756 3888 33760
rect 3824 33700 3828 33756
rect 3828 33700 3884 33756
rect 3884 33700 3888 33756
rect 3824 33696 3888 33700
rect 3904 33756 3968 33760
rect 3904 33700 3908 33756
rect 3908 33700 3964 33756
rect 3964 33700 3968 33756
rect 3904 33696 3968 33700
rect 11438 33756 11502 33760
rect 11438 33700 11442 33756
rect 11442 33700 11498 33756
rect 11498 33700 11502 33756
rect 11438 33696 11502 33700
rect 11518 33756 11582 33760
rect 11518 33700 11522 33756
rect 11522 33700 11578 33756
rect 11578 33700 11582 33756
rect 11518 33696 11582 33700
rect 11598 33756 11662 33760
rect 11598 33700 11602 33756
rect 11602 33700 11658 33756
rect 11658 33700 11662 33756
rect 11598 33696 11662 33700
rect 11678 33756 11742 33760
rect 11678 33700 11682 33756
rect 11682 33700 11738 33756
rect 11738 33700 11742 33756
rect 11678 33696 11742 33700
rect 19212 33756 19276 33760
rect 19212 33700 19216 33756
rect 19216 33700 19272 33756
rect 19272 33700 19276 33756
rect 19212 33696 19276 33700
rect 19292 33756 19356 33760
rect 19292 33700 19296 33756
rect 19296 33700 19352 33756
rect 19352 33700 19356 33756
rect 19292 33696 19356 33700
rect 19372 33756 19436 33760
rect 19372 33700 19376 33756
rect 19376 33700 19432 33756
rect 19432 33700 19436 33756
rect 19372 33696 19436 33700
rect 19452 33756 19516 33760
rect 19452 33700 19456 33756
rect 19456 33700 19512 33756
rect 19512 33700 19516 33756
rect 19452 33696 19516 33700
rect 26986 33756 27050 33760
rect 26986 33700 26990 33756
rect 26990 33700 27046 33756
rect 27046 33700 27050 33756
rect 26986 33696 27050 33700
rect 27066 33756 27130 33760
rect 27066 33700 27070 33756
rect 27070 33700 27126 33756
rect 27126 33700 27130 33756
rect 27066 33696 27130 33700
rect 27146 33756 27210 33760
rect 27146 33700 27150 33756
rect 27150 33700 27206 33756
rect 27206 33700 27210 33756
rect 27146 33696 27210 33700
rect 27226 33756 27290 33760
rect 27226 33700 27230 33756
rect 27230 33700 27286 33756
rect 27286 33700 27290 33756
rect 27226 33696 27290 33700
rect 4324 33212 4388 33216
rect 4324 33156 4328 33212
rect 4328 33156 4384 33212
rect 4384 33156 4388 33212
rect 4324 33152 4388 33156
rect 4404 33212 4468 33216
rect 4404 33156 4408 33212
rect 4408 33156 4464 33212
rect 4464 33156 4468 33212
rect 4404 33152 4468 33156
rect 4484 33212 4548 33216
rect 4484 33156 4488 33212
rect 4488 33156 4544 33212
rect 4544 33156 4548 33212
rect 4484 33152 4548 33156
rect 4564 33212 4628 33216
rect 4564 33156 4568 33212
rect 4568 33156 4624 33212
rect 4624 33156 4628 33212
rect 4564 33152 4628 33156
rect 12098 33212 12162 33216
rect 12098 33156 12102 33212
rect 12102 33156 12158 33212
rect 12158 33156 12162 33212
rect 12098 33152 12162 33156
rect 12178 33212 12242 33216
rect 12178 33156 12182 33212
rect 12182 33156 12238 33212
rect 12238 33156 12242 33212
rect 12178 33152 12242 33156
rect 12258 33212 12322 33216
rect 12258 33156 12262 33212
rect 12262 33156 12318 33212
rect 12318 33156 12322 33212
rect 12258 33152 12322 33156
rect 12338 33212 12402 33216
rect 12338 33156 12342 33212
rect 12342 33156 12398 33212
rect 12398 33156 12402 33212
rect 12338 33152 12402 33156
rect 19872 33212 19936 33216
rect 19872 33156 19876 33212
rect 19876 33156 19932 33212
rect 19932 33156 19936 33212
rect 19872 33152 19936 33156
rect 19952 33212 20016 33216
rect 19952 33156 19956 33212
rect 19956 33156 20012 33212
rect 20012 33156 20016 33212
rect 19952 33152 20016 33156
rect 20032 33212 20096 33216
rect 20032 33156 20036 33212
rect 20036 33156 20092 33212
rect 20092 33156 20096 33212
rect 20032 33152 20096 33156
rect 20112 33212 20176 33216
rect 20112 33156 20116 33212
rect 20116 33156 20172 33212
rect 20172 33156 20176 33212
rect 20112 33152 20176 33156
rect 27646 33212 27710 33216
rect 27646 33156 27650 33212
rect 27650 33156 27706 33212
rect 27706 33156 27710 33212
rect 27646 33152 27710 33156
rect 27726 33212 27790 33216
rect 27726 33156 27730 33212
rect 27730 33156 27786 33212
rect 27786 33156 27790 33212
rect 27726 33152 27790 33156
rect 27806 33212 27870 33216
rect 27806 33156 27810 33212
rect 27810 33156 27866 33212
rect 27866 33156 27870 33212
rect 27806 33152 27870 33156
rect 27886 33212 27950 33216
rect 27886 33156 27890 33212
rect 27890 33156 27946 33212
rect 27946 33156 27950 33212
rect 27886 33152 27950 33156
rect 3664 32668 3728 32672
rect 3664 32612 3668 32668
rect 3668 32612 3724 32668
rect 3724 32612 3728 32668
rect 3664 32608 3728 32612
rect 3744 32668 3808 32672
rect 3744 32612 3748 32668
rect 3748 32612 3804 32668
rect 3804 32612 3808 32668
rect 3744 32608 3808 32612
rect 3824 32668 3888 32672
rect 3824 32612 3828 32668
rect 3828 32612 3884 32668
rect 3884 32612 3888 32668
rect 3824 32608 3888 32612
rect 3904 32668 3968 32672
rect 3904 32612 3908 32668
rect 3908 32612 3964 32668
rect 3964 32612 3968 32668
rect 3904 32608 3968 32612
rect 11438 32668 11502 32672
rect 11438 32612 11442 32668
rect 11442 32612 11498 32668
rect 11498 32612 11502 32668
rect 11438 32608 11502 32612
rect 11518 32668 11582 32672
rect 11518 32612 11522 32668
rect 11522 32612 11578 32668
rect 11578 32612 11582 32668
rect 11518 32608 11582 32612
rect 11598 32668 11662 32672
rect 11598 32612 11602 32668
rect 11602 32612 11658 32668
rect 11658 32612 11662 32668
rect 11598 32608 11662 32612
rect 11678 32668 11742 32672
rect 11678 32612 11682 32668
rect 11682 32612 11738 32668
rect 11738 32612 11742 32668
rect 11678 32608 11742 32612
rect 19212 32668 19276 32672
rect 19212 32612 19216 32668
rect 19216 32612 19272 32668
rect 19272 32612 19276 32668
rect 19212 32608 19276 32612
rect 19292 32668 19356 32672
rect 19292 32612 19296 32668
rect 19296 32612 19352 32668
rect 19352 32612 19356 32668
rect 19292 32608 19356 32612
rect 19372 32668 19436 32672
rect 19372 32612 19376 32668
rect 19376 32612 19432 32668
rect 19432 32612 19436 32668
rect 19372 32608 19436 32612
rect 19452 32668 19516 32672
rect 19452 32612 19456 32668
rect 19456 32612 19512 32668
rect 19512 32612 19516 32668
rect 19452 32608 19516 32612
rect 26986 32668 27050 32672
rect 26986 32612 26990 32668
rect 26990 32612 27046 32668
rect 27046 32612 27050 32668
rect 26986 32608 27050 32612
rect 27066 32668 27130 32672
rect 27066 32612 27070 32668
rect 27070 32612 27126 32668
rect 27126 32612 27130 32668
rect 27066 32608 27130 32612
rect 27146 32668 27210 32672
rect 27146 32612 27150 32668
rect 27150 32612 27206 32668
rect 27206 32612 27210 32668
rect 27146 32608 27210 32612
rect 27226 32668 27290 32672
rect 27226 32612 27230 32668
rect 27230 32612 27286 32668
rect 27286 32612 27290 32668
rect 27226 32608 27290 32612
rect 4324 32124 4388 32128
rect 4324 32068 4328 32124
rect 4328 32068 4384 32124
rect 4384 32068 4388 32124
rect 4324 32064 4388 32068
rect 4404 32124 4468 32128
rect 4404 32068 4408 32124
rect 4408 32068 4464 32124
rect 4464 32068 4468 32124
rect 4404 32064 4468 32068
rect 4484 32124 4548 32128
rect 4484 32068 4488 32124
rect 4488 32068 4544 32124
rect 4544 32068 4548 32124
rect 4484 32064 4548 32068
rect 4564 32124 4628 32128
rect 4564 32068 4568 32124
rect 4568 32068 4624 32124
rect 4624 32068 4628 32124
rect 4564 32064 4628 32068
rect 12098 32124 12162 32128
rect 12098 32068 12102 32124
rect 12102 32068 12158 32124
rect 12158 32068 12162 32124
rect 12098 32064 12162 32068
rect 12178 32124 12242 32128
rect 12178 32068 12182 32124
rect 12182 32068 12238 32124
rect 12238 32068 12242 32124
rect 12178 32064 12242 32068
rect 12258 32124 12322 32128
rect 12258 32068 12262 32124
rect 12262 32068 12318 32124
rect 12318 32068 12322 32124
rect 12258 32064 12322 32068
rect 12338 32124 12402 32128
rect 12338 32068 12342 32124
rect 12342 32068 12398 32124
rect 12398 32068 12402 32124
rect 12338 32064 12402 32068
rect 19872 32124 19936 32128
rect 19872 32068 19876 32124
rect 19876 32068 19932 32124
rect 19932 32068 19936 32124
rect 19872 32064 19936 32068
rect 19952 32124 20016 32128
rect 19952 32068 19956 32124
rect 19956 32068 20012 32124
rect 20012 32068 20016 32124
rect 19952 32064 20016 32068
rect 20032 32124 20096 32128
rect 20032 32068 20036 32124
rect 20036 32068 20092 32124
rect 20092 32068 20096 32124
rect 20032 32064 20096 32068
rect 20112 32124 20176 32128
rect 20112 32068 20116 32124
rect 20116 32068 20172 32124
rect 20172 32068 20176 32124
rect 20112 32064 20176 32068
rect 27646 32124 27710 32128
rect 27646 32068 27650 32124
rect 27650 32068 27706 32124
rect 27706 32068 27710 32124
rect 27646 32064 27710 32068
rect 27726 32124 27790 32128
rect 27726 32068 27730 32124
rect 27730 32068 27786 32124
rect 27786 32068 27790 32124
rect 27726 32064 27790 32068
rect 27806 32124 27870 32128
rect 27806 32068 27810 32124
rect 27810 32068 27866 32124
rect 27866 32068 27870 32124
rect 27806 32064 27870 32068
rect 27886 32124 27950 32128
rect 27886 32068 27890 32124
rect 27890 32068 27946 32124
rect 27946 32068 27950 32124
rect 27886 32064 27950 32068
rect 16988 31860 17052 31924
rect 20300 31920 20364 31924
rect 20300 31864 20350 31920
rect 20350 31864 20364 31920
rect 20300 31860 20364 31864
rect 20300 31648 20364 31652
rect 20300 31592 20350 31648
rect 20350 31592 20364 31648
rect 20300 31588 20364 31592
rect 3664 31580 3728 31584
rect 3664 31524 3668 31580
rect 3668 31524 3724 31580
rect 3724 31524 3728 31580
rect 3664 31520 3728 31524
rect 3744 31580 3808 31584
rect 3744 31524 3748 31580
rect 3748 31524 3804 31580
rect 3804 31524 3808 31580
rect 3744 31520 3808 31524
rect 3824 31580 3888 31584
rect 3824 31524 3828 31580
rect 3828 31524 3884 31580
rect 3884 31524 3888 31580
rect 3824 31520 3888 31524
rect 3904 31580 3968 31584
rect 3904 31524 3908 31580
rect 3908 31524 3964 31580
rect 3964 31524 3968 31580
rect 3904 31520 3968 31524
rect 11438 31580 11502 31584
rect 11438 31524 11442 31580
rect 11442 31524 11498 31580
rect 11498 31524 11502 31580
rect 11438 31520 11502 31524
rect 11518 31580 11582 31584
rect 11518 31524 11522 31580
rect 11522 31524 11578 31580
rect 11578 31524 11582 31580
rect 11518 31520 11582 31524
rect 11598 31580 11662 31584
rect 11598 31524 11602 31580
rect 11602 31524 11658 31580
rect 11658 31524 11662 31580
rect 11598 31520 11662 31524
rect 11678 31580 11742 31584
rect 11678 31524 11682 31580
rect 11682 31524 11738 31580
rect 11738 31524 11742 31580
rect 11678 31520 11742 31524
rect 19212 31580 19276 31584
rect 19212 31524 19216 31580
rect 19216 31524 19272 31580
rect 19272 31524 19276 31580
rect 19212 31520 19276 31524
rect 19292 31580 19356 31584
rect 19292 31524 19296 31580
rect 19296 31524 19352 31580
rect 19352 31524 19356 31580
rect 19292 31520 19356 31524
rect 19372 31580 19436 31584
rect 19372 31524 19376 31580
rect 19376 31524 19432 31580
rect 19432 31524 19436 31580
rect 19372 31520 19436 31524
rect 19452 31580 19516 31584
rect 19452 31524 19456 31580
rect 19456 31524 19512 31580
rect 19512 31524 19516 31580
rect 19452 31520 19516 31524
rect 26986 31580 27050 31584
rect 26986 31524 26990 31580
rect 26990 31524 27046 31580
rect 27046 31524 27050 31580
rect 26986 31520 27050 31524
rect 27066 31580 27130 31584
rect 27066 31524 27070 31580
rect 27070 31524 27126 31580
rect 27126 31524 27130 31580
rect 27066 31520 27130 31524
rect 27146 31580 27210 31584
rect 27146 31524 27150 31580
rect 27150 31524 27206 31580
rect 27206 31524 27210 31580
rect 27146 31520 27210 31524
rect 27226 31580 27290 31584
rect 27226 31524 27230 31580
rect 27230 31524 27286 31580
rect 27286 31524 27290 31580
rect 27226 31520 27290 31524
rect 4324 31036 4388 31040
rect 4324 30980 4328 31036
rect 4328 30980 4384 31036
rect 4384 30980 4388 31036
rect 4324 30976 4388 30980
rect 4404 31036 4468 31040
rect 4404 30980 4408 31036
rect 4408 30980 4464 31036
rect 4464 30980 4468 31036
rect 4404 30976 4468 30980
rect 4484 31036 4548 31040
rect 4484 30980 4488 31036
rect 4488 30980 4544 31036
rect 4544 30980 4548 31036
rect 4484 30976 4548 30980
rect 4564 31036 4628 31040
rect 4564 30980 4568 31036
rect 4568 30980 4624 31036
rect 4624 30980 4628 31036
rect 4564 30976 4628 30980
rect 12098 31036 12162 31040
rect 12098 30980 12102 31036
rect 12102 30980 12158 31036
rect 12158 30980 12162 31036
rect 12098 30976 12162 30980
rect 12178 31036 12242 31040
rect 12178 30980 12182 31036
rect 12182 30980 12238 31036
rect 12238 30980 12242 31036
rect 12178 30976 12242 30980
rect 12258 31036 12322 31040
rect 12258 30980 12262 31036
rect 12262 30980 12318 31036
rect 12318 30980 12322 31036
rect 12258 30976 12322 30980
rect 12338 31036 12402 31040
rect 12338 30980 12342 31036
rect 12342 30980 12398 31036
rect 12398 30980 12402 31036
rect 12338 30976 12402 30980
rect 19872 31036 19936 31040
rect 19872 30980 19876 31036
rect 19876 30980 19932 31036
rect 19932 30980 19936 31036
rect 19872 30976 19936 30980
rect 19952 31036 20016 31040
rect 19952 30980 19956 31036
rect 19956 30980 20012 31036
rect 20012 30980 20016 31036
rect 19952 30976 20016 30980
rect 20032 31036 20096 31040
rect 20032 30980 20036 31036
rect 20036 30980 20092 31036
rect 20092 30980 20096 31036
rect 20032 30976 20096 30980
rect 20112 31036 20176 31040
rect 20112 30980 20116 31036
rect 20116 30980 20172 31036
rect 20172 30980 20176 31036
rect 20112 30976 20176 30980
rect 27646 31036 27710 31040
rect 27646 30980 27650 31036
rect 27650 30980 27706 31036
rect 27706 30980 27710 31036
rect 27646 30976 27710 30980
rect 27726 31036 27790 31040
rect 27726 30980 27730 31036
rect 27730 30980 27786 31036
rect 27786 30980 27790 31036
rect 27726 30976 27790 30980
rect 27806 31036 27870 31040
rect 27806 30980 27810 31036
rect 27810 30980 27866 31036
rect 27866 30980 27870 31036
rect 27806 30976 27870 30980
rect 27886 31036 27950 31040
rect 27886 30980 27890 31036
rect 27890 30980 27946 31036
rect 27946 30980 27950 31036
rect 27886 30976 27950 30980
rect 26740 30696 26804 30700
rect 26740 30640 26754 30696
rect 26754 30640 26804 30696
rect 26740 30636 26804 30640
rect 3664 30492 3728 30496
rect 3664 30436 3668 30492
rect 3668 30436 3724 30492
rect 3724 30436 3728 30492
rect 3664 30432 3728 30436
rect 3744 30492 3808 30496
rect 3744 30436 3748 30492
rect 3748 30436 3804 30492
rect 3804 30436 3808 30492
rect 3744 30432 3808 30436
rect 3824 30492 3888 30496
rect 3824 30436 3828 30492
rect 3828 30436 3884 30492
rect 3884 30436 3888 30492
rect 3824 30432 3888 30436
rect 3904 30492 3968 30496
rect 3904 30436 3908 30492
rect 3908 30436 3964 30492
rect 3964 30436 3968 30492
rect 3904 30432 3968 30436
rect 11438 30492 11502 30496
rect 11438 30436 11442 30492
rect 11442 30436 11498 30492
rect 11498 30436 11502 30492
rect 11438 30432 11502 30436
rect 11518 30492 11582 30496
rect 11518 30436 11522 30492
rect 11522 30436 11578 30492
rect 11578 30436 11582 30492
rect 11518 30432 11582 30436
rect 11598 30492 11662 30496
rect 11598 30436 11602 30492
rect 11602 30436 11658 30492
rect 11658 30436 11662 30492
rect 11598 30432 11662 30436
rect 11678 30492 11742 30496
rect 11678 30436 11682 30492
rect 11682 30436 11738 30492
rect 11738 30436 11742 30492
rect 11678 30432 11742 30436
rect 19212 30492 19276 30496
rect 19212 30436 19216 30492
rect 19216 30436 19272 30492
rect 19272 30436 19276 30492
rect 19212 30432 19276 30436
rect 19292 30492 19356 30496
rect 19292 30436 19296 30492
rect 19296 30436 19352 30492
rect 19352 30436 19356 30492
rect 19292 30432 19356 30436
rect 19372 30492 19436 30496
rect 19372 30436 19376 30492
rect 19376 30436 19432 30492
rect 19432 30436 19436 30492
rect 19372 30432 19436 30436
rect 19452 30492 19516 30496
rect 19452 30436 19456 30492
rect 19456 30436 19512 30492
rect 19512 30436 19516 30492
rect 19452 30432 19516 30436
rect 26986 30492 27050 30496
rect 26986 30436 26990 30492
rect 26990 30436 27046 30492
rect 27046 30436 27050 30492
rect 26986 30432 27050 30436
rect 27066 30492 27130 30496
rect 27066 30436 27070 30492
rect 27070 30436 27126 30492
rect 27126 30436 27130 30492
rect 27066 30432 27130 30436
rect 27146 30492 27210 30496
rect 27146 30436 27150 30492
rect 27150 30436 27206 30492
rect 27206 30436 27210 30492
rect 27146 30432 27210 30436
rect 27226 30492 27290 30496
rect 27226 30436 27230 30492
rect 27230 30436 27286 30492
rect 27286 30436 27290 30492
rect 27226 30432 27290 30436
rect 23612 30288 23676 30292
rect 23612 30232 23626 30288
rect 23626 30232 23676 30288
rect 23612 30228 23676 30232
rect 4324 29948 4388 29952
rect 4324 29892 4328 29948
rect 4328 29892 4384 29948
rect 4384 29892 4388 29948
rect 4324 29888 4388 29892
rect 4404 29948 4468 29952
rect 4404 29892 4408 29948
rect 4408 29892 4464 29948
rect 4464 29892 4468 29948
rect 4404 29888 4468 29892
rect 4484 29948 4548 29952
rect 4484 29892 4488 29948
rect 4488 29892 4544 29948
rect 4544 29892 4548 29948
rect 4484 29888 4548 29892
rect 4564 29948 4628 29952
rect 4564 29892 4568 29948
rect 4568 29892 4624 29948
rect 4624 29892 4628 29948
rect 4564 29888 4628 29892
rect 12098 29948 12162 29952
rect 12098 29892 12102 29948
rect 12102 29892 12158 29948
rect 12158 29892 12162 29948
rect 12098 29888 12162 29892
rect 12178 29948 12242 29952
rect 12178 29892 12182 29948
rect 12182 29892 12238 29948
rect 12238 29892 12242 29948
rect 12178 29888 12242 29892
rect 12258 29948 12322 29952
rect 12258 29892 12262 29948
rect 12262 29892 12318 29948
rect 12318 29892 12322 29948
rect 12258 29888 12322 29892
rect 12338 29948 12402 29952
rect 12338 29892 12342 29948
rect 12342 29892 12398 29948
rect 12398 29892 12402 29948
rect 12338 29888 12402 29892
rect 19872 29948 19936 29952
rect 19872 29892 19876 29948
rect 19876 29892 19932 29948
rect 19932 29892 19936 29948
rect 19872 29888 19936 29892
rect 19952 29948 20016 29952
rect 19952 29892 19956 29948
rect 19956 29892 20012 29948
rect 20012 29892 20016 29948
rect 19952 29888 20016 29892
rect 20032 29948 20096 29952
rect 20032 29892 20036 29948
rect 20036 29892 20092 29948
rect 20092 29892 20096 29948
rect 20032 29888 20096 29892
rect 20112 29948 20176 29952
rect 20112 29892 20116 29948
rect 20116 29892 20172 29948
rect 20172 29892 20176 29948
rect 20112 29888 20176 29892
rect 27646 29948 27710 29952
rect 27646 29892 27650 29948
rect 27650 29892 27706 29948
rect 27706 29892 27710 29948
rect 27646 29888 27710 29892
rect 27726 29948 27790 29952
rect 27726 29892 27730 29948
rect 27730 29892 27786 29948
rect 27786 29892 27790 29948
rect 27726 29888 27790 29892
rect 27806 29948 27870 29952
rect 27806 29892 27810 29948
rect 27810 29892 27866 29948
rect 27866 29892 27870 29948
rect 27806 29888 27870 29892
rect 27886 29948 27950 29952
rect 27886 29892 27890 29948
rect 27890 29892 27946 29948
rect 27946 29892 27950 29948
rect 27886 29888 27950 29892
rect 3664 29404 3728 29408
rect 3664 29348 3668 29404
rect 3668 29348 3724 29404
rect 3724 29348 3728 29404
rect 3664 29344 3728 29348
rect 3744 29404 3808 29408
rect 3744 29348 3748 29404
rect 3748 29348 3804 29404
rect 3804 29348 3808 29404
rect 3744 29344 3808 29348
rect 3824 29404 3888 29408
rect 3824 29348 3828 29404
rect 3828 29348 3884 29404
rect 3884 29348 3888 29404
rect 3824 29344 3888 29348
rect 3904 29404 3968 29408
rect 3904 29348 3908 29404
rect 3908 29348 3964 29404
rect 3964 29348 3968 29404
rect 3904 29344 3968 29348
rect 11438 29404 11502 29408
rect 11438 29348 11442 29404
rect 11442 29348 11498 29404
rect 11498 29348 11502 29404
rect 11438 29344 11502 29348
rect 11518 29404 11582 29408
rect 11518 29348 11522 29404
rect 11522 29348 11578 29404
rect 11578 29348 11582 29404
rect 11518 29344 11582 29348
rect 11598 29404 11662 29408
rect 11598 29348 11602 29404
rect 11602 29348 11658 29404
rect 11658 29348 11662 29404
rect 11598 29344 11662 29348
rect 11678 29404 11742 29408
rect 11678 29348 11682 29404
rect 11682 29348 11738 29404
rect 11738 29348 11742 29404
rect 11678 29344 11742 29348
rect 19212 29404 19276 29408
rect 19212 29348 19216 29404
rect 19216 29348 19272 29404
rect 19272 29348 19276 29404
rect 19212 29344 19276 29348
rect 19292 29404 19356 29408
rect 19292 29348 19296 29404
rect 19296 29348 19352 29404
rect 19352 29348 19356 29404
rect 19292 29344 19356 29348
rect 19372 29404 19436 29408
rect 19372 29348 19376 29404
rect 19376 29348 19432 29404
rect 19432 29348 19436 29404
rect 19372 29344 19436 29348
rect 19452 29404 19516 29408
rect 19452 29348 19456 29404
rect 19456 29348 19512 29404
rect 19512 29348 19516 29404
rect 19452 29344 19516 29348
rect 26986 29404 27050 29408
rect 26986 29348 26990 29404
rect 26990 29348 27046 29404
rect 27046 29348 27050 29404
rect 26986 29344 27050 29348
rect 27066 29404 27130 29408
rect 27066 29348 27070 29404
rect 27070 29348 27126 29404
rect 27126 29348 27130 29404
rect 27066 29344 27130 29348
rect 27146 29404 27210 29408
rect 27146 29348 27150 29404
rect 27150 29348 27206 29404
rect 27206 29348 27210 29404
rect 27146 29344 27210 29348
rect 27226 29404 27290 29408
rect 27226 29348 27230 29404
rect 27230 29348 27286 29404
rect 27286 29348 27290 29404
rect 27226 29344 27290 29348
rect 20668 29140 20732 29204
rect 4324 28860 4388 28864
rect 4324 28804 4328 28860
rect 4328 28804 4384 28860
rect 4384 28804 4388 28860
rect 4324 28800 4388 28804
rect 4404 28860 4468 28864
rect 4404 28804 4408 28860
rect 4408 28804 4464 28860
rect 4464 28804 4468 28860
rect 4404 28800 4468 28804
rect 4484 28860 4548 28864
rect 4484 28804 4488 28860
rect 4488 28804 4544 28860
rect 4544 28804 4548 28860
rect 4484 28800 4548 28804
rect 4564 28860 4628 28864
rect 4564 28804 4568 28860
rect 4568 28804 4624 28860
rect 4624 28804 4628 28860
rect 4564 28800 4628 28804
rect 12098 28860 12162 28864
rect 12098 28804 12102 28860
rect 12102 28804 12158 28860
rect 12158 28804 12162 28860
rect 12098 28800 12162 28804
rect 12178 28860 12242 28864
rect 12178 28804 12182 28860
rect 12182 28804 12238 28860
rect 12238 28804 12242 28860
rect 12178 28800 12242 28804
rect 12258 28860 12322 28864
rect 12258 28804 12262 28860
rect 12262 28804 12318 28860
rect 12318 28804 12322 28860
rect 12258 28800 12322 28804
rect 12338 28860 12402 28864
rect 12338 28804 12342 28860
rect 12342 28804 12398 28860
rect 12398 28804 12402 28860
rect 12338 28800 12402 28804
rect 19872 28860 19936 28864
rect 19872 28804 19876 28860
rect 19876 28804 19932 28860
rect 19932 28804 19936 28860
rect 19872 28800 19936 28804
rect 19952 28860 20016 28864
rect 19952 28804 19956 28860
rect 19956 28804 20012 28860
rect 20012 28804 20016 28860
rect 19952 28800 20016 28804
rect 20032 28860 20096 28864
rect 20032 28804 20036 28860
rect 20036 28804 20092 28860
rect 20092 28804 20096 28860
rect 20032 28800 20096 28804
rect 20112 28860 20176 28864
rect 20112 28804 20116 28860
rect 20116 28804 20172 28860
rect 20172 28804 20176 28860
rect 20112 28800 20176 28804
rect 27646 28860 27710 28864
rect 27646 28804 27650 28860
rect 27650 28804 27706 28860
rect 27706 28804 27710 28860
rect 27646 28800 27710 28804
rect 27726 28860 27790 28864
rect 27726 28804 27730 28860
rect 27730 28804 27786 28860
rect 27786 28804 27790 28860
rect 27726 28800 27790 28804
rect 27806 28860 27870 28864
rect 27806 28804 27810 28860
rect 27810 28804 27866 28860
rect 27866 28804 27870 28860
rect 27806 28800 27870 28804
rect 27886 28860 27950 28864
rect 27886 28804 27890 28860
rect 27890 28804 27946 28860
rect 27946 28804 27950 28860
rect 27886 28800 27950 28804
rect 13676 28732 13740 28796
rect 21956 28656 22020 28660
rect 21956 28600 21970 28656
rect 21970 28600 22020 28656
rect 21956 28596 22020 28600
rect 28764 28460 28828 28524
rect 3664 28316 3728 28320
rect 3664 28260 3668 28316
rect 3668 28260 3724 28316
rect 3724 28260 3728 28316
rect 3664 28256 3728 28260
rect 3744 28316 3808 28320
rect 3744 28260 3748 28316
rect 3748 28260 3804 28316
rect 3804 28260 3808 28316
rect 3744 28256 3808 28260
rect 3824 28316 3888 28320
rect 3824 28260 3828 28316
rect 3828 28260 3884 28316
rect 3884 28260 3888 28316
rect 3824 28256 3888 28260
rect 3904 28316 3968 28320
rect 3904 28260 3908 28316
rect 3908 28260 3964 28316
rect 3964 28260 3968 28316
rect 3904 28256 3968 28260
rect 11438 28316 11502 28320
rect 11438 28260 11442 28316
rect 11442 28260 11498 28316
rect 11498 28260 11502 28316
rect 11438 28256 11502 28260
rect 11518 28316 11582 28320
rect 11518 28260 11522 28316
rect 11522 28260 11578 28316
rect 11578 28260 11582 28316
rect 11518 28256 11582 28260
rect 11598 28316 11662 28320
rect 11598 28260 11602 28316
rect 11602 28260 11658 28316
rect 11658 28260 11662 28316
rect 11598 28256 11662 28260
rect 11678 28316 11742 28320
rect 11678 28260 11682 28316
rect 11682 28260 11738 28316
rect 11738 28260 11742 28316
rect 11678 28256 11742 28260
rect 19212 28316 19276 28320
rect 19212 28260 19216 28316
rect 19216 28260 19272 28316
rect 19272 28260 19276 28316
rect 19212 28256 19276 28260
rect 19292 28316 19356 28320
rect 19292 28260 19296 28316
rect 19296 28260 19352 28316
rect 19352 28260 19356 28316
rect 19292 28256 19356 28260
rect 19372 28316 19436 28320
rect 19372 28260 19376 28316
rect 19376 28260 19432 28316
rect 19432 28260 19436 28316
rect 19372 28256 19436 28260
rect 19452 28316 19516 28320
rect 19452 28260 19456 28316
rect 19456 28260 19512 28316
rect 19512 28260 19516 28316
rect 19452 28256 19516 28260
rect 26986 28316 27050 28320
rect 26986 28260 26990 28316
rect 26990 28260 27046 28316
rect 27046 28260 27050 28316
rect 26986 28256 27050 28260
rect 27066 28316 27130 28320
rect 27066 28260 27070 28316
rect 27070 28260 27126 28316
rect 27126 28260 27130 28316
rect 27066 28256 27130 28260
rect 27146 28316 27210 28320
rect 27146 28260 27150 28316
rect 27150 28260 27206 28316
rect 27206 28260 27210 28316
rect 27146 28256 27210 28260
rect 27226 28316 27290 28320
rect 27226 28260 27230 28316
rect 27230 28260 27286 28316
rect 27286 28260 27290 28316
rect 27226 28256 27290 28260
rect 24532 28112 24596 28116
rect 24532 28056 24546 28112
rect 24546 28056 24596 28112
rect 24532 28052 24596 28056
rect 4324 27772 4388 27776
rect 4324 27716 4328 27772
rect 4328 27716 4384 27772
rect 4384 27716 4388 27772
rect 4324 27712 4388 27716
rect 4404 27772 4468 27776
rect 4404 27716 4408 27772
rect 4408 27716 4464 27772
rect 4464 27716 4468 27772
rect 4404 27712 4468 27716
rect 4484 27772 4548 27776
rect 4484 27716 4488 27772
rect 4488 27716 4544 27772
rect 4544 27716 4548 27772
rect 4484 27712 4548 27716
rect 4564 27772 4628 27776
rect 4564 27716 4568 27772
rect 4568 27716 4624 27772
rect 4624 27716 4628 27772
rect 4564 27712 4628 27716
rect 12098 27772 12162 27776
rect 12098 27716 12102 27772
rect 12102 27716 12158 27772
rect 12158 27716 12162 27772
rect 12098 27712 12162 27716
rect 12178 27772 12242 27776
rect 12178 27716 12182 27772
rect 12182 27716 12238 27772
rect 12238 27716 12242 27772
rect 12178 27712 12242 27716
rect 12258 27772 12322 27776
rect 12258 27716 12262 27772
rect 12262 27716 12318 27772
rect 12318 27716 12322 27772
rect 12258 27712 12322 27716
rect 12338 27772 12402 27776
rect 12338 27716 12342 27772
rect 12342 27716 12398 27772
rect 12398 27716 12402 27772
rect 12338 27712 12402 27716
rect 19872 27772 19936 27776
rect 19872 27716 19876 27772
rect 19876 27716 19932 27772
rect 19932 27716 19936 27772
rect 19872 27712 19936 27716
rect 19952 27772 20016 27776
rect 19952 27716 19956 27772
rect 19956 27716 20012 27772
rect 20012 27716 20016 27772
rect 19952 27712 20016 27716
rect 20032 27772 20096 27776
rect 20032 27716 20036 27772
rect 20036 27716 20092 27772
rect 20092 27716 20096 27772
rect 20032 27712 20096 27716
rect 20112 27772 20176 27776
rect 20112 27716 20116 27772
rect 20116 27716 20172 27772
rect 20172 27716 20176 27772
rect 20112 27712 20176 27716
rect 27646 27772 27710 27776
rect 27646 27716 27650 27772
rect 27650 27716 27706 27772
rect 27706 27716 27710 27772
rect 27646 27712 27710 27716
rect 27726 27772 27790 27776
rect 27726 27716 27730 27772
rect 27730 27716 27786 27772
rect 27786 27716 27790 27772
rect 27726 27712 27790 27716
rect 27806 27772 27870 27776
rect 27806 27716 27810 27772
rect 27810 27716 27866 27772
rect 27866 27716 27870 27772
rect 27806 27712 27870 27716
rect 27886 27772 27950 27776
rect 27886 27716 27890 27772
rect 27890 27716 27946 27772
rect 27946 27716 27950 27772
rect 27886 27712 27950 27716
rect 3664 27228 3728 27232
rect 3664 27172 3668 27228
rect 3668 27172 3724 27228
rect 3724 27172 3728 27228
rect 3664 27168 3728 27172
rect 3744 27228 3808 27232
rect 3744 27172 3748 27228
rect 3748 27172 3804 27228
rect 3804 27172 3808 27228
rect 3744 27168 3808 27172
rect 3824 27228 3888 27232
rect 3824 27172 3828 27228
rect 3828 27172 3884 27228
rect 3884 27172 3888 27228
rect 3824 27168 3888 27172
rect 3904 27228 3968 27232
rect 3904 27172 3908 27228
rect 3908 27172 3964 27228
rect 3964 27172 3968 27228
rect 3904 27168 3968 27172
rect 11438 27228 11502 27232
rect 11438 27172 11442 27228
rect 11442 27172 11498 27228
rect 11498 27172 11502 27228
rect 11438 27168 11502 27172
rect 11518 27228 11582 27232
rect 11518 27172 11522 27228
rect 11522 27172 11578 27228
rect 11578 27172 11582 27228
rect 11518 27168 11582 27172
rect 11598 27228 11662 27232
rect 11598 27172 11602 27228
rect 11602 27172 11658 27228
rect 11658 27172 11662 27228
rect 11598 27168 11662 27172
rect 11678 27228 11742 27232
rect 11678 27172 11682 27228
rect 11682 27172 11738 27228
rect 11738 27172 11742 27228
rect 11678 27168 11742 27172
rect 19212 27228 19276 27232
rect 19212 27172 19216 27228
rect 19216 27172 19272 27228
rect 19272 27172 19276 27228
rect 19212 27168 19276 27172
rect 19292 27228 19356 27232
rect 19292 27172 19296 27228
rect 19296 27172 19352 27228
rect 19352 27172 19356 27228
rect 19292 27168 19356 27172
rect 19372 27228 19436 27232
rect 19372 27172 19376 27228
rect 19376 27172 19432 27228
rect 19432 27172 19436 27228
rect 19372 27168 19436 27172
rect 19452 27228 19516 27232
rect 19452 27172 19456 27228
rect 19456 27172 19512 27228
rect 19512 27172 19516 27228
rect 19452 27168 19516 27172
rect 26986 27228 27050 27232
rect 26986 27172 26990 27228
rect 26990 27172 27046 27228
rect 27046 27172 27050 27228
rect 26986 27168 27050 27172
rect 27066 27228 27130 27232
rect 27066 27172 27070 27228
rect 27070 27172 27126 27228
rect 27126 27172 27130 27228
rect 27066 27168 27130 27172
rect 27146 27228 27210 27232
rect 27146 27172 27150 27228
rect 27150 27172 27206 27228
rect 27206 27172 27210 27228
rect 27146 27168 27210 27172
rect 27226 27228 27290 27232
rect 27226 27172 27230 27228
rect 27230 27172 27286 27228
rect 27286 27172 27290 27228
rect 27226 27168 27290 27172
rect 4324 26684 4388 26688
rect 4324 26628 4328 26684
rect 4328 26628 4384 26684
rect 4384 26628 4388 26684
rect 4324 26624 4388 26628
rect 4404 26684 4468 26688
rect 4404 26628 4408 26684
rect 4408 26628 4464 26684
rect 4464 26628 4468 26684
rect 4404 26624 4468 26628
rect 4484 26684 4548 26688
rect 4484 26628 4488 26684
rect 4488 26628 4544 26684
rect 4544 26628 4548 26684
rect 4484 26624 4548 26628
rect 4564 26684 4628 26688
rect 4564 26628 4568 26684
rect 4568 26628 4624 26684
rect 4624 26628 4628 26684
rect 4564 26624 4628 26628
rect 12098 26684 12162 26688
rect 12098 26628 12102 26684
rect 12102 26628 12158 26684
rect 12158 26628 12162 26684
rect 12098 26624 12162 26628
rect 12178 26684 12242 26688
rect 12178 26628 12182 26684
rect 12182 26628 12238 26684
rect 12238 26628 12242 26684
rect 12178 26624 12242 26628
rect 12258 26684 12322 26688
rect 12258 26628 12262 26684
rect 12262 26628 12318 26684
rect 12318 26628 12322 26684
rect 12258 26624 12322 26628
rect 12338 26684 12402 26688
rect 12338 26628 12342 26684
rect 12342 26628 12398 26684
rect 12398 26628 12402 26684
rect 12338 26624 12402 26628
rect 19872 26684 19936 26688
rect 19872 26628 19876 26684
rect 19876 26628 19932 26684
rect 19932 26628 19936 26684
rect 19872 26624 19936 26628
rect 19952 26684 20016 26688
rect 19952 26628 19956 26684
rect 19956 26628 20012 26684
rect 20012 26628 20016 26684
rect 19952 26624 20016 26628
rect 20032 26684 20096 26688
rect 20032 26628 20036 26684
rect 20036 26628 20092 26684
rect 20092 26628 20096 26684
rect 20032 26624 20096 26628
rect 20112 26684 20176 26688
rect 20112 26628 20116 26684
rect 20116 26628 20172 26684
rect 20172 26628 20176 26684
rect 20112 26624 20176 26628
rect 27646 26684 27710 26688
rect 27646 26628 27650 26684
rect 27650 26628 27706 26684
rect 27706 26628 27710 26684
rect 27646 26624 27710 26628
rect 27726 26684 27790 26688
rect 27726 26628 27730 26684
rect 27730 26628 27786 26684
rect 27786 26628 27790 26684
rect 27726 26624 27790 26628
rect 27806 26684 27870 26688
rect 27806 26628 27810 26684
rect 27810 26628 27866 26684
rect 27866 26628 27870 26684
rect 27806 26624 27870 26628
rect 27886 26684 27950 26688
rect 27886 26628 27890 26684
rect 27890 26628 27946 26684
rect 27946 26628 27950 26684
rect 27886 26624 27950 26628
rect 3664 26140 3728 26144
rect 3664 26084 3668 26140
rect 3668 26084 3724 26140
rect 3724 26084 3728 26140
rect 3664 26080 3728 26084
rect 3744 26140 3808 26144
rect 3744 26084 3748 26140
rect 3748 26084 3804 26140
rect 3804 26084 3808 26140
rect 3744 26080 3808 26084
rect 3824 26140 3888 26144
rect 3824 26084 3828 26140
rect 3828 26084 3884 26140
rect 3884 26084 3888 26140
rect 3824 26080 3888 26084
rect 3904 26140 3968 26144
rect 3904 26084 3908 26140
rect 3908 26084 3964 26140
rect 3964 26084 3968 26140
rect 3904 26080 3968 26084
rect 11438 26140 11502 26144
rect 11438 26084 11442 26140
rect 11442 26084 11498 26140
rect 11498 26084 11502 26140
rect 11438 26080 11502 26084
rect 11518 26140 11582 26144
rect 11518 26084 11522 26140
rect 11522 26084 11578 26140
rect 11578 26084 11582 26140
rect 11518 26080 11582 26084
rect 11598 26140 11662 26144
rect 11598 26084 11602 26140
rect 11602 26084 11658 26140
rect 11658 26084 11662 26140
rect 11598 26080 11662 26084
rect 11678 26140 11742 26144
rect 11678 26084 11682 26140
rect 11682 26084 11738 26140
rect 11738 26084 11742 26140
rect 11678 26080 11742 26084
rect 19212 26140 19276 26144
rect 19212 26084 19216 26140
rect 19216 26084 19272 26140
rect 19272 26084 19276 26140
rect 19212 26080 19276 26084
rect 19292 26140 19356 26144
rect 19292 26084 19296 26140
rect 19296 26084 19352 26140
rect 19352 26084 19356 26140
rect 19292 26080 19356 26084
rect 19372 26140 19436 26144
rect 19372 26084 19376 26140
rect 19376 26084 19432 26140
rect 19432 26084 19436 26140
rect 19372 26080 19436 26084
rect 19452 26140 19516 26144
rect 19452 26084 19456 26140
rect 19456 26084 19512 26140
rect 19512 26084 19516 26140
rect 19452 26080 19516 26084
rect 26986 26140 27050 26144
rect 26986 26084 26990 26140
rect 26990 26084 27046 26140
rect 27046 26084 27050 26140
rect 26986 26080 27050 26084
rect 27066 26140 27130 26144
rect 27066 26084 27070 26140
rect 27070 26084 27126 26140
rect 27126 26084 27130 26140
rect 27066 26080 27130 26084
rect 27146 26140 27210 26144
rect 27146 26084 27150 26140
rect 27150 26084 27206 26140
rect 27206 26084 27210 26140
rect 27146 26080 27210 26084
rect 27226 26140 27290 26144
rect 27226 26084 27230 26140
rect 27230 26084 27286 26140
rect 27286 26084 27290 26140
rect 27226 26080 27290 26084
rect 4324 25596 4388 25600
rect 4324 25540 4328 25596
rect 4328 25540 4384 25596
rect 4384 25540 4388 25596
rect 4324 25536 4388 25540
rect 4404 25596 4468 25600
rect 4404 25540 4408 25596
rect 4408 25540 4464 25596
rect 4464 25540 4468 25596
rect 4404 25536 4468 25540
rect 4484 25596 4548 25600
rect 4484 25540 4488 25596
rect 4488 25540 4544 25596
rect 4544 25540 4548 25596
rect 4484 25536 4548 25540
rect 4564 25596 4628 25600
rect 4564 25540 4568 25596
rect 4568 25540 4624 25596
rect 4624 25540 4628 25596
rect 4564 25536 4628 25540
rect 12098 25596 12162 25600
rect 12098 25540 12102 25596
rect 12102 25540 12158 25596
rect 12158 25540 12162 25596
rect 12098 25536 12162 25540
rect 12178 25596 12242 25600
rect 12178 25540 12182 25596
rect 12182 25540 12238 25596
rect 12238 25540 12242 25596
rect 12178 25536 12242 25540
rect 12258 25596 12322 25600
rect 12258 25540 12262 25596
rect 12262 25540 12318 25596
rect 12318 25540 12322 25596
rect 12258 25536 12322 25540
rect 12338 25596 12402 25600
rect 12338 25540 12342 25596
rect 12342 25540 12398 25596
rect 12398 25540 12402 25596
rect 12338 25536 12402 25540
rect 19872 25596 19936 25600
rect 19872 25540 19876 25596
rect 19876 25540 19932 25596
rect 19932 25540 19936 25596
rect 19872 25536 19936 25540
rect 19952 25596 20016 25600
rect 19952 25540 19956 25596
rect 19956 25540 20012 25596
rect 20012 25540 20016 25596
rect 19952 25536 20016 25540
rect 20032 25596 20096 25600
rect 20032 25540 20036 25596
rect 20036 25540 20092 25596
rect 20092 25540 20096 25596
rect 20032 25536 20096 25540
rect 20112 25596 20176 25600
rect 20112 25540 20116 25596
rect 20116 25540 20172 25596
rect 20172 25540 20176 25596
rect 20112 25536 20176 25540
rect 27646 25596 27710 25600
rect 27646 25540 27650 25596
rect 27650 25540 27706 25596
rect 27706 25540 27710 25596
rect 27646 25536 27710 25540
rect 27726 25596 27790 25600
rect 27726 25540 27730 25596
rect 27730 25540 27786 25596
rect 27786 25540 27790 25596
rect 27726 25536 27790 25540
rect 27806 25596 27870 25600
rect 27806 25540 27810 25596
rect 27810 25540 27866 25596
rect 27866 25540 27870 25596
rect 27806 25536 27870 25540
rect 27886 25596 27950 25600
rect 27886 25540 27890 25596
rect 27890 25540 27946 25596
rect 27946 25540 27950 25596
rect 27886 25536 27950 25540
rect 3664 25052 3728 25056
rect 3664 24996 3668 25052
rect 3668 24996 3724 25052
rect 3724 24996 3728 25052
rect 3664 24992 3728 24996
rect 3744 25052 3808 25056
rect 3744 24996 3748 25052
rect 3748 24996 3804 25052
rect 3804 24996 3808 25052
rect 3744 24992 3808 24996
rect 3824 25052 3888 25056
rect 3824 24996 3828 25052
rect 3828 24996 3884 25052
rect 3884 24996 3888 25052
rect 3824 24992 3888 24996
rect 3904 25052 3968 25056
rect 3904 24996 3908 25052
rect 3908 24996 3964 25052
rect 3964 24996 3968 25052
rect 3904 24992 3968 24996
rect 11438 25052 11502 25056
rect 11438 24996 11442 25052
rect 11442 24996 11498 25052
rect 11498 24996 11502 25052
rect 11438 24992 11502 24996
rect 11518 25052 11582 25056
rect 11518 24996 11522 25052
rect 11522 24996 11578 25052
rect 11578 24996 11582 25052
rect 11518 24992 11582 24996
rect 11598 25052 11662 25056
rect 11598 24996 11602 25052
rect 11602 24996 11658 25052
rect 11658 24996 11662 25052
rect 11598 24992 11662 24996
rect 11678 25052 11742 25056
rect 11678 24996 11682 25052
rect 11682 24996 11738 25052
rect 11738 24996 11742 25052
rect 11678 24992 11742 24996
rect 19212 25052 19276 25056
rect 19212 24996 19216 25052
rect 19216 24996 19272 25052
rect 19272 24996 19276 25052
rect 19212 24992 19276 24996
rect 19292 25052 19356 25056
rect 19292 24996 19296 25052
rect 19296 24996 19352 25052
rect 19352 24996 19356 25052
rect 19292 24992 19356 24996
rect 19372 25052 19436 25056
rect 19372 24996 19376 25052
rect 19376 24996 19432 25052
rect 19432 24996 19436 25052
rect 19372 24992 19436 24996
rect 19452 25052 19516 25056
rect 19452 24996 19456 25052
rect 19456 24996 19512 25052
rect 19512 24996 19516 25052
rect 19452 24992 19516 24996
rect 26986 25052 27050 25056
rect 26986 24996 26990 25052
rect 26990 24996 27046 25052
rect 27046 24996 27050 25052
rect 26986 24992 27050 24996
rect 27066 25052 27130 25056
rect 27066 24996 27070 25052
rect 27070 24996 27126 25052
rect 27126 24996 27130 25052
rect 27066 24992 27130 24996
rect 27146 25052 27210 25056
rect 27146 24996 27150 25052
rect 27150 24996 27206 25052
rect 27206 24996 27210 25052
rect 27146 24992 27210 24996
rect 27226 25052 27290 25056
rect 27226 24996 27230 25052
rect 27230 24996 27286 25052
rect 27286 24996 27290 25052
rect 27226 24992 27290 24996
rect 4324 24508 4388 24512
rect 4324 24452 4328 24508
rect 4328 24452 4384 24508
rect 4384 24452 4388 24508
rect 4324 24448 4388 24452
rect 4404 24508 4468 24512
rect 4404 24452 4408 24508
rect 4408 24452 4464 24508
rect 4464 24452 4468 24508
rect 4404 24448 4468 24452
rect 4484 24508 4548 24512
rect 4484 24452 4488 24508
rect 4488 24452 4544 24508
rect 4544 24452 4548 24508
rect 4484 24448 4548 24452
rect 4564 24508 4628 24512
rect 4564 24452 4568 24508
rect 4568 24452 4624 24508
rect 4624 24452 4628 24508
rect 4564 24448 4628 24452
rect 12098 24508 12162 24512
rect 12098 24452 12102 24508
rect 12102 24452 12158 24508
rect 12158 24452 12162 24508
rect 12098 24448 12162 24452
rect 12178 24508 12242 24512
rect 12178 24452 12182 24508
rect 12182 24452 12238 24508
rect 12238 24452 12242 24508
rect 12178 24448 12242 24452
rect 12258 24508 12322 24512
rect 12258 24452 12262 24508
rect 12262 24452 12318 24508
rect 12318 24452 12322 24508
rect 12258 24448 12322 24452
rect 12338 24508 12402 24512
rect 12338 24452 12342 24508
rect 12342 24452 12398 24508
rect 12398 24452 12402 24508
rect 12338 24448 12402 24452
rect 19872 24508 19936 24512
rect 19872 24452 19876 24508
rect 19876 24452 19932 24508
rect 19932 24452 19936 24508
rect 19872 24448 19936 24452
rect 19952 24508 20016 24512
rect 19952 24452 19956 24508
rect 19956 24452 20012 24508
rect 20012 24452 20016 24508
rect 19952 24448 20016 24452
rect 20032 24508 20096 24512
rect 20032 24452 20036 24508
rect 20036 24452 20092 24508
rect 20092 24452 20096 24508
rect 20032 24448 20096 24452
rect 20112 24508 20176 24512
rect 20112 24452 20116 24508
rect 20116 24452 20172 24508
rect 20172 24452 20176 24508
rect 20112 24448 20176 24452
rect 27646 24508 27710 24512
rect 27646 24452 27650 24508
rect 27650 24452 27706 24508
rect 27706 24452 27710 24508
rect 27646 24448 27710 24452
rect 27726 24508 27790 24512
rect 27726 24452 27730 24508
rect 27730 24452 27786 24508
rect 27786 24452 27790 24508
rect 27726 24448 27790 24452
rect 27806 24508 27870 24512
rect 27806 24452 27810 24508
rect 27810 24452 27866 24508
rect 27866 24452 27870 24508
rect 27806 24448 27870 24452
rect 27886 24508 27950 24512
rect 27886 24452 27890 24508
rect 27890 24452 27946 24508
rect 27946 24452 27950 24508
rect 27886 24448 27950 24452
rect 3664 23964 3728 23968
rect 3664 23908 3668 23964
rect 3668 23908 3724 23964
rect 3724 23908 3728 23964
rect 3664 23904 3728 23908
rect 3744 23964 3808 23968
rect 3744 23908 3748 23964
rect 3748 23908 3804 23964
rect 3804 23908 3808 23964
rect 3744 23904 3808 23908
rect 3824 23964 3888 23968
rect 3824 23908 3828 23964
rect 3828 23908 3884 23964
rect 3884 23908 3888 23964
rect 3824 23904 3888 23908
rect 3904 23964 3968 23968
rect 3904 23908 3908 23964
rect 3908 23908 3964 23964
rect 3964 23908 3968 23964
rect 3904 23904 3968 23908
rect 11438 23964 11502 23968
rect 11438 23908 11442 23964
rect 11442 23908 11498 23964
rect 11498 23908 11502 23964
rect 11438 23904 11502 23908
rect 11518 23964 11582 23968
rect 11518 23908 11522 23964
rect 11522 23908 11578 23964
rect 11578 23908 11582 23964
rect 11518 23904 11582 23908
rect 11598 23964 11662 23968
rect 11598 23908 11602 23964
rect 11602 23908 11658 23964
rect 11658 23908 11662 23964
rect 11598 23904 11662 23908
rect 11678 23964 11742 23968
rect 11678 23908 11682 23964
rect 11682 23908 11738 23964
rect 11738 23908 11742 23964
rect 11678 23904 11742 23908
rect 19212 23964 19276 23968
rect 19212 23908 19216 23964
rect 19216 23908 19272 23964
rect 19272 23908 19276 23964
rect 19212 23904 19276 23908
rect 19292 23964 19356 23968
rect 19292 23908 19296 23964
rect 19296 23908 19352 23964
rect 19352 23908 19356 23964
rect 19292 23904 19356 23908
rect 19372 23964 19436 23968
rect 19372 23908 19376 23964
rect 19376 23908 19432 23964
rect 19432 23908 19436 23964
rect 19372 23904 19436 23908
rect 19452 23964 19516 23968
rect 19452 23908 19456 23964
rect 19456 23908 19512 23964
rect 19512 23908 19516 23964
rect 19452 23904 19516 23908
rect 26986 23964 27050 23968
rect 26986 23908 26990 23964
rect 26990 23908 27046 23964
rect 27046 23908 27050 23964
rect 26986 23904 27050 23908
rect 27066 23964 27130 23968
rect 27066 23908 27070 23964
rect 27070 23908 27126 23964
rect 27126 23908 27130 23964
rect 27066 23904 27130 23908
rect 27146 23964 27210 23968
rect 27146 23908 27150 23964
rect 27150 23908 27206 23964
rect 27206 23908 27210 23964
rect 27146 23904 27210 23908
rect 27226 23964 27290 23968
rect 27226 23908 27230 23964
rect 27230 23908 27286 23964
rect 27286 23908 27290 23964
rect 27226 23904 27290 23908
rect 20484 23836 20548 23900
rect 4324 23420 4388 23424
rect 4324 23364 4328 23420
rect 4328 23364 4384 23420
rect 4384 23364 4388 23420
rect 4324 23360 4388 23364
rect 4404 23420 4468 23424
rect 4404 23364 4408 23420
rect 4408 23364 4464 23420
rect 4464 23364 4468 23420
rect 4404 23360 4468 23364
rect 4484 23420 4548 23424
rect 4484 23364 4488 23420
rect 4488 23364 4544 23420
rect 4544 23364 4548 23420
rect 4484 23360 4548 23364
rect 4564 23420 4628 23424
rect 4564 23364 4568 23420
rect 4568 23364 4624 23420
rect 4624 23364 4628 23420
rect 4564 23360 4628 23364
rect 12098 23420 12162 23424
rect 12098 23364 12102 23420
rect 12102 23364 12158 23420
rect 12158 23364 12162 23420
rect 12098 23360 12162 23364
rect 12178 23420 12242 23424
rect 12178 23364 12182 23420
rect 12182 23364 12238 23420
rect 12238 23364 12242 23420
rect 12178 23360 12242 23364
rect 12258 23420 12322 23424
rect 12258 23364 12262 23420
rect 12262 23364 12318 23420
rect 12318 23364 12322 23420
rect 12258 23360 12322 23364
rect 12338 23420 12402 23424
rect 12338 23364 12342 23420
rect 12342 23364 12398 23420
rect 12398 23364 12402 23420
rect 12338 23360 12402 23364
rect 19872 23420 19936 23424
rect 19872 23364 19876 23420
rect 19876 23364 19932 23420
rect 19932 23364 19936 23420
rect 19872 23360 19936 23364
rect 19952 23420 20016 23424
rect 19952 23364 19956 23420
rect 19956 23364 20012 23420
rect 20012 23364 20016 23420
rect 19952 23360 20016 23364
rect 20032 23420 20096 23424
rect 20032 23364 20036 23420
rect 20036 23364 20092 23420
rect 20092 23364 20096 23420
rect 20032 23360 20096 23364
rect 20112 23420 20176 23424
rect 20112 23364 20116 23420
rect 20116 23364 20172 23420
rect 20172 23364 20176 23420
rect 20112 23360 20176 23364
rect 27646 23420 27710 23424
rect 27646 23364 27650 23420
rect 27650 23364 27706 23420
rect 27706 23364 27710 23420
rect 27646 23360 27710 23364
rect 27726 23420 27790 23424
rect 27726 23364 27730 23420
rect 27730 23364 27786 23420
rect 27786 23364 27790 23420
rect 27726 23360 27790 23364
rect 27806 23420 27870 23424
rect 27806 23364 27810 23420
rect 27810 23364 27866 23420
rect 27866 23364 27870 23420
rect 27806 23360 27870 23364
rect 27886 23420 27950 23424
rect 27886 23364 27890 23420
rect 27890 23364 27946 23420
rect 27946 23364 27950 23420
rect 27886 23360 27950 23364
rect 3664 22876 3728 22880
rect 3664 22820 3668 22876
rect 3668 22820 3724 22876
rect 3724 22820 3728 22876
rect 3664 22816 3728 22820
rect 3744 22876 3808 22880
rect 3744 22820 3748 22876
rect 3748 22820 3804 22876
rect 3804 22820 3808 22876
rect 3744 22816 3808 22820
rect 3824 22876 3888 22880
rect 3824 22820 3828 22876
rect 3828 22820 3884 22876
rect 3884 22820 3888 22876
rect 3824 22816 3888 22820
rect 3904 22876 3968 22880
rect 3904 22820 3908 22876
rect 3908 22820 3964 22876
rect 3964 22820 3968 22876
rect 3904 22816 3968 22820
rect 11438 22876 11502 22880
rect 11438 22820 11442 22876
rect 11442 22820 11498 22876
rect 11498 22820 11502 22876
rect 11438 22816 11502 22820
rect 11518 22876 11582 22880
rect 11518 22820 11522 22876
rect 11522 22820 11578 22876
rect 11578 22820 11582 22876
rect 11518 22816 11582 22820
rect 11598 22876 11662 22880
rect 11598 22820 11602 22876
rect 11602 22820 11658 22876
rect 11658 22820 11662 22876
rect 11598 22816 11662 22820
rect 11678 22876 11742 22880
rect 11678 22820 11682 22876
rect 11682 22820 11738 22876
rect 11738 22820 11742 22876
rect 11678 22816 11742 22820
rect 19212 22876 19276 22880
rect 19212 22820 19216 22876
rect 19216 22820 19272 22876
rect 19272 22820 19276 22876
rect 19212 22816 19276 22820
rect 19292 22876 19356 22880
rect 19292 22820 19296 22876
rect 19296 22820 19352 22876
rect 19352 22820 19356 22876
rect 19292 22816 19356 22820
rect 19372 22876 19436 22880
rect 19372 22820 19376 22876
rect 19376 22820 19432 22876
rect 19432 22820 19436 22876
rect 19372 22816 19436 22820
rect 19452 22876 19516 22880
rect 19452 22820 19456 22876
rect 19456 22820 19512 22876
rect 19512 22820 19516 22876
rect 19452 22816 19516 22820
rect 26986 22876 27050 22880
rect 26986 22820 26990 22876
rect 26990 22820 27046 22876
rect 27046 22820 27050 22876
rect 26986 22816 27050 22820
rect 27066 22876 27130 22880
rect 27066 22820 27070 22876
rect 27070 22820 27126 22876
rect 27126 22820 27130 22876
rect 27066 22816 27130 22820
rect 27146 22876 27210 22880
rect 27146 22820 27150 22876
rect 27150 22820 27206 22876
rect 27206 22820 27210 22876
rect 27146 22816 27210 22820
rect 27226 22876 27290 22880
rect 27226 22820 27230 22876
rect 27230 22820 27286 22876
rect 27286 22820 27290 22876
rect 27226 22816 27290 22820
rect 4324 22332 4388 22336
rect 4324 22276 4328 22332
rect 4328 22276 4384 22332
rect 4384 22276 4388 22332
rect 4324 22272 4388 22276
rect 4404 22332 4468 22336
rect 4404 22276 4408 22332
rect 4408 22276 4464 22332
rect 4464 22276 4468 22332
rect 4404 22272 4468 22276
rect 4484 22332 4548 22336
rect 4484 22276 4488 22332
rect 4488 22276 4544 22332
rect 4544 22276 4548 22332
rect 4484 22272 4548 22276
rect 4564 22332 4628 22336
rect 4564 22276 4568 22332
rect 4568 22276 4624 22332
rect 4624 22276 4628 22332
rect 4564 22272 4628 22276
rect 12098 22332 12162 22336
rect 12098 22276 12102 22332
rect 12102 22276 12158 22332
rect 12158 22276 12162 22332
rect 12098 22272 12162 22276
rect 12178 22332 12242 22336
rect 12178 22276 12182 22332
rect 12182 22276 12238 22332
rect 12238 22276 12242 22332
rect 12178 22272 12242 22276
rect 12258 22332 12322 22336
rect 12258 22276 12262 22332
rect 12262 22276 12318 22332
rect 12318 22276 12322 22332
rect 12258 22272 12322 22276
rect 12338 22332 12402 22336
rect 12338 22276 12342 22332
rect 12342 22276 12398 22332
rect 12398 22276 12402 22332
rect 12338 22272 12402 22276
rect 19872 22332 19936 22336
rect 19872 22276 19876 22332
rect 19876 22276 19932 22332
rect 19932 22276 19936 22332
rect 19872 22272 19936 22276
rect 19952 22332 20016 22336
rect 19952 22276 19956 22332
rect 19956 22276 20012 22332
rect 20012 22276 20016 22332
rect 19952 22272 20016 22276
rect 20032 22332 20096 22336
rect 20032 22276 20036 22332
rect 20036 22276 20092 22332
rect 20092 22276 20096 22332
rect 20032 22272 20096 22276
rect 20112 22332 20176 22336
rect 20112 22276 20116 22332
rect 20116 22276 20172 22332
rect 20172 22276 20176 22332
rect 20112 22272 20176 22276
rect 27646 22332 27710 22336
rect 27646 22276 27650 22332
rect 27650 22276 27706 22332
rect 27706 22276 27710 22332
rect 27646 22272 27710 22276
rect 27726 22332 27790 22336
rect 27726 22276 27730 22332
rect 27730 22276 27786 22332
rect 27786 22276 27790 22332
rect 27726 22272 27790 22276
rect 27806 22332 27870 22336
rect 27806 22276 27810 22332
rect 27810 22276 27866 22332
rect 27866 22276 27870 22332
rect 27806 22272 27870 22276
rect 27886 22332 27950 22336
rect 27886 22276 27890 22332
rect 27890 22276 27946 22332
rect 27946 22276 27950 22332
rect 27886 22272 27950 22276
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 11438 21788 11502 21792
rect 11438 21732 11442 21788
rect 11442 21732 11498 21788
rect 11498 21732 11502 21788
rect 11438 21728 11502 21732
rect 11518 21788 11582 21792
rect 11518 21732 11522 21788
rect 11522 21732 11578 21788
rect 11578 21732 11582 21788
rect 11518 21728 11582 21732
rect 11598 21788 11662 21792
rect 11598 21732 11602 21788
rect 11602 21732 11658 21788
rect 11658 21732 11662 21788
rect 11598 21728 11662 21732
rect 11678 21788 11742 21792
rect 11678 21732 11682 21788
rect 11682 21732 11738 21788
rect 11738 21732 11742 21788
rect 11678 21728 11742 21732
rect 19212 21788 19276 21792
rect 19212 21732 19216 21788
rect 19216 21732 19272 21788
rect 19272 21732 19276 21788
rect 19212 21728 19276 21732
rect 19292 21788 19356 21792
rect 19292 21732 19296 21788
rect 19296 21732 19352 21788
rect 19352 21732 19356 21788
rect 19292 21728 19356 21732
rect 19372 21788 19436 21792
rect 19372 21732 19376 21788
rect 19376 21732 19432 21788
rect 19432 21732 19436 21788
rect 19372 21728 19436 21732
rect 19452 21788 19516 21792
rect 19452 21732 19456 21788
rect 19456 21732 19512 21788
rect 19512 21732 19516 21788
rect 19452 21728 19516 21732
rect 26986 21788 27050 21792
rect 26986 21732 26990 21788
rect 26990 21732 27046 21788
rect 27046 21732 27050 21788
rect 26986 21728 27050 21732
rect 27066 21788 27130 21792
rect 27066 21732 27070 21788
rect 27070 21732 27126 21788
rect 27126 21732 27130 21788
rect 27066 21728 27130 21732
rect 27146 21788 27210 21792
rect 27146 21732 27150 21788
rect 27150 21732 27206 21788
rect 27206 21732 27210 21788
rect 27146 21728 27210 21732
rect 27226 21788 27290 21792
rect 27226 21732 27230 21788
rect 27230 21732 27286 21788
rect 27286 21732 27290 21788
rect 27226 21728 27290 21732
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 12098 21244 12162 21248
rect 12098 21188 12102 21244
rect 12102 21188 12158 21244
rect 12158 21188 12162 21244
rect 12098 21184 12162 21188
rect 12178 21244 12242 21248
rect 12178 21188 12182 21244
rect 12182 21188 12238 21244
rect 12238 21188 12242 21244
rect 12178 21184 12242 21188
rect 12258 21244 12322 21248
rect 12258 21188 12262 21244
rect 12262 21188 12318 21244
rect 12318 21188 12322 21244
rect 12258 21184 12322 21188
rect 12338 21244 12402 21248
rect 12338 21188 12342 21244
rect 12342 21188 12398 21244
rect 12398 21188 12402 21244
rect 12338 21184 12402 21188
rect 19872 21244 19936 21248
rect 19872 21188 19876 21244
rect 19876 21188 19932 21244
rect 19932 21188 19936 21244
rect 19872 21184 19936 21188
rect 19952 21244 20016 21248
rect 19952 21188 19956 21244
rect 19956 21188 20012 21244
rect 20012 21188 20016 21244
rect 19952 21184 20016 21188
rect 20032 21244 20096 21248
rect 20032 21188 20036 21244
rect 20036 21188 20092 21244
rect 20092 21188 20096 21244
rect 20032 21184 20096 21188
rect 20112 21244 20176 21248
rect 20112 21188 20116 21244
rect 20116 21188 20172 21244
rect 20172 21188 20176 21244
rect 20112 21184 20176 21188
rect 27646 21244 27710 21248
rect 27646 21188 27650 21244
rect 27650 21188 27706 21244
rect 27706 21188 27710 21244
rect 27646 21184 27710 21188
rect 27726 21244 27790 21248
rect 27726 21188 27730 21244
rect 27730 21188 27786 21244
rect 27786 21188 27790 21244
rect 27726 21184 27790 21188
rect 27806 21244 27870 21248
rect 27806 21188 27810 21244
rect 27810 21188 27866 21244
rect 27866 21188 27870 21244
rect 27806 21184 27870 21188
rect 27886 21244 27950 21248
rect 27886 21188 27890 21244
rect 27890 21188 27946 21244
rect 27946 21188 27950 21244
rect 27886 21184 27950 21188
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 11438 20700 11502 20704
rect 11438 20644 11442 20700
rect 11442 20644 11498 20700
rect 11498 20644 11502 20700
rect 11438 20640 11502 20644
rect 11518 20700 11582 20704
rect 11518 20644 11522 20700
rect 11522 20644 11578 20700
rect 11578 20644 11582 20700
rect 11518 20640 11582 20644
rect 11598 20700 11662 20704
rect 11598 20644 11602 20700
rect 11602 20644 11658 20700
rect 11658 20644 11662 20700
rect 11598 20640 11662 20644
rect 11678 20700 11742 20704
rect 11678 20644 11682 20700
rect 11682 20644 11738 20700
rect 11738 20644 11742 20700
rect 11678 20640 11742 20644
rect 19212 20700 19276 20704
rect 19212 20644 19216 20700
rect 19216 20644 19272 20700
rect 19272 20644 19276 20700
rect 19212 20640 19276 20644
rect 19292 20700 19356 20704
rect 19292 20644 19296 20700
rect 19296 20644 19352 20700
rect 19352 20644 19356 20700
rect 19292 20640 19356 20644
rect 19372 20700 19436 20704
rect 19372 20644 19376 20700
rect 19376 20644 19432 20700
rect 19432 20644 19436 20700
rect 19372 20640 19436 20644
rect 19452 20700 19516 20704
rect 19452 20644 19456 20700
rect 19456 20644 19512 20700
rect 19512 20644 19516 20700
rect 19452 20640 19516 20644
rect 26986 20700 27050 20704
rect 26986 20644 26990 20700
rect 26990 20644 27046 20700
rect 27046 20644 27050 20700
rect 26986 20640 27050 20644
rect 27066 20700 27130 20704
rect 27066 20644 27070 20700
rect 27070 20644 27126 20700
rect 27126 20644 27130 20700
rect 27066 20640 27130 20644
rect 27146 20700 27210 20704
rect 27146 20644 27150 20700
rect 27150 20644 27206 20700
rect 27206 20644 27210 20700
rect 27146 20640 27210 20644
rect 27226 20700 27290 20704
rect 27226 20644 27230 20700
rect 27230 20644 27286 20700
rect 27286 20644 27290 20700
rect 27226 20640 27290 20644
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 12098 20156 12162 20160
rect 12098 20100 12102 20156
rect 12102 20100 12158 20156
rect 12158 20100 12162 20156
rect 12098 20096 12162 20100
rect 12178 20156 12242 20160
rect 12178 20100 12182 20156
rect 12182 20100 12238 20156
rect 12238 20100 12242 20156
rect 12178 20096 12242 20100
rect 12258 20156 12322 20160
rect 12258 20100 12262 20156
rect 12262 20100 12318 20156
rect 12318 20100 12322 20156
rect 12258 20096 12322 20100
rect 12338 20156 12402 20160
rect 12338 20100 12342 20156
rect 12342 20100 12398 20156
rect 12398 20100 12402 20156
rect 12338 20096 12402 20100
rect 19872 20156 19936 20160
rect 19872 20100 19876 20156
rect 19876 20100 19932 20156
rect 19932 20100 19936 20156
rect 19872 20096 19936 20100
rect 19952 20156 20016 20160
rect 19952 20100 19956 20156
rect 19956 20100 20012 20156
rect 20012 20100 20016 20156
rect 19952 20096 20016 20100
rect 20032 20156 20096 20160
rect 20032 20100 20036 20156
rect 20036 20100 20092 20156
rect 20092 20100 20096 20156
rect 20032 20096 20096 20100
rect 20112 20156 20176 20160
rect 20112 20100 20116 20156
rect 20116 20100 20172 20156
rect 20172 20100 20176 20156
rect 20112 20096 20176 20100
rect 27646 20156 27710 20160
rect 27646 20100 27650 20156
rect 27650 20100 27706 20156
rect 27706 20100 27710 20156
rect 27646 20096 27710 20100
rect 27726 20156 27790 20160
rect 27726 20100 27730 20156
rect 27730 20100 27786 20156
rect 27786 20100 27790 20156
rect 27726 20096 27790 20100
rect 27806 20156 27870 20160
rect 27806 20100 27810 20156
rect 27810 20100 27866 20156
rect 27866 20100 27870 20156
rect 27806 20096 27870 20100
rect 27886 20156 27950 20160
rect 27886 20100 27890 20156
rect 27890 20100 27946 20156
rect 27946 20100 27950 20156
rect 27886 20096 27950 20100
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 11438 19612 11502 19616
rect 11438 19556 11442 19612
rect 11442 19556 11498 19612
rect 11498 19556 11502 19612
rect 11438 19552 11502 19556
rect 11518 19612 11582 19616
rect 11518 19556 11522 19612
rect 11522 19556 11578 19612
rect 11578 19556 11582 19612
rect 11518 19552 11582 19556
rect 11598 19612 11662 19616
rect 11598 19556 11602 19612
rect 11602 19556 11658 19612
rect 11658 19556 11662 19612
rect 11598 19552 11662 19556
rect 11678 19612 11742 19616
rect 11678 19556 11682 19612
rect 11682 19556 11738 19612
rect 11738 19556 11742 19612
rect 11678 19552 11742 19556
rect 19212 19612 19276 19616
rect 19212 19556 19216 19612
rect 19216 19556 19272 19612
rect 19272 19556 19276 19612
rect 19212 19552 19276 19556
rect 19292 19612 19356 19616
rect 19292 19556 19296 19612
rect 19296 19556 19352 19612
rect 19352 19556 19356 19612
rect 19292 19552 19356 19556
rect 19372 19612 19436 19616
rect 19372 19556 19376 19612
rect 19376 19556 19432 19612
rect 19432 19556 19436 19612
rect 19372 19552 19436 19556
rect 19452 19612 19516 19616
rect 19452 19556 19456 19612
rect 19456 19556 19512 19612
rect 19512 19556 19516 19612
rect 19452 19552 19516 19556
rect 26986 19612 27050 19616
rect 26986 19556 26990 19612
rect 26990 19556 27046 19612
rect 27046 19556 27050 19612
rect 26986 19552 27050 19556
rect 27066 19612 27130 19616
rect 27066 19556 27070 19612
rect 27070 19556 27126 19612
rect 27126 19556 27130 19612
rect 27066 19552 27130 19556
rect 27146 19612 27210 19616
rect 27146 19556 27150 19612
rect 27150 19556 27206 19612
rect 27206 19556 27210 19612
rect 27146 19552 27210 19556
rect 27226 19612 27290 19616
rect 27226 19556 27230 19612
rect 27230 19556 27286 19612
rect 27286 19556 27290 19612
rect 27226 19552 27290 19556
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 12098 19068 12162 19072
rect 12098 19012 12102 19068
rect 12102 19012 12158 19068
rect 12158 19012 12162 19068
rect 12098 19008 12162 19012
rect 12178 19068 12242 19072
rect 12178 19012 12182 19068
rect 12182 19012 12238 19068
rect 12238 19012 12242 19068
rect 12178 19008 12242 19012
rect 12258 19068 12322 19072
rect 12258 19012 12262 19068
rect 12262 19012 12318 19068
rect 12318 19012 12322 19068
rect 12258 19008 12322 19012
rect 12338 19068 12402 19072
rect 12338 19012 12342 19068
rect 12342 19012 12398 19068
rect 12398 19012 12402 19068
rect 12338 19008 12402 19012
rect 19872 19068 19936 19072
rect 19872 19012 19876 19068
rect 19876 19012 19932 19068
rect 19932 19012 19936 19068
rect 19872 19008 19936 19012
rect 19952 19068 20016 19072
rect 19952 19012 19956 19068
rect 19956 19012 20012 19068
rect 20012 19012 20016 19068
rect 19952 19008 20016 19012
rect 20032 19068 20096 19072
rect 20032 19012 20036 19068
rect 20036 19012 20092 19068
rect 20092 19012 20096 19068
rect 20032 19008 20096 19012
rect 20112 19068 20176 19072
rect 20112 19012 20116 19068
rect 20116 19012 20172 19068
rect 20172 19012 20176 19068
rect 20112 19008 20176 19012
rect 27646 19068 27710 19072
rect 27646 19012 27650 19068
rect 27650 19012 27706 19068
rect 27706 19012 27710 19068
rect 27646 19008 27710 19012
rect 27726 19068 27790 19072
rect 27726 19012 27730 19068
rect 27730 19012 27786 19068
rect 27786 19012 27790 19068
rect 27726 19008 27790 19012
rect 27806 19068 27870 19072
rect 27806 19012 27810 19068
rect 27810 19012 27866 19068
rect 27866 19012 27870 19068
rect 27806 19008 27870 19012
rect 27886 19068 27950 19072
rect 27886 19012 27890 19068
rect 27890 19012 27946 19068
rect 27946 19012 27950 19068
rect 27886 19008 27950 19012
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 11438 18524 11502 18528
rect 11438 18468 11442 18524
rect 11442 18468 11498 18524
rect 11498 18468 11502 18524
rect 11438 18464 11502 18468
rect 11518 18524 11582 18528
rect 11518 18468 11522 18524
rect 11522 18468 11578 18524
rect 11578 18468 11582 18524
rect 11518 18464 11582 18468
rect 11598 18524 11662 18528
rect 11598 18468 11602 18524
rect 11602 18468 11658 18524
rect 11658 18468 11662 18524
rect 11598 18464 11662 18468
rect 11678 18524 11742 18528
rect 11678 18468 11682 18524
rect 11682 18468 11738 18524
rect 11738 18468 11742 18524
rect 11678 18464 11742 18468
rect 19212 18524 19276 18528
rect 19212 18468 19216 18524
rect 19216 18468 19272 18524
rect 19272 18468 19276 18524
rect 19212 18464 19276 18468
rect 19292 18524 19356 18528
rect 19292 18468 19296 18524
rect 19296 18468 19352 18524
rect 19352 18468 19356 18524
rect 19292 18464 19356 18468
rect 19372 18524 19436 18528
rect 19372 18468 19376 18524
rect 19376 18468 19432 18524
rect 19432 18468 19436 18524
rect 19372 18464 19436 18468
rect 19452 18524 19516 18528
rect 19452 18468 19456 18524
rect 19456 18468 19512 18524
rect 19512 18468 19516 18524
rect 19452 18464 19516 18468
rect 26986 18524 27050 18528
rect 26986 18468 26990 18524
rect 26990 18468 27046 18524
rect 27046 18468 27050 18524
rect 26986 18464 27050 18468
rect 27066 18524 27130 18528
rect 27066 18468 27070 18524
rect 27070 18468 27126 18524
rect 27126 18468 27130 18524
rect 27066 18464 27130 18468
rect 27146 18524 27210 18528
rect 27146 18468 27150 18524
rect 27150 18468 27206 18524
rect 27206 18468 27210 18524
rect 27146 18464 27210 18468
rect 27226 18524 27290 18528
rect 27226 18468 27230 18524
rect 27230 18468 27286 18524
rect 27286 18468 27290 18524
rect 27226 18464 27290 18468
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 12098 17980 12162 17984
rect 12098 17924 12102 17980
rect 12102 17924 12158 17980
rect 12158 17924 12162 17980
rect 12098 17920 12162 17924
rect 12178 17980 12242 17984
rect 12178 17924 12182 17980
rect 12182 17924 12238 17980
rect 12238 17924 12242 17980
rect 12178 17920 12242 17924
rect 12258 17980 12322 17984
rect 12258 17924 12262 17980
rect 12262 17924 12318 17980
rect 12318 17924 12322 17980
rect 12258 17920 12322 17924
rect 12338 17980 12402 17984
rect 12338 17924 12342 17980
rect 12342 17924 12398 17980
rect 12398 17924 12402 17980
rect 12338 17920 12402 17924
rect 19872 17980 19936 17984
rect 19872 17924 19876 17980
rect 19876 17924 19932 17980
rect 19932 17924 19936 17980
rect 19872 17920 19936 17924
rect 19952 17980 20016 17984
rect 19952 17924 19956 17980
rect 19956 17924 20012 17980
rect 20012 17924 20016 17980
rect 19952 17920 20016 17924
rect 20032 17980 20096 17984
rect 20032 17924 20036 17980
rect 20036 17924 20092 17980
rect 20092 17924 20096 17980
rect 20032 17920 20096 17924
rect 20112 17980 20176 17984
rect 20112 17924 20116 17980
rect 20116 17924 20172 17980
rect 20172 17924 20176 17980
rect 20112 17920 20176 17924
rect 27646 17980 27710 17984
rect 27646 17924 27650 17980
rect 27650 17924 27706 17980
rect 27706 17924 27710 17980
rect 27646 17920 27710 17924
rect 27726 17980 27790 17984
rect 27726 17924 27730 17980
rect 27730 17924 27786 17980
rect 27786 17924 27790 17980
rect 27726 17920 27790 17924
rect 27806 17980 27870 17984
rect 27806 17924 27810 17980
rect 27810 17924 27866 17980
rect 27866 17924 27870 17980
rect 27806 17920 27870 17924
rect 27886 17980 27950 17984
rect 27886 17924 27890 17980
rect 27890 17924 27946 17980
rect 27946 17924 27950 17980
rect 27886 17920 27950 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 11438 17436 11502 17440
rect 11438 17380 11442 17436
rect 11442 17380 11498 17436
rect 11498 17380 11502 17436
rect 11438 17376 11502 17380
rect 11518 17436 11582 17440
rect 11518 17380 11522 17436
rect 11522 17380 11578 17436
rect 11578 17380 11582 17436
rect 11518 17376 11582 17380
rect 11598 17436 11662 17440
rect 11598 17380 11602 17436
rect 11602 17380 11658 17436
rect 11658 17380 11662 17436
rect 11598 17376 11662 17380
rect 11678 17436 11742 17440
rect 11678 17380 11682 17436
rect 11682 17380 11738 17436
rect 11738 17380 11742 17436
rect 11678 17376 11742 17380
rect 19212 17436 19276 17440
rect 19212 17380 19216 17436
rect 19216 17380 19272 17436
rect 19272 17380 19276 17436
rect 19212 17376 19276 17380
rect 19292 17436 19356 17440
rect 19292 17380 19296 17436
rect 19296 17380 19352 17436
rect 19352 17380 19356 17436
rect 19292 17376 19356 17380
rect 19372 17436 19436 17440
rect 19372 17380 19376 17436
rect 19376 17380 19432 17436
rect 19432 17380 19436 17436
rect 19372 17376 19436 17380
rect 19452 17436 19516 17440
rect 19452 17380 19456 17436
rect 19456 17380 19512 17436
rect 19512 17380 19516 17436
rect 19452 17376 19516 17380
rect 26986 17436 27050 17440
rect 26986 17380 26990 17436
rect 26990 17380 27046 17436
rect 27046 17380 27050 17436
rect 26986 17376 27050 17380
rect 27066 17436 27130 17440
rect 27066 17380 27070 17436
rect 27070 17380 27126 17436
rect 27126 17380 27130 17436
rect 27066 17376 27130 17380
rect 27146 17436 27210 17440
rect 27146 17380 27150 17436
rect 27150 17380 27206 17436
rect 27206 17380 27210 17436
rect 27146 17376 27210 17380
rect 27226 17436 27290 17440
rect 27226 17380 27230 17436
rect 27230 17380 27286 17436
rect 27286 17380 27290 17436
rect 27226 17376 27290 17380
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 12098 16892 12162 16896
rect 12098 16836 12102 16892
rect 12102 16836 12158 16892
rect 12158 16836 12162 16892
rect 12098 16832 12162 16836
rect 12178 16892 12242 16896
rect 12178 16836 12182 16892
rect 12182 16836 12238 16892
rect 12238 16836 12242 16892
rect 12178 16832 12242 16836
rect 12258 16892 12322 16896
rect 12258 16836 12262 16892
rect 12262 16836 12318 16892
rect 12318 16836 12322 16892
rect 12258 16832 12322 16836
rect 12338 16892 12402 16896
rect 12338 16836 12342 16892
rect 12342 16836 12398 16892
rect 12398 16836 12402 16892
rect 12338 16832 12402 16836
rect 19872 16892 19936 16896
rect 19872 16836 19876 16892
rect 19876 16836 19932 16892
rect 19932 16836 19936 16892
rect 19872 16832 19936 16836
rect 19952 16892 20016 16896
rect 19952 16836 19956 16892
rect 19956 16836 20012 16892
rect 20012 16836 20016 16892
rect 19952 16832 20016 16836
rect 20032 16892 20096 16896
rect 20032 16836 20036 16892
rect 20036 16836 20092 16892
rect 20092 16836 20096 16892
rect 20032 16832 20096 16836
rect 20112 16892 20176 16896
rect 20112 16836 20116 16892
rect 20116 16836 20172 16892
rect 20172 16836 20176 16892
rect 20112 16832 20176 16836
rect 27646 16892 27710 16896
rect 27646 16836 27650 16892
rect 27650 16836 27706 16892
rect 27706 16836 27710 16892
rect 27646 16832 27710 16836
rect 27726 16892 27790 16896
rect 27726 16836 27730 16892
rect 27730 16836 27786 16892
rect 27786 16836 27790 16892
rect 27726 16832 27790 16836
rect 27806 16892 27870 16896
rect 27806 16836 27810 16892
rect 27810 16836 27866 16892
rect 27866 16836 27870 16892
rect 27806 16832 27870 16836
rect 27886 16892 27950 16896
rect 27886 16836 27890 16892
rect 27890 16836 27946 16892
rect 27946 16836 27950 16892
rect 27886 16832 27950 16836
rect 26740 16628 26804 16692
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 11438 16348 11502 16352
rect 11438 16292 11442 16348
rect 11442 16292 11498 16348
rect 11498 16292 11502 16348
rect 11438 16288 11502 16292
rect 11518 16348 11582 16352
rect 11518 16292 11522 16348
rect 11522 16292 11578 16348
rect 11578 16292 11582 16348
rect 11518 16288 11582 16292
rect 11598 16348 11662 16352
rect 11598 16292 11602 16348
rect 11602 16292 11658 16348
rect 11658 16292 11662 16348
rect 11598 16288 11662 16292
rect 11678 16348 11742 16352
rect 11678 16292 11682 16348
rect 11682 16292 11738 16348
rect 11738 16292 11742 16348
rect 11678 16288 11742 16292
rect 19212 16348 19276 16352
rect 19212 16292 19216 16348
rect 19216 16292 19272 16348
rect 19272 16292 19276 16348
rect 19212 16288 19276 16292
rect 19292 16348 19356 16352
rect 19292 16292 19296 16348
rect 19296 16292 19352 16348
rect 19352 16292 19356 16348
rect 19292 16288 19356 16292
rect 19372 16348 19436 16352
rect 19372 16292 19376 16348
rect 19376 16292 19432 16348
rect 19432 16292 19436 16348
rect 19372 16288 19436 16292
rect 19452 16348 19516 16352
rect 19452 16292 19456 16348
rect 19456 16292 19512 16348
rect 19512 16292 19516 16348
rect 19452 16288 19516 16292
rect 26986 16348 27050 16352
rect 26986 16292 26990 16348
rect 26990 16292 27046 16348
rect 27046 16292 27050 16348
rect 26986 16288 27050 16292
rect 27066 16348 27130 16352
rect 27066 16292 27070 16348
rect 27070 16292 27126 16348
rect 27126 16292 27130 16348
rect 27066 16288 27130 16292
rect 27146 16348 27210 16352
rect 27146 16292 27150 16348
rect 27150 16292 27206 16348
rect 27206 16292 27210 16348
rect 27146 16288 27210 16292
rect 27226 16348 27290 16352
rect 27226 16292 27230 16348
rect 27230 16292 27286 16348
rect 27286 16292 27290 16348
rect 27226 16288 27290 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 12098 15804 12162 15808
rect 12098 15748 12102 15804
rect 12102 15748 12158 15804
rect 12158 15748 12162 15804
rect 12098 15744 12162 15748
rect 12178 15804 12242 15808
rect 12178 15748 12182 15804
rect 12182 15748 12238 15804
rect 12238 15748 12242 15804
rect 12178 15744 12242 15748
rect 12258 15804 12322 15808
rect 12258 15748 12262 15804
rect 12262 15748 12318 15804
rect 12318 15748 12322 15804
rect 12258 15744 12322 15748
rect 12338 15804 12402 15808
rect 12338 15748 12342 15804
rect 12342 15748 12398 15804
rect 12398 15748 12402 15804
rect 12338 15744 12402 15748
rect 19872 15804 19936 15808
rect 19872 15748 19876 15804
rect 19876 15748 19932 15804
rect 19932 15748 19936 15804
rect 19872 15744 19936 15748
rect 19952 15804 20016 15808
rect 19952 15748 19956 15804
rect 19956 15748 20012 15804
rect 20012 15748 20016 15804
rect 19952 15744 20016 15748
rect 20032 15804 20096 15808
rect 20032 15748 20036 15804
rect 20036 15748 20092 15804
rect 20092 15748 20096 15804
rect 20032 15744 20096 15748
rect 20112 15804 20176 15808
rect 20112 15748 20116 15804
rect 20116 15748 20172 15804
rect 20172 15748 20176 15804
rect 20112 15744 20176 15748
rect 27646 15804 27710 15808
rect 27646 15748 27650 15804
rect 27650 15748 27706 15804
rect 27706 15748 27710 15804
rect 27646 15744 27710 15748
rect 27726 15804 27790 15808
rect 27726 15748 27730 15804
rect 27730 15748 27786 15804
rect 27786 15748 27790 15804
rect 27726 15744 27790 15748
rect 27806 15804 27870 15808
rect 27806 15748 27810 15804
rect 27810 15748 27866 15804
rect 27866 15748 27870 15804
rect 27806 15744 27870 15748
rect 27886 15804 27950 15808
rect 27886 15748 27890 15804
rect 27890 15748 27946 15804
rect 27946 15748 27950 15804
rect 27886 15744 27950 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 11438 15260 11502 15264
rect 11438 15204 11442 15260
rect 11442 15204 11498 15260
rect 11498 15204 11502 15260
rect 11438 15200 11502 15204
rect 11518 15260 11582 15264
rect 11518 15204 11522 15260
rect 11522 15204 11578 15260
rect 11578 15204 11582 15260
rect 11518 15200 11582 15204
rect 11598 15260 11662 15264
rect 11598 15204 11602 15260
rect 11602 15204 11658 15260
rect 11658 15204 11662 15260
rect 11598 15200 11662 15204
rect 11678 15260 11742 15264
rect 11678 15204 11682 15260
rect 11682 15204 11738 15260
rect 11738 15204 11742 15260
rect 11678 15200 11742 15204
rect 19212 15260 19276 15264
rect 19212 15204 19216 15260
rect 19216 15204 19272 15260
rect 19272 15204 19276 15260
rect 19212 15200 19276 15204
rect 19292 15260 19356 15264
rect 19292 15204 19296 15260
rect 19296 15204 19352 15260
rect 19352 15204 19356 15260
rect 19292 15200 19356 15204
rect 19372 15260 19436 15264
rect 19372 15204 19376 15260
rect 19376 15204 19432 15260
rect 19432 15204 19436 15260
rect 19372 15200 19436 15204
rect 19452 15260 19516 15264
rect 19452 15204 19456 15260
rect 19456 15204 19512 15260
rect 19512 15204 19516 15260
rect 19452 15200 19516 15204
rect 26986 15260 27050 15264
rect 26986 15204 26990 15260
rect 26990 15204 27046 15260
rect 27046 15204 27050 15260
rect 26986 15200 27050 15204
rect 27066 15260 27130 15264
rect 27066 15204 27070 15260
rect 27070 15204 27126 15260
rect 27126 15204 27130 15260
rect 27066 15200 27130 15204
rect 27146 15260 27210 15264
rect 27146 15204 27150 15260
rect 27150 15204 27206 15260
rect 27206 15204 27210 15260
rect 27146 15200 27210 15204
rect 27226 15260 27290 15264
rect 27226 15204 27230 15260
rect 27230 15204 27286 15260
rect 27286 15204 27290 15260
rect 27226 15200 27290 15204
rect 16988 15192 17052 15196
rect 16988 15136 17002 15192
rect 17002 15136 17052 15192
rect 16988 15132 17052 15136
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 12098 14716 12162 14720
rect 12098 14660 12102 14716
rect 12102 14660 12158 14716
rect 12158 14660 12162 14716
rect 12098 14656 12162 14660
rect 12178 14716 12242 14720
rect 12178 14660 12182 14716
rect 12182 14660 12238 14716
rect 12238 14660 12242 14716
rect 12178 14656 12242 14660
rect 12258 14716 12322 14720
rect 12258 14660 12262 14716
rect 12262 14660 12318 14716
rect 12318 14660 12322 14716
rect 12258 14656 12322 14660
rect 12338 14716 12402 14720
rect 12338 14660 12342 14716
rect 12342 14660 12398 14716
rect 12398 14660 12402 14716
rect 12338 14656 12402 14660
rect 19872 14716 19936 14720
rect 19872 14660 19876 14716
rect 19876 14660 19932 14716
rect 19932 14660 19936 14716
rect 19872 14656 19936 14660
rect 19952 14716 20016 14720
rect 19952 14660 19956 14716
rect 19956 14660 20012 14716
rect 20012 14660 20016 14716
rect 19952 14656 20016 14660
rect 20032 14716 20096 14720
rect 20032 14660 20036 14716
rect 20036 14660 20092 14716
rect 20092 14660 20096 14716
rect 20032 14656 20096 14660
rect 20112 14716 20176 14720
rect 20112 14660 20116 14716
rect 20116 14660 20172 14716
rect 20172 14660 20176 14716
rect 20112 14656 20176 14660
rect 27646 14716 27710 14720
rect 27646 14660 27650 14716
rect 27650 14660 27706 14716
rect 27706 14660 27710 14716
rect 27646 14656 27710 14660
rect 27726 14716 27790 14720
rect 27726 14660 27730 14716
rect 27730 14660 27786 14716
rect 27786 14660 27790 14716
rect 27726 14656 27790 14660
rect 27806 14716 27870 14720
rect 27806 14660 27810 14716
rect 27810 14660 27866 14716
rect 27866 14660 27870 14716
rect 27806 14656 27870 14660
rect 27886 14716 27950 14720
rect 27886 14660 27890 14716
rect 27890 14660 27946 14716
rect 27946 14660 27950 14716
rect 27886 14656 27950 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 11438 14172 11502 14176
rect 11438 14116 11442 14172
rect 11442 14116 11498 14172
rect 11498 14116 11502 14172
rect 11438 14112 11502 14116
rect 11518 14172 11582 14176
rect 11518 14116 11522 14172
rect 11522 14116 11578 14172
rect 11578 14116 11582 14172
rect 11518 14112 11582 14116
rect 11598 14172 11662 14176
rect 11598 14116 11602 14172
rect 11602 14116 11658 14172
rect 11658 14116 11662 14172
rect 11598 14112 11662 14116
rect 11678 14172 11742 14176
rect 11678 14116 11682 14172
rect 11682 14116 11738 14172
rect 11738 14116 11742 14172
rect 11678 14112 11742 14116
rect 19212 14172 19276 14176
rect 19212 14116 19216 14172
rect 19216 14116 19272 14172
rect 19272 14116 19276 14172
rect 19212 14112 19276 14116
rect 19292 14172 19356 14176
rect 19292 14116 19296 14172
rect 19296 14116 19352 14172
rect 19352 14116 19356 14172
rect 19292 14112 19356 14116
rect 19372 14172 19436 14176
rect 19372 14116 19376 14172
rect 19376 14116 19432 14172
rect 19432 14116 19436 14172
rect 19372 14112 19436 14116
rect 19452 14172 19516 14176
rect 19452 14116 19456 14172
rect 19456 14116 19512 14172
rect 19512 14116 19516 14172
rect 19452 14112 19516 14116
rect 26986 14172 27050 14176
rect 26986 14116 26990 14172
rect 26990 14116 27046 14172
rect 27046 14116 27050 14172
rect 26986 14112 27050 14116
rect 27066 14172 27130 14176
rect 27066 14116 27070 14172
rect 27070 14116 27126 14172
rect 27126 14116 27130 14172
rect 27066 14112 27130 14116
rect 27146 14172 27210 14176
rect 27146 14116 27150 14172
rect 27150 14116 27206 14172
rect 27206 14116 27210 14172
rect 27146 14112 27210 14116
rect 27226 14172 27290 14176
rect 27226 14116 27230 14172
rect 27230 14116 27286 14172
rect 27286 14116 27290 14172
rect 27226 14112 27290 14116
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 12098 13628 12162 13632
rect 12098 13572 12102 13628
rect 12102 13572 12158 13628
rect 12158 13572 12162 13628
rect 12098 13568 12162 13572
rect 12178 13628 12242 13632
rect 12178 13572 12182 13628
rect 12182 13572 12238 13628
rect 12238 13572 12242 13628
rect 12178 13568 12242 13572
rect 12258 13628 12322 13632
rect 12258 13572 12262 13628
rect 12262 13572 12318 13628
rect 12318 13572 12322 13628
rect 12258 13568 12322 13572
rect 12338 13628 12402 13632
rect 12338 13572 12342 13628
rect 12342 13572 12398 13628
rect 12398 13572 12402 13628
rect 12338 13568 12402 13572
rect 19872 13628 19936 13632
rect 19872 13572 19876 13628
rect 19876 13572 19932 13628
rect 19932 13572 19936 13628
rect 19872 13568 19936 13572
rect 19952 13628 20016 13632
rect 19952 13572 19956 13628
rect 19956 13572 20012 13628
rect 20012 13572 20016 13628
rect 19952 13568 20016 13572
rect 20032 13628 20096 13632
rect 20032 13572 20036 13628
rect 20036 13572 20092 13628
rect 20092 13572 20096 13628
rect 20032 13568 20096 13572
rect 20112 13628 20176 13632
rect 20112 13572 20116 13628
rect 20116 13572 20172 13628
rect 20172 13572 20176 13628
rect 20112 13568 20176 13572
rect 27646 13628 27710 13632
rect 27646 13572 27650 13628
rect 27650 13572 27706 13628
rect 27706 13572 27710 13628
rect 27646 13568 27710 13572
rect 27726 13628 27790 13632
rect 27726 13572 27730 13628
rect 27730 13572 27786 13628
rect 27786 13572 27790 13628
rect 27726 13568 27790 13572
rect 27806 13628 27870 13632
rect 27806 13572 27810 13628
rect 27810 13572 27866 13628
rect 27866 13572 27870 13628
rect 27806 13568 27870 13572
rect 27886 13628 27950 13632
rect 27886 13572 27890 13628
rect 27890 13572 27946 13628
rect 27946 13572 27950 13628
rect 27886 13568 27950 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 11438 13084 11502 13088
rect 11438 13028 11442 13084
rect 11442 13028 11498 13084
rect 11498 13028 11502 13084
rect 11438 13024 11502 13028
rect 11518 13084 11582 13088
rect 11518 13028 11522 13084
rect 11522 13028 11578 13084
rect 11578 13028 11582 13084
rect 11518 13024 11582 13028
rect 11598 13084 11662 13088
rect 11598 13028 11602 13084
rect 11602 13028 11658 13084
rect 11658 13028 11662 13084
rect 11598 13024 11662 13028
rect 11678 13084 11742 13088
rect 11678 13028 11682 13084
rect 11682 13028 11738 13084
rect 11738 13028 11742 13084
rect 11678 13024 11742 13028
rect 19212 13084 19276 13088
rect 19212 13028 19216 13084
rect 19216 13028 19272 13084
rect 19272 13028 19276 13084
rect 19212 13024 19276 13028
rect 19292 13084 19356 13088
rect 19292 13028 19296 13084
rect 19296 13028 19352 13084
rect 19352 13028 19356 13084
rect 19292 13024 19356 13028
rect 19372 13084 19436 13088
rect 19372 13028 19376 13084
rect 19376 13028 19432 13084
rect 19432 13028 19436 13084
rect 19372 13024 19436 13028
rect 19452 13084 19516 13088
rect 19452 13028 19456 13084
rect 19456 13028 19512 13084
rect 19512 13028 19516 13084
rect 19452 13024 19516 13028
rect 26986 13084 27050 13088
rect 26986 13028 26990 13084
rect 26990 13028 27046 13084
rect 27046 13028 27050 13084
rect 26986 13024 27050 13028
rect 27066 13084 27130 13088
rect 27066 13028 27070 13084
rect 27070 13028 27126 13084
rect 27126 13028 27130 13084
rect 27066 13024 27130 13028
rect 27146 13084 27210 13088
rect 27146 13028 27150 13084
rect 27150 13028 27206 13084
rect 27206 13028 27210 13084
rect 27146 13024 27210 13028
rect 27226 13084 27290 13088
rect 27226 13028 27230 13084
rect 27230 13028 27286 13084
rect 27286 13028 27290 13084
rect 27226 13024 27290 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 12098 12540 12162 12544
rect 12098 12484 12102 12540
rect 12102 12484 12158 12540
rect 12158 12484 12162 12540
rect 12098 12480 12162 12484
rect 12178 12540 12242 12544
rect 12178 12484 12182 12540
rect 12182 12484 12238 12540
rect 12238 12484 12242 12540
rect 12178 12480 12242 12484
rect 12258 12540 12322 12544
rect 12258 12484 12262 12540
rect 12262 12484 12318 12540
rect 12318 12484 12322 12540
rect 12258 12480 12322 12484
rect 12338 12540 12402 12544
rect 12338 12484 12342 12540
rect 12342 12484 12398 12540
rect 12398 12484 12402 12540
rect 12338 12480 12402 12484
rect 19872 12540 19936 12544
rect 19872 12484 19876 12540
rect 19876 12484 19932 12540
rect 19932 12484 19936 12540
rect 19872 12480 19936 12484
rect 19952 12540 20016 12544
rect 19952 12484 19956 12540
rect 19956 12484 20012 12540
rect 20012 12484 20016 12540
rect 19952 12480 20016 12484
rect 20032 12540 20096 12544
rect 20032 12484 20036 12540
rect 20036 12484 20092 12540
rect 20092 12484 20096 12540
rect 20032 12480 20096 12484
rect 20112 12540 20176 12544
rect 20112 12484 20116 12540
rect 20116 12484 20172 12540
rect 20172 12484 20176 12540
rect 20112 12480 20176 12484
rect 27646 12540 27710 12544
rect 27646 12484 27650 12540
rect 27650 12484 27706 12540
rect 27706 12484 27710 12540
rect 27646 12480 27710 12484
rect 27726 12540 27790 12544
rect 27726 12484 27730 12540
rect 27730 12484 27786 12540
rect 27786 12484 27790 12540
rect 27726 12480 27790 12484
rect 27806 12540 27870 12544
rect 27806 12484 27810 12540
rect 27810 12484 27866 12540
rect 27866 12484 27870 12540
rect 27806 12480 27870 12484
rect 27886 12540 27950 12544
rect 27886 12484 27890 12540
rect 27890 12484 27946 12540
rect 27946 12484 27950 12540
rect 27886 12480 27950 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 11438 11996 11502 12000
rect 11438 11940 11442 11996
rect 11442 11940 11498 11996
rect 11498 11940 11502 11996
rect 11438 11936 11502 11940
rect 11518 11996 11582 12000
rect 11518 11940 11522 11996
rect 11522 11940 11578 11996
rect 11578 11940 11582 11996
rect 11518 11936 11582 11940
rect 11598 11996 11662 12000
rect 11598 11940 11602 11996
rect 11602 11940 11658 11996
rect 11658 11940 11662 11996
rect 11598 11936 11662 11940
rect 11678 11996 11742 12000
rect 11678 11940 11682 11996
rect 11682 11940 11738 11996
rect 11738 11940 11742 11996
rect 11678 11936 11742 11940
rect 19212 11996 19276 12000
rect 19212 11940 19216 11996
rect 19216 11940 19272 11996
rect 19272 11940 19276 11996
rect 19212 11936 19276 11940
rect 19292 11996 19356 12000
rect 19292 11940 19296 11996
rect 19296 11940 19352 11996
rect 19352 11940 19356 11996
rect 19292 11936 19356 11940
rect 19372 11996 19436 12000
rect 19372 11940 19376 11996
rect 19376 11940 19432 11996
rect 19432 11940 19436 11996
rect 19372 11936 19436 11940
rect 19452 11996 19516 12000
rect 19452 11940 19456 11996
rect 19456 11940 19512 11996
rect 19512 11940 19516 11996
rect 19452 11936 19516 11940
rect 26986 11996 27050 12000
rect 26986 11940 26990 11996
rect 26990 11940 27046 11996
rect 27046 11940 27050 11996
rect 26986 11936 27050 11940
rect 27066 11996 27130 12000
rect 27066 11940 27070 11996
rect 27070 11940 27126 11996
rect 27126 11940 27130 11996
rect 27066 11936 27130 11940
rect 27146 11996 27210 12000
rect 27146 11940 27150 11996
rect 27150 11940 27206 11996
rect 27206 11940 27210 11996
rect 27146 11936 27210 11940
rect 27226 11996 27290 12000
rect 27226 11940 27230 11996
rect 27230 11940 27286 11996
rect 27286 11940 27290 11996
rect 27226 11936 27290 11940
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 12098 11452 12162 11456
rect 12098 11396 12102 11452
rect 12102 11396 12158 11452
rect 12158 11396 12162 11452
rect 12098 11392 12162 11396
rect 12178 11452 12242 11456
rect 12178 11396 12182 11452
rect 12182 11396 12238 11452
rect 12238 11396 12242 11452
rect 12178 11392 12242 11396
rect 12258 11452 12322 11456
rect 12258 11396 12262 11452
rect 12262 11396 12318 11452
rect 12318 11396 12322 11452
rect 12258 11392 12322 11396
rect 12338 11452 12402 11456
rect 12338 11396 12342 11452
rect 12342 11396 12398 11452
rect 12398 11396 12402 11452
rect 12338 11392 12402 11396
rect 19872 11452 19936 11456
rect 19872 11396 19876 11452
rect 19876 11396 19932 11452
rect 19932 11396 19936 11452
rect 19872 11392 19936 11396
rect 19952 11452 20016 11456
rect 19952 11396 19956 11452
rect 19956 11396 20012 11452
rect 20012 11396 20016 11452
rect 19952 11392 20016 11396
rect 20032 11452 20096 11456
rect 20032 11396 20036 11452
rect 20036 11396 20092 11452
rect 20092 11396 20096 11452
rect 20032 11392 20096 11396
rect 20112 11452 20176 11456
rect 20112 11396 20116 11452
rect 20116 11396 20172 11452
rect 20172 11396 20176 11452
rect 20112 11392 20176 11396
rect 27646 11452 27710 11456
rect 27646 11396 27650 11452
rect 27650 11396 27706 11452
rect 27706 11396 27710 11452
rect 27646 11392 27710 11396
rect 27726 11452 27790 11456
rect 27726 11396 27730 11452
rect 27730 11396 27786 11452
rect 27786 11396 27790 11452
rect 27726 11392 27790 11396
rect 27806 11452 27870 11456
rect 27806 11396 27810 11452
rect 27810 11396 27866 11452
rect 27866 11396 27870 11452
rect 27806 11392 27870 11396
rect 27886 11452 27950 11456
rect 27886 11396 27890 11452
rect 27890 11396 27946 11452
rect 27946 11396 27950 11452
rect 27886 11392 27950 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 11438 10908 11502 10912
rect 11438 10852 11442 10908
rect 11442 10852 11498 10908
rect 11498 10852 11502 10908
rect 11438 10848 11502 10852
rect 11518 10908 11582 10912
rect 11518 10852 11522 10908
rect 11522 10852 11578 10908
rect 11578 10852 11582 10908
rect 11518 10848 11582 10852
rect 11598 10908 11662 10912
rect 11598 10852 11602 10908
rect 11602 10852 11658 10908
rect 11658 10852 11662 10908
rect 11598 10848 11662 10852
rect 11678 10908 11742 10912
rect 11678 10852 11682 10908
rect 11682 10852 11738 10908
rect 11738 10852 11742 10908
rect 11678 10848 11742 10852
rect 19212 10908 19276 10912
rect 19212 10852 19216 10908
rect 19216 10852 19272 10908
rect 19272 10852 19276 10908
rect 19212 10848 19276 10852
rect 19292 10908 19356 10912
rect 19292 10852 19296 10908
rect 19296 10852 19352 10908
rect 19352 10852 19356 10908
rect 19292 10848 19356 10852
rect 19372 10908 19436 10912
rect 19372 10852 19376 10908
rect 19376 10852 19432 10908
rect 19432 10852 19436 10908
rect 19372 10848 19436 10852
rect 19452 10908 19516 10912
rect 19452 10852 19456 10908
rect 19456 10852 19512 10908
rect 19512 10852 19516 10908
rect 19452 10848 19516 10852
rect 26986 10908 27050 10912
rect 26986 10852 26990 10908
rect 26990 10852 27046 10908
rect 27046 10852 27050 10908
rect 26986 10848 27050 10852
rect 27066 10908 27130 10912
rect 27066 10852 27070 10908
rect 27070 10852 27126 10908
rect 27126 10852 27130 10908
rect 27066 10848 27130 10852
rect 27146 10908 27210 10912
rect 27146 10852 27150 10908
rect 27150 10852 27206 10908
rect 27206 10852 27210 10908
rect 27146 10848 27210 10852
rect 27226 10908 27290 10912
rect 27226 10852 27230 10908
rect 27230 10852 27286 10908
rect 27286 10852 27290 10908
rect 27226 10848 27290 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 12098 10364 12162 10368
rect 12098 10308 12102 10364
rect 12102 10308 12158 10364
rect 12158 10308 12162 10364
rect 12098 10304 12162 10308
rect 12178 10364 12242 10368
rect 12178 10308 12182 10364
rect 12182 10308 12238 10364
rect 12238 10308 12242 10364
rect 12178 10304 12242 10308
rect 12258 10364 12322 10368
rect 12258 10308 12262 10364
rect 12262 10308 12318 10364
rect 12318 10308 12322 10364
rect 12258 10304 12322 10308
rect 12338 10364 12402 10368
rect 12338 10308 12342 10364
rect 12342 10308 12398 10364
rect 12398 10308 12402 10364
rect 12338 10304 12402 10308
rect 19872 10364 19936 10368
rect 19872 10308 19876 10364
rect 19876 10308 19932 10364
rect 19932 10308 19936 10364
rect 19872 10304 19936 10308
rect 19952 10364 20016 10368
rect 19952 10308 19956 10364
rect 19956 10308 20012 10364
rect 20012 10308 20016 10364
rect 19952 10304 20016 10308
rect 20032 10364 20096 10368
rect 20032 10308 20036 10364
rect 20036 10308 20092 10364
rect 20092 10308 20096 10364
rect 20032 10304 20096 10308
rect 20112 10364 20176 10368
rect 20112 10308 20116 10364
rect 20116 10308 20172 10364
rect 20172 10308 20176 10364
rect 20112 10304 20176 10308
rect 27646 10364 27710 10368
rect 27646 10308 27650 10364
rect 27650 10308 27706 10364
rect 27706 10308 27710 10364
rect 27646 10304 27710 10308
rect 27726 10364 27790 10368
rect 27726 10308 27730 10364
rect 27730 10308 27786 10364
rect 27786 10308 27790 10364
rect 27726 10304 27790 10308
rect 27806 10364 27870 10368
rect 27806 10308 27810 10364
rect 27810 10308 27866 10364
rect 27866 10308 27870 10364
rect 27806 10304 27870 10308
rect 27886 10364 27950 10368
rect 27886 10308 27890 10364
rect 27890 10308 27946 10364
rect 27946 10308 27950 10364
rect 27886 10304 27950 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 11438 9820 11502 9824
rect 11438 9764 11442 9820
rect 11442 9764 11498 9820
rect 11498 9764 11502 9820
rect 11438 9760 11502 9764
rect 11518 9820 11582 9824
rect 11518 9764 11522 9820
rect 11522 9764 11578 9820
rect 11578 9764 11582 9820
rect 11518 9760 11582 9764
rect 11598 9820 11662 9824
rect 11598 9764 11602 9820
rect 11602 9764 11658 9820
rect 11658 9764 11662 9820
rect 11598 9760 11662 9764
rect 11678 9820 11742 9824
rect 11678 9764 11682 9820
rect 11682 9764 11738 9820
rect 11738 9764 11742 9820
rect 11678 9760 11742 9764
rect 19212 9820 19276 9824
rect 19212 9764 19216 9820
rect 19216 9764 19272 9820
rect 19272 9764 19276 9820
rect 19212 9760 19276 9764
rect 19292 9820 19356 9824
rect 19292 9764 19296 9820
rect 19296 9764 19352 9820
rect 19352 9764 19356 9820
rect 19292 9760 19356 9764
rect 19372 9820 19436 9824
rect 19372 9764 19376 9820
rect 19376 9764 19432 9820
rect 19432 9764 19436 9820
rect 19372 9760 19436 9764
rect 19452 9820 19516 9824
rect 19452 9764 19456 9820
rect 19456 9764 19512 9820
rect 19512 9764 19516 9820
rect 19452 9760 19516 9764
rect 26986 9820 27050 9824
rect 26986 9764 26990 9820
rect 26990 9764 27046 9820
rect 27046 9764 27050 9820
rect 26986 9760 27050 9764
rect 27066 9820 27130 9824
rect 27066 9764 27070 9820
rect 27070 9764 27126 9820
rect 27126 9764 27130 9820
rect 27066 9760 27130 9764
rect 27146 9820 27210 9824
rect 27146 9764 27150 9820
rect 27150 9764 27206 9820
rect 27206 9764 27210 9820
rect 27146 9760 27210 9764
rect 27226 9820 27290 9824
rect 27226 9764 27230 9820
rect 27230 9764 27286 9820
rect 27286 9764 27290 9820
rect 27226 9760 27290 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 12098 9276 12162 9280
rect 12098 9220 12102 9276
rect 12102 9220 12158 9276
rect 12158 9220 12162 9276
rect 12098 9216 12162 9220
rect 12178 9276 12242 9280
rect 12178 9220 12182 9276
rect 12182 9220 12238 9276
rect 12238 9220 12242 9276
rect 12178 9216 12242 9220
rect 12258 9276 12322 9280
rect 12258 9220 12262 9276
rect 12262 9220 12318 9276
rect 12318 9220 12322 9276
rect 12258 9216 12322 9220
rect 12338 9276 12402 9280
rect 12338 9220 12342 9276
rect 12342 9220 12398 9276
rect 12398 9220 12402 9276
rect 12338 9216 12402 9220
rect 19872 9276 19936 9280
rect 19872 9220 19876 9276
rect 19876 9220 19932 9276
rect 19932 9220 19936 9276
rect 19872 9216 19936 9220
rect 19952 9276 20016 9280
rect 19952 9220 19956 9276
rect 19956 9220 20012 9276
rect 20012 9220 20016 9276
rect 19952 9216 20016 9220
rect 20032 9276 20096 9280
rect 20032 9220 20036 9276
rect 20036 9220 20092 9276
rect 20092 9220 20096 9276
rect 20032 9216 20096 9220
rect 20112 9276 20176 9280
rect 20112 9220 20116 9276
rect 20116 9220 20172 9276
rect 20172 9220 20176 9276
rect 20112 9216 20176 9220
rect 27646 9276 27710 9280
rect 27646 9220 27650 9276
rect 27650 9220 27706 9276
rect 27706 9220 27710 9276
rect 27646 9216 27710 9220
rect 27726 9276 27790 9280
rect 27726 9220 27730 9276
rect 27730 9220 27786 9276
rect 27786 9220 27790 9276
rect 27726 9216 27790 9220
rect 27806 9276 27870 9280
rect 27806 9220 27810 9276
rect 27810 9220 27866 9276
rect 27866 9220 27870 9276
rect 27806 9216 27870 9220
rect 27886 9276 27950 9280
rect 27886 9220 27890 9276
rect 27890 9220 27946 9276
rect 27946 9220 27950 9276
rect 27886 9216 27950 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 11438 8732 11502 8736
rect 11438 8676 11442 8732
rect 11442 8676 11498 8732
rect 11498 8676 11502 8732
rect 11438 8672 11502 8676
rect 11518 8732 11582 8736
rect 11518 8676 11522 8732
rect 11522 8676 11578 8732
rect 11578 8676 11582 8732
rect 11518 8672 11582 8676
rect 11598 8732 11662 8736
rect 11598 8676 11602 8732
rect 11602 8676 11658 8732
rect 11658 8676 11662 8732
rect 11598 8672 11662 8676
rect 11678 8732 11742 8736
rect 11678 8676 11682 8732
rect 11682 8676 11738 8732
rect 11738 8676 11742 8732
rect 11678 8672 11742 8676
rect 19212 8732 19276 8736
rect 19212 8676 19216 8732
rect 19216 8676 19272 8732
rect 19272 8676 19276 8732
rect 19212 8672 19276 8676
rect 19292 8732 19356 8736
rect 19292 8676 19296 8732
rect 19296 8676 19352 8732
rect 19352 8676 19356 8732
rect 19292 8672 19356 8676
rect 19372 8732 19436 8736
rect 19372 8676 19376 8732
rect 19376 8676 19432 8732
rect 19432 8676 19436 8732
rect 19372 8672 19436 8676
rect 19452 8732 19516 8736
rect 19452 8676 19456 8732
rect 19456 8676 19512 8732
rect 19512 8676 19516 8732
rect 19452 8672 19516 8676
rect 26986 8732 27050 8736
rect 26986 8676 26990 8732
rect 26990 8676 27046 8732
rect 27046 8676 27050 8732
rect 26986 8672 27050 8676
rect 27066 8732 27130 8736
rect 27066 8676 27070 8732
rect 27070 8676 27126 8732
rect 27126 8676 27130 8732
rect 27066 8672 27130 8676
rect 27146 8732 27210 8736
rect 27146 8676 27150 8732
rect 27150 8676 27206 8732
rect 27206 8676 27210 8732
rect 27146 8672 27210 8676
rect 27226 8732 27290 8736
rect 27226 8676 27230 8732
rect 27230 8676 27286 8732
rect 27286 8676 27290 8732
rect 27226 8672 27290 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 12098 8188 12162 8192
rect 12098 8132 12102 8188
rect 12102 8132 12158 8188
rect 12158 8132 12162 8188
rect 12098 8128 12162 8132
rect 12178 8188 12242 8192
rect 12178 8132 12182 8188
rect 12182 8132 12238 8188
rect 12238 8132 12242 8188
rect 12178 8128 12242 8132
rect 12258 8188 12322 8192
rect 12258 8132 12262 8188
rect 12262 8132 12318 8188
rect 12318 8132 12322 8188
rect 12258 8128 12322 8132
rect 12338 8188 12402 8192
rect 12338 8132 12342 8188
rect 12342 8132 12398 8188
rect 12398 8132 12402 8188
rect 12338 8128 12402 8132
rect 19872 8188 19936 8192
rect 19872 8132 19876 8188
rect 19876 8132 19932 8188
rect 19932 8132 19936 8188
rect 19872 8128 19936 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 27646 8188 27710 8192
rect 27646 8132 27650 8188
rect 27650 8132 27706 8188
rect 27706 8132 27710 8188
rect 27646 8128 27710 8132
rect 27726 8188 27790 8192
rect 27726 8132 27730 8188
rect 27730 8132 27786 8188
rect 27786 8132 27790 8188
rect 27726 8128 27790 8132
rect 27806 8188 27870 8192
rect 27806 8132 27810 8188
rect 27810 8132 27866 8188
rect 27866 8132 27870 8188
rect 27806 8128 27870 8132
rect 27886 8188 27950 8192
rect 27886 8132 27890 8188
rect 27890 8132 27946 8188
rect 27946 8132 27950 8188
rect 27886 8128 27950 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 11438 7644 11502 7648
rect 11438 7588 11442 7644
rect 11442 7588 11498 7644
rect 11498 7588 11502 7644
rect 11438 7584 11502 7588
rect 11518 7644 11582 7648
rect 11518 7588 11522 7644
rect 11522 7588 11578 7644
rect 11578 7588 11582 7644
rect 11518 7584 11582 7588
rect 11598 7644 11662 7648
rect 11598 7588 11602 7644
rect 11602 7588 11658 7644
rect 11658 7588 11662 7644
rect 11598 7584 11662 7588
rect 11678 7644 11742 7648
rect 11678 7588 11682 7644
rect 11682 7588 11738 7644
rect 11738 7588 11742 7644
rect 11678 7584 11742 7588
rect 19212 7644 19276 7648
rect 19212 7588 19216 7644
rect 19216 7588 19272 7644
rect 19272 7588 19276 7644
rect 19212 7584 19276 7588
rect 19292 7644 19356 7648
rect 19292 7588 19296 7644
rect 19296 7588 19352 7644
rect 19352 7588 19356 7644
rect 19292 7584 19356 7588
rect 19372 7644 19436 7648
rect 19372 7588 19376 7644
rect 19376 7588 19432 7644
rect 19432 7588 19436 7644
rect 19372 7584 19436 7588
rect 19452 7644 19516 7648
rect 19452 7588 19456 7644
rect 19456 7588 19512 7644
rect 19512 7588 19516 7644
rect 19452 7584 19516 7588
rect 26986 7644 27050 7648
rect 26986 7588 26990 7644
rect 26990 7588 27046 7644
rect 27046 7588 27050 7644
rect 26986 7584 27050 7588
rect 27066 7644 27130 7648
rect 27066 7588 27070 7644
rect 27070 7588 27126 7644
rect 27126 7588 27130 7644
rect 27066 7584 27130 7588
rect 27146 7644 27210 7648
rect 27146 7588 27150 7644
rect 27150 7588 27206 7644
rect 27206 7588 27210 7644
rect 27146 7584 27210 7588
rect 27226 7644 27290 7648
rect 27226 7588 27230 7644
rect 27230 7588 27286 7644
rect 27286 7588 27290 7644
rect 27226 7584 27290 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 12098 7100 12162 7104
rect 12098 7044 12102 7100
rect 12102 7044 12158 7100
rect 12158 7044 12162 7100
rect 12098 7040 12162 7044
rect 12178 7100 12242 7104
rect 12178 7044 12182 7100
rect 12182 7044 12238 7100
rect 12238 7044 12242 7100
rect 12178 7040 12242 7044
rect 12258 7100 12322 7104
rect 12258 7044 12262 7100
rect 12262 7044 12318 7100
rect 12318 7044 12322 7100
rect 12258 7040 12322 7044
rect 12338 7100 12402 7104
rect 12338 7044 12342 7100
rect 12342 7044 12398 7100
rect 12398 7044 12402 7100
rect 12338 7040 12402 7044
rect 19872 7100 19936 7104
rect 19872 7044 19876 7100
rect 19876 7044 19932 7100
rect 19932 7044 19936 7100
rect 19872 7040 19936 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 27646 7100 27710 7104
rect 27646 7044 27650 7100
rect 27650 7044 27706 7100
rect 27706 7044 27710 7100
rect 27646 7040 27710 7044
rect 27726 7100 27790 7104
rect 27726 7044 27730 7100
rect 27730 7044 27786 7100
rect 27786 7044 27790 7100
rect 27726 7040 27790 7044
rect 27806 7100 27870 7104
rect 27806 7044 27810 7100
rect 27810 7044 27866 7100
rect 27866 7044 27870 7100
rect 27806 7040 27870 7044
rect 27886 7100 27950 7104
rect 27886 7044 27890 7100
rect 27890 7044 27946 7100
rect 27946 7044 27950 7100
rect 27886 7040 27950 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 11438 6556 11502 6560
rect 11438 6500 11442 6556
rect 11442 6500 11498 6556
rect 11498 6500 11502 6556
rect 11438 6496 11502 6500
rect 11518 6556 11582 6560
rect 11518 6500 11522 6556
rect 11522 6500 11578 6556
rect 11578 6500 11582 6556
rect 11518 6496 11582 6500
rect 11598 6556 11662 6560
rect 11598 6500 11602 6556
rect 11602 6500 11658 6556
rect 11658 6500 11662 6556
rect 11598 6496 11662 6500
rect 11678 6556 11742 6560
rect 11678 6500 11682 6556
rect 11682 6500 11738 6556
rect 11738 6500 11742 6556
rect 11678 6496 11742 6500
rect 19212 6556 19276 6560
rect 19212 6500 19216 6556
rect 19216 6500 19272 6556
rect 19272 6500 19276 6556
rect 19212 6496 19276 6500
rect 19292 6556 19356 6560
rect 19292 6500 19296 6556
rect 19296 6500 19352 6556
rect 19352 6500 19356 6556
rect 19292 6496 19356 6500
rect 19372 6556 19436 6560
rect 19372 6500 19376 6556
rect 19376 6500 19432 6556
rect 19432 6500 19436 6556
rect 19372 6496 19436 6500
rect 19452 6556 19516 6560
rect 19452 6500 19456 6556
rect 19456 6500 19512 6556
rect 19512 6500 19516 6556
rect 19452 6496 19516 6500
rect 26986 6556 27050 6560
rect 26986 6500 26990 6556
rect 26990 6500 27046 6556
rect 27046 6500 27050 6556
rect 26986 6496 27050 6500
rect 27066 6556 27130 6560
rect 27066 6500 27070 6556
rect 27070 6500 27126 6556
rect 27126 6500 27130 6556
rect 27066 6496 27130 6500
rect 27146 6556 27210 6560
rect 27146 6500 27150 6556
rect 27150 6500 27206 6556
rect 27206 6500 27210 6556
rect 27146 6496 27210 6500
rect 27226 6556 27290 6560
rect 27226 6500 27230 6556
rect 27230 6500 27286 6556
rect 27286 6500 27290 6556
rect 27226 6496 27290 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 12098 6012 12162 6016
rect 12098 5956 12102 6012
rect 12102 5956 12158 6012
rect 12158 5956 12162 6012
rect 12098 5952 12162 5956
rect 12178 6012 12242 6016
rect 12178 5956 12182 6012
rect 12182 5956 12238 6012
rect 12238 5956 12242 6012
rect 12178 5952 12242 5956
rect 12258 6012 12322 6016
rect 12258 5956 12262 6012
rect 12262 5956 12318 6012
rect 12318 5956 12322 6012
rect 12258 5952 12322 5956
rect 12338 6012 12402 6016
rect 12338 5956 12342 6012
rect 12342 5956 12398 6012
rect 12398 5956 12402 6012
rect 12338 5952 12402 5956
rect 19872 6012 19936 6016
rect 19872 5956 19876 6012
rect 19876 5956 19932 6012
rect 19932 5956 19936 6012
rect 19872 5952 19936 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 27646 6012 27710 6016
rect 27646 5956 27650 6012
rect 27650 5956 27706 6012
rect 27706 5956 27710 6012
rect 27646 5952 27710 5956
rect 27726 6012 27790 6016
rect 27726 5956 27730 6012
rect 27730 5956 27786 6012
rect 27786 5956 27790 6012
rect 27726 5952 27790 5956
rect 27806 6012 27870 6016
rect 27806 5956 27810 6012
rect 27810 5956 27866 6012
rect 27866 5956 27870 6012
rect 27806 5952 27870 5956
rect 27886 6012 27950 6016
rect 27886 5956 27890 6012
rect 27890 5956 27946 6012
rect 27946 5956 27950 6012
rect 27886 5952 27950 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 11438 5468 11502 5472
rect 11438 5412 11442 5468
rect 11442 5412 11498 5468
rect 11498 5412 11502 5468
rect 11438 5408 11502 5412
rect 11518 5468 11582 5472
rect 11518 5412 11522 5468
rect 11522 5412 11578 5468
rect 11578 5412 11582 5468
rect 11518 5408 11582 5412
rect 11598 5468 11662 5472
rect 11598 5412 11602 5468
rect 11602 5412 11658 5468
rect 11658 5412 11662 5468
rect 11598 5408 11662 5412
rect 11678 5468 11742 5472
rect 11678 5412 11682 5468
rect 11682 5412 11738 5468
rect 11738 5412 11742 5468
rect 11678 5408 11742 5412
rect 19212 5468 19276 5472
rect 19212 5412 19216 5468
rect 19216 5412 19272 5468
rect 19272 5412 19276 5468
rect 19212 5408 19276 5412
rect 19292 5468 19356 5472
rect 19292 5412 19296 5468
rect 19296 5412 19352 5468
rect 19352 5412 19356 5468
rect 19292 5408 19356 5412
rect 19372 5468 19436 5472
rect 19372 5412 19376 5468
rect 19376 5412 19432 5468
rect 19432 5412 19436 5468
rect 19372 5408 19436 5412
rect 19452 5468 19516 5472
rect 19452 5412 19456 5468
rect 19456 5412 19512 5468
rect 19512 5412 19516 5468
rect 19452 5408 19516 5412
rect 26986 5468 27050 5472
rect 26986 5412 26990 5468
rect 26990 5412 27046 5468
rect 27046 5412 27050 5468
rect 26986 5408 27050 5412
rect 27066 5468 27130 5472
rect 27066 5412 27070 5468
rect 27070 5412 27126 5468
rect 27126 5412 27130 5468
rect 27066 5408 27130 5412
rect 27146 5468 27210 5472
rect 27146 5412 27150 5468
rect 27150 5412 27206 5468
rect 27206 5412 27210 5468
rect 27146 5408 27210 5412
rect 27226 5468 27290 5472
rect 27226 5412 27230 5468
rect 27230 5412 27286 5468
rect 27286 5412 27290 5468
rect 27226 5408 27290 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 12098 4924 12162 4928
rect 12098 4868 12102 4924
rect 12102 4868 12158 4924
rect 12158 4868 12162 4924
rect 12098 4864 12162 4868
rect 12178 4924 12242 4928
rect 12178 4868 12182 4924
rect 12182 4868 12238 4924
rect 12238 4868 12242 4924
rect 12178 4864 12242 4868
rect 12258 4924 12322 4928
rect 12258 4868 12262 4924
rect 12262 4868 12318 4924
rect 12318 4868 12322 4924
rect 12258 4864 12322 4868
rect 12338 4924 12402 4928
rect 12338 4868 12342 4924
rect 12342 4868 12398 4924
rect 12398 4868 12402 4924
rect 12338 4864 12402 4868
rect 19872 4924 19936 4928
rect 19872 4868 19876 4924
rect 19876 4868 19932 4924
rect 19932 4868 19936 4924
rect 19872 4864 19936 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 27646 4924 27710 4928
rect 27646 4868 27650 4924
rect 27650 4868 27706 4924
rect 27706 4868 27710 4924
rect 27646 4864 27710 4868
rect 27726 4924 27790 4928
rect 27726 4868 27730 4924
rect 27730 4868 27786 4924
rect 27786 4868 27790 4924
rect 27726 4864 27790 4868
rect 27806 4924 27870 4928
rect 27806 4868 27810 4924
rect 27810 4868 27866 4924
rect 27866 4868 27870 4924
rect 27806 4864 27870 4868
rect 27886 4924 27950 4928
rect 27886 4868 27890 4924
rect 27890 4868 27946 4924
rect 27946 4868 27950 4924
rect 27886 4864 27950 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 11438 4380 11502 4384
rect 11438 4324 11442 4380
rect 11442 4324 11498 4380
rect 11498 4324 11502 4380
rect 11438 4320 11502 4324
rect 11518 4380 11582 4384
rect 11518 4324 11522 4380
rect 11522 4324 11578 4380
rect 11578 4324 11582 4380
rect 11518 4320 11582 4324
rect 11598 4380 11662 4384
rect 11598 4324 11602 4380
rect 11602 4324 11658 4380
rect 11658 4324 11662 4380
rect 11598 4320 11662 4324
rect 11678 4380 11742 4384
rect 11678 4324 11682 4380
rect 11682 4324 11738 4380
rect 11738 4324 11742 4380
rect 11678 4320 11742 4324
rect 19212 4380 19276 4384
rect 19212 4324 19216 4380
rect 19216 4324 19272 4380
rect 19272 4324 19276 4380
rect 19212 4320 19276 4324
rect 19292 4380 19356 4384
rect 19292 4324 19296 4380
rect 19296 4324 19352 4380
rect 19352 4324 19356 4380
rect 19292 4320 19356 4324
rect 19372 4380 19436 4384
rect 19372 4324 19376 4380
rect 19376 4324 19432 4380
rect 19432 4324 19436 4380
rect 19372 4320 19436 4324
rect 19452 4380 19516 4384
rect 19452 4324 19456 4380
rect 19456 4324 19512 4380
rect 19512 4324 19516 4380
rect 19452 4320 19516 4324
rect 26986 4380 27050 4384
rect 26986 4324 26990 4380
rect 26990 4324 27046 4380
rect 27046 4324 27050 4380
rect 26986 4320 27050 4324
rect 27066 4380 27130 4384
rect 27066 4324 27070 4380
rect 27070 4324 27126 4380
rect 27126 4324 27130 4380
rect 27066 4320 27130 4324
rect 27146 4380 27210 4384
rect 27146 4324 27150 4380
rect 27150 4324 27206 4380
rect 27206 4324 27210 4380
rect 27146 4320 27210 4324
rect 27226 4380 27290 4384
rect 27226 4324 27230 4380
rect 27230 4324 27286 4380
rect 27286 4324 27290 4380
rect 27226 4320 27290 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 12098 3836 12162 3840
rect 12098 3780 12102 3836
rect 12102 3780 12158 3836
rect 12158 3780 12162 3836
rect 12098 3776 12162 3780
rect 12178 3836 12242 3840
rect 12178 3780 12182 3836
rect 12182 3780 12238 3836
rect 12238 3780 12242 3836
rect 12178 3776 12242 3780
rect 12258 3836 12322 3840
rect 12258 3780 12262 3836
rect 12262 3780 12318 3836
rect 12318 3780 12322 3836
rect 12258 3776 12322 3780
rect 12338 3836 12402 3840
rect 12338 3780 12342 3836
rect 12342 3780 12398 3836
rect 12398 3780 12402 3836
rect 12338 3776 12402 3780
rect 19872 3836 19936 3840
rect 19872 3780 19876 3836
rect 19876 3780 19932 3836
rect 19932 3780 19936 3836
rect 19872 3776 19936 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 27646 3836 27710 3840
rect 27646 3780 27650 3836
rect 27650 3780 27706 3836
rect 27706 3780 27710 3836
rect 27646 3776 27710 3780
rect 27726 3836 27790 3840
rect 27726 3780 27730 3836
rect 27730 3780 27786 3836
rect 27786 3780 27790 3836
rect 27726 3776 27790 3780
rect 27806 3836 27870 3840
rect 27806 3780 27810 3836
rect 27810 3780 27866 3836
rect 27866 3780 27870 3836
rect 27806 3776 27870 3780
rect 27886 3836 27950 3840
rect 27886 3780 27890 3836
rect 27890 3780 27946 3836
rect 27946 3780 27950 3836
rect 27886 3776 27950 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 11438 3292 11502 3296
rect 11438 3236 11442 3292
rect 11442 3236 11498 3292
rect 11498 3236 11502 3292
rect 11438 3232 11502 3236
rect 11518 3292 11582 3296
rect 11518 3236 11522 3292
rect 11522 3236 11578 3292
rect 11578 3236 11582 3292
rect 11518 3232 11582 3236
rect 11598 3292 11662 3296
rect 11598 3236 11602 3292
rect 11602 3236 11658 3292
rect 11658 3236 11662 3292
rect 11598 3232 11662 3236
rect 11678 3292 11742 3296
rect 11678 3236 11682 3292
rect 11682 3236 11738 3292
rect 11738 3236 11742 3292
rect 11678 3232 11742 3236
rect 19212 3292 19276 3296
rect 19212 3236 19216 3292
rect 19216 3236 19272 3292
rect 19272 3236 19276 3292
rect 19212 3232 19276 3236
rect 19292 3292 19356 3296
rect 19292 3236 19296 3292
rect 19296 3236 19352 3292
rect 19352 3236 19356 3292
rect 19292 3232 19356 3236
rect 19372 3292 19436 3296
rect 19372 3236 19376 3292
rect 19376 3236 19432 3292
rect 19432 3236 19436 3292
rect 19372 3232 19436 3236
rect 19452 3292 19516 3296
rect 19452 3236 19456 3292
rect 19456 3236 19512 3292
rect 19512 3236 19516 3292
rect 19452 3232 19516 3236
rect 26986 3292 27050 3296
rect 26986 3236 26990 3292
rect 26990 3236 27046 3292
rect 27046 3236 27050 3292
rect 26986 3232 27050 3236
rect 27066 3292 27130 3296
rect 27066 3236 27070 3292
rect 27070 3236 27126 3292
rect 27126 3236 27130 3292
rect 27066 3232 27130 3236
rect 27146 3292 27210 3296
rect 27146 3236 27150 3292
rect 27150 3236 27206 3292
rect 27206 3236 27210 3292
rect 27146 3232 27210 3236
rect 27226 3292 27290 3296
rect 27226 3236 27230 3292
rect 27230 3236 27286 3292
rect 27286 3236 27290 3292
rect 27226 3232 27290 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 12098 2748 12162 2752
rect 12098 2692 12102 2748
rect 12102 2692 12158 2748
rect 12158 2692 12162 2748
rect 12098 2688 12162 2692
rect 12178 2748 12242 2752
rect 12178 2692 12182 2748
rect 12182 2692 12238 2748
rect 12238 2692 12242 2748
rect 12178 2688 12242 2692
rect 12258 2748 12322 2752
rect 12258 2692 12262 2748
rect 12262 2692 12318 2748
rect 12318 2692 12322 2748
rect 12258 2688 12322 2692
rect 12338 2748 12402 2752
rect 12338 2692 12342 2748
rect 12342 2692 12398 2748
rect 12398 2692 12402 2748
rect 12338 2688 12402 2692
rect 19872 2748 19936 2752
rect 19872 2692 19876 2748
rect 19876 2692 19932 2748
rect 19932 2692 19936 2748
rect 19872 2688 19936 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 27646 2748 27710 2752
rect 27646 2692 27650 2748
rect 27650 2692 27706 2748
rect 27706 2692 27710 2748
rect 27646 2688 27710 2692
rect 27726 2748 27790 2752
rect 27726 2692 27730 2748
rect 27730 2692 27786 2748
rect 27786 2692 27790 2748
rect 27726 2688 27790 2692
rect 27806 2748 27870 2752
rect 27806 2692 27810 2748
rect 27810 2692 27866 2748
rect 27866 2692 27870 2748
rect 27806 2688 27870 2692
rect 27886 2748 27950 2752
rect 27886 2692 27890 2748
rect 27890 2692 27946 2748
rect 27946 2692 27950 2748
rect 27886 2688 27950 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 11438 2204 11502 2208
rect 11438 2148 11442 2204
rect 11442 2148 11498 2204
rect 11498 2148 11502 2204
rect 11438 2144 11502 2148
rect 11518 2204 11582 2208
rect 11518 2148 11522 2204
rect 11522 2148 11578 2204
rect 11578 2148 11582 2204
rect 11518 2144 11582 2148
rect 11598 2204 11662 2208
rect 11598 2148 11602 2204
rect 11602 2148 11658 2204
rect 11658 2148 11662 2204
rect 11598 2144 11662 2148
rect 11678 2204 11742 2208
rect 11678 2148 11682 2204
rect 11682 2148 11738 2204
rect 11738 2148 11742 2204
rect 11678 2144 11742 2148
rect 19212 2204 19276 2208
rect 19212 2148 19216 2204
rect 19216 2148 19272 2204
rect 19272 2148 19276 2204
rect 19212 2144 19276 2148
rect 19292 2204 19356 2208
rect 19292 2148 19296 2204
rect 19296 2148 19352 2204
rect 19352 2148 19356 2204
rect 19292 2144 19356 2148
rect 19372 2204 19436 2208
rect 19372 2148 19376 2204
rect 19376 2148 19432 2204
rect 19432 2148 19436 2204
rect 19372 2144 19436 2148
rect 19452 2204 19516 2208
rect 19452 2148 19456 2204
rect 19456 2148 19512 2204
rect 19512 2148 19516 2204
rect 19452 2144 19516 2148
rect 26986 2204 27050 2208
rect 26986 2148 26990 2204
rect 26990 2148 27046 2204
rect 27046 2148 27050 2204
rect 26986 2144 27050 2148
rect 27066 2204 27130 2208
rect 27066 2148 27070 2204
rect 27070 2148 27126 2204
rect 27126 2148 27130 2204
rect 27066 2144 27130 2148
rect 27146 2204 27210 2208
rect 27146 2148 27150 2204
rect 27150 2148 27206 2204
rect 27206 2148 27210 2204
rect 27146 2144 27210 2148
rect 27226 2204 27290 2208
rect 27226 2148 27230 2204
rect 27230 2148 27286 2204
rect 27286 2148 27290 2204
rect 27226 2144 27290 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 12098 1660 12162 1664
rect 12098 1604 12102 1660
rect 12102 1604 12158 1660
rect 12158 1604 12162 1660
rect 12098 1600 12162 1604
rect 12178 1660 12242 1664
rect 12178 1604 12182 1660
rect 12182 1604 12238 1660
rect 12238 1604 12242 1660
rect 12178 1600 12242 1604
rect 12258 1660 12322 1664
rect 12258 1604 12262 1660
rect 12262 1604 12318 1660
rect 12318 1604 12322 1660
rect 12258 1600 12322 1604
rect 12338 1660 12402 1664
rect 12338 1604 12342 1660
rect 12342 1604 12398 1660
rect 12398 1604 12402 1660
rect 12338 1600 12402 1604
rect 19872 1660 19936 1664
rect 19872 1604 19876 1660
rect 19876 1604 19932 1660
rect 19932 1604 19936 1660
rect 19872 1600 19936 1604
rect 19952 1660 20016 1664
rect 19952 1604 19956 1660
rect 19956 1604 20012 1660
rect 20012 1604 20016 1660
rect 19952 1600 20016 1604
rect 20032 1660 20096 1664
rect 20032 1604 20036 1660
rect 20036 1604 20092 1660
rect 20092 1604 20096 1660
rect 20032 1600 20096 1604
rect 20112 1660 20176 1664
rect 20112 1604 20116 1660
rect 20116 1604 20172 1660
rect 20172 1604 20176 1660
rect 20112 1600 20176 1604
rect 27646 1660 27710 1664
rect 27646 1604 27650 1660
rect 27650 1604 27706 1660
rect 27706 1604 27710 1660
rect 27646 1600 27710 1604
rect 27726 1660 27790 1664
rect 27726 1604 27730 1660
rect 27730 1604 27786 1660
rect 27786 1604 27790 1660
rect 27726 1600 27790 1604
rect 27806 1660 27870 1664
rect 27806 1604 27810 1660
rect 27810 1604 27866 1660
rect 27866 1604 27870 1660
rect 27806 1600 27870 1604
rect 27886 1660 27950 1664
rect 27886 1604 27890 1660
rect 27890 1604 27946 1660
rect 27946 1604 27950 1660
rect 27886 1600 27950 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 11438 1116 11502 1120
rect 11438 1060 11442 1116
rect 11442 1060 11498 1116
rect 11498 1060 11502 1116
rect 11438 1056 11502 1060
rect 11518 1116 11582 1120
rect 11518 1060 11522 1116
rect 11522 1060 11578 1116
rect 11578 1060 11582 1116
rect 11518 1056 11582 1060
rect 11598 1116 11662 1120
rect 11598 1060 11602 1116
rect 11602 1060 11658 1116
rect 11658 1060 11662 1116
rect 11598 1056 11662 1060
rect 11678 1116 11742 1120
rect 11678 1060 11682 1116
rect 11682 1060 11738 1116
rect 11738 1060 11742 1116
rect 11678 1056 11742 1060
rect 19212 1116 19276 1120
rect 19212 1060 19216 1116
rect 19216 1060 19272 1116
rect 19272 1060 19276 1116
rect 19212 1056 19276 1060
rect 19292 1116 19356 1120
rect 19292 1060 19296 1116
rect 19296 1060 19352 1116
rect 19352 1060 19356 1116
rect 19292 1056 19356 1060
rect 19372 1116 19436 1120
rect 19372 1060 19376 1116
rect 19376 1060 19432 1116
rect 19432 1060 19436 1116
rect 19372 1056 19436 1060
rect 19452 1116 19516 1120
rect 19452 1060 19456 1116
rect 19456 1060 19512 1116
rect 19512 1060 19516 1116
rect 19452 1056 19516 1060
rect 26986 1116 27050 1120
rect 26986 1060 26990 1116
rect 26990 1060 27046 1116
rect 27046 1060 27050 1116
rect 26986 1056 27050 1060
rect 27066 1116 27130 1120
rect 27066 1060 27070 1116
rect 27070 1060 27126 1116
rect 27126 1060 27130 1116
rect 27066 1056 27130 1060
rect 27146 1116 27210 1120
rect 27146 1060 27150 1116
rect 27150 1060 27206 1116
rect 27206 1060 27210 1116
rect 27146 1056 27210 1060
rect 27226 1116 27290 1120
rect 27226 1060 27230 1116
rect 27230 1060 27286 1116
rect 27286 1060 27290 1116
rect 27226 1056 27290 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 12098 572 12162 576
rect 12098 516 12102 572
rect 12102 516 12158 572
rect 12158 516 12162 572
rect 12098 512 12162 516
rect 12178 572 12242 576
rect 12178 516 12182 572
rect 12182 516 12238 572
rect 12238 516 12242 572
rect 12178 512 12242 516
rect 12258 572 12322 576
rect 12258 516 12262 572
rect 12262 516 12318 572
rect 12318 516 12322 572
rect 12258 512 12322 516
rect 12338 572 12402 576
rect 12338 516 12342 572
rect 12342 516 12398 572
rect 12398 516 12402 572
rect 12338 512 12402 516
rect 19872 572 19936 576
rect 19872 516 19876 572
rect 19876 516 19932 572
rect 19932 516 19936 572
rect 19872 512 19936 516
rect 19952 572 20016 576
rect 19952 516 19956 572
rect 19956 516 20012 572
rect 20012 516 20016 572
rect 19952 512 20016 516
rect 20032 572 20096 576
rect 20032 516 20036 572
rect 20036 516 20092 572
rect 20092 516 20096 572
rect 20032 512 20096 516
rect 20112 572 20176 576
rect 20112 516 20116 572
rect 20116 516 20172 572
rect 20172 516 20176 572
rect 20112 512 20176 516
rect 27646 572 27710 576
rect 27646 516 27650 572
rect 27650 516 27706 572
rect 27706 516 27710 572
rect 27646 512 27710 516
rect 27726 572 27790 576
rect 27726 516 27730 572
rect 27730 516 27786 572
rect 27786 516 27790 572
rect 27726 512 27790 516
rect 27806 572 27870 576
rect 27806 516 27810 572
rect 27810 516 27866 572
rect 27866 516 27870 572
rect 27806 512 27870 516
rect 27886 572 27950 576
rect 27886 516 27890 572
rect 27890 516 27946 572
rect 27946 516 27950 572
rect 27886 512 27950 516
<< metal4 >>
rect 3656 44640 3976 44656
rect 3656 44576 3664 44640
rect 3728 44576 3744 44640
rect 3808 44576 3824 44640
rect 3888 44576 3904 44640
rect 3968 44576 3976 44640
rect 3656 43552 3976 44576
rect 3656 43488 3664 43552
rect 3728 43488 3744 43552
rect 3808 43488 3824 43552
rect 3888 43488 3904 43552
rect 3968 43488 3976 43552
rect 3656 42464 3976 43488
rect 3656 42400 3664 42464
rect 3728 42400 3744 42464
rect 3808 42400 3824 42464
rect 3888 42400 3904 42464
rect 3968 42400 3976 42464
rect 3656 41376 3976 42400
rect 3656 41312 3664 41376
rect 3728 41312 3744 41376
rect 3808 41312 3824 41376
rect 3888 41312 3904 41376
rect 3968 41312 3976 41376
rect 3656 40288 3976 41312
rect 3656 40224 3664 40288
rect 3728 40224 3744 40288
rect 3808 40224 3824 40288
rect 3888 40224 3904 40288
rect 3968 40224 3976 40288
rect 3656 39200 3976 40224
rect 3656 39136 3664 39200
rect 3728 39136 3744 39200
rect 3808 39136 3824 39200
rect 3888 39136 3904 39200
rect 3968 39136 3976 39200
rect 3656 38112 3976 39136
rect 3656 38048 3664 38112
rect 3728 38048 3744 38112
rect 3808 38048 3824 38112
rect 3888 38048 3904 38112
rect 3968 38048 3976 38112
rect 3656 37024 3976 38048
rect 3656 36960 3664 37024
rect 3728 36960 3744 37024
rect 3808 36960 3824 37024
rect 3888 36960 3904 37024
rect 3968 36960 3976 37024
rect 3656 35936 3976 36960
rect 3656 35872 3664 35936
rect 3728 35872 3744 35936
rect 3808 35872 3824 35936
rect 3888 35872 3904 35936
rect 3968 35872 3976 35936
rect 3656 34848 3976 35872
rect 3656 34784 3664 34848
rect 3728 34784 3744 34848
rect 3808 34784 3824 34848
rect 3888 34784 3904 34848
rect 3968 34784 3976 34848
rect 3656 33760 3976 34784
rect 3656 33696 3664 33760
rect 3728 33696 3744 33760
rect 3808 33696 3824 33760
rect 3888 33696 3904 33760
rect 3968 33696 3976 33760
rect 3656 32672 3976 33696
rect 3656 32608 3664 32672
rect 3728 32608 3744 32672
rect 3808 32608 3824 32672
rect 3888 32608 3904 32672
rect 3968 32608 3976 32672
rect 3656 31584 3976 32608
rect 3656 31520 3664 31584
rect 3728 31520 3744 31584
rect 3808 31520 3824 31584
rect 3888 31520 3904 31584
rect 3968 31520 3976 31584
rect 3656 30496 3976 31520
rect 3656 30432 3664 30496
rect 3728 30432 3744 30496
rect 3808 30432 3824 30496
rect 3888 30432 3904 30496
rect 3968 30432 3976 30496
rect 3656 29408 3976 30432
rect 3656 29344 3664 29408
rect 3728 29344 3744 29408
rect 3808 29344 3824 29408
rect 3888 29344 3904 29408
rect 3968 29344 3976 29408
rect 3656 28320 3976 29344
rect 3656 28256 3664 28320
rect 3728 28256 3744 28320
rect 3808 28256 3824 28320
rect 3888 28256 3904 28320
rect 3968 28256 3976 28320
rect 3656 27232 3976 28256
rect 3656 27168 3664 27232
rect 3728 27168 3744 27232
rect 3808 27168 3824 27232
rect 3888 27168 3904 27232
rect 3968 27168 3976 27232
rect 3656 26144 3976 27168
rect 3656 26080 3664 26144
rect 3728 26080 3744 26144
rect 3808 26080 3824 26144
rect 3888 26080 3904 26144
rect 3968 26080 3976 26144
rect 3656 25056 3976 26080
rect 3656 24992 3664 25056
rect 3728 24992 3744 25056
rect 3808 24992 3824 25056
rect 3888 24992 3904 25056
rect 3968 24992 3976 25056
rect 3656 23968 3976 24992
rect 3656 23904 3664 23968
rect 3728 23904 3744 23968
rect 3808 23904 3824 23968
rect 3888 23904 3904 23968
rect 3968 23904 3976 23968
rect 3656 22880 3976 23904
rect 3656 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3976 22880
rect 3656 21792 3976 22816
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 44096 4636 44656
rect 4316 44032 4324 44096
rect 4388 44032 4404 44096
rect 4468 44032 4484 44096
rect 4548 44032 4564 44096
rect 4628 44032 4636 44096
rect 4316 43008 4636 44032
rect 6134 44029 6194 45152
rect 6686 44029 6746 45152
rect 7238 44573 7298 45152
rect 7790 44573 7850 45152
rect 8342 44573 8402 45152
rect 8894 44573 8954 45152
rect 9446 44573 9506 45152
rect 7235 44572 7301 44573
rect 7235 44508 7236 44572
rect 7300 44508 7301 44572
rect 7235 44507 7301 44508
rect 7787 44572 7853 44573
rect 7787 44508 7788 44572
rect 7852 44508 7853 44572
rect 7787 44507 7853 44508
rect 8339 44572 8405 44573
rect 8339 44508 8340 44572
rect 8404 44508 8405 44572
rect 8339 44507 8405 44508
rect 8891 44572 8957 44573
rect 8891 44508 8892 44572
rect 8956 44508 8957 44572
rect 8891 44507 8957 44508
rect 9443 44572 9509 44573
rect 9443 44508 9444 44572
rect 9508 44508 9509 44572
rect 9443 44507 9509 44508
rect 9998 44029 10058 45152
rect 6131 44028 6197 44029
rect 6131 43964 6132 44028
rect 6196 43964 6197 44028
rect 6131 43963 6197 43964
rect 6683 44028 6749 44029
rect 6683 43964 6684 44028
rect 6748 43964 6749 44028
rect 6683 43963 6749 43964
rect 9995 44028 10061 44029
rect 9995 43964 9996 44028
rect 10060 43964 10061 44028
rect 9995 43963 10061 43964
rect 4316 42944 4324 43008
rect 4388 42944 4404 43008
rect 4468 42944 4484 43008
rect 4548 42944 4564 43008
rect 4628 42944 4636 43008
rect 4316 41920 4636 42944
rect 4316 41856 4324 41920
rect 4388 41856 4404 41920
rect 4468 41856 4484 41920
rect 4548 41856 4564 41920
rect 4628 41856 4636 41920
rect 4316 40832 4636 41856
rect 4316 40768 4324 40832
rect 4388 40768 4404 40832
rect 4468 40768 4484 40832
rect 4548 40768 4564 40832
rect 4628 40768 4636 40832
rect 4316 39744 4636 40768
rect 4316 39680 4324 39744
rect 4388 39680 4404 39744
rect 4468 39680 4484 39744
rect 4548 39680 4564 39744
rect 4628 39680 4636 39744
rect 4316 38656 4636 39680
rect 4316 38592 4324 38656
rect 4388 38592 4404 38656
rect 4468 38592 4484 38656
rect 4548 38592 4564 38656
rect 4628 38592 4636 38656
rect 4316 37568 4636 38592
rect 4316 37504 4324 37568
rect 4388 37504 4404 37568
rect 4468 37504 4484 37568
rect 4548 37504 4564 37568
rect 4628 37504 4636 37568
rect 4316 36480 4636 37504
rect 4316 36416 4324 36480
rect 4388 36416 4404 36480
rect 4468 36416 4484 36480
rect 4548 36416 4564 36480
rect 4628 36416 4636 36480
rect 4316 35392 4636 36416
rect 10550 36141 10610 45152
rect 11102 43893 11162 45152
rect 11654 44845 11714 45152
rect 12206 44845 12266 45152
rect 11651 44844 11717 44845
rect 11651 44780 11652 44844
rect 11716 44780 11717 44844
rect 11651 44779 11717 44780
rect 12203 44844 12269 44845
rect 12203 44780 12204 44844
rect 12268 44780 12269 44844
rect 12203 44779 12269 44780
rect 11430 44640 11750 44656
rect 11430 44576 11438 44640
rect 11502 44576 11518 44640
rect 11582 44576 11598 44640
rect 11662 44576 11678 44640
rect 11742 44576 11750 44640
rect 11099 43892 11165 43893
rect 11099 43828 11100 43892
rect 11164 43828 11165 43892
rect 11099 43827 11165 43828
rect 11430 43552 11750 44576
rect 11430 43488 11438 43552
rect 11502 43488 11518 43552
rect 11582 43488 11598 43552
rect 11662 43488 11678 43552
rect 11742 43488 11750 43552
rect 11430 42464 11750 43488
rect 11430 42400 11438 42464
rect 11502 42400 11518 42464
rect 11582 42400 11598 42464
rect 11662 42400 11678 42464
rect 11742 42400 11750 42464
rect 11430 41376 11750 42400
rect 11430 41312 11438 41376
rect 11502 41312 11518 41376
rect 11582 41312 11598 41376
rect 11662 41312 11678 41376
rect 11742 41312 11750 41376
rect 11430 40288 11750 41312
rect 11430 40224 11438 40288
rect 11502 40224 11518 40288
rect 11582 40224 11598 40288
rect 11662 40224 11678 40288
rect 11742 40224 11750 40288
rect 11430 39200 11750 40224
rect 11430 39136 11438 39200
rect 11502 39136 11518 39200
rect 11582 39136 11598 39200
rect 11662 39136 11678 39200
rect 11742 39136 11750 39200
rect 11430 38112 11750 39136
rect 11430 38048 11438 38112
rect 11502 38048 11518 38112
rect 11582 38048 11598 38112
rect 11662 38048 11678 38112
rect 11742 38048 11750 38112
rect 11430 37024 11750 38048
rect 11430 36960 11438 37024
rect 11502 36960 11518 37024
rect 11582 36960 11598 37024
rect 11662 36960 11678 37024
rect 11742 36960 11750 37024
rect 10547 36140 10613 36141
rect 10547 36076 10548 36140
rect 10612 36076 10613 36140
rect 10547 36075 10613 36076
rect 4316 35328 4324 35392
rect 4388 35328 4404 35392
rect 4468 35328 4484 35392
rect 4548 35328 4564 35392
rect 4628 35328 4636 35392
rect 4316 34304 4636 35328
rect 4316 34240 4324 34304
rect 4388 34240 4404 34304
rect 4468 34240 4484 34304
rect 4548 34240 4564 34304
rect 4628 34240 4636 34304
rect 4316 33216 4636 34240
rect 4316 33152 4324 33216
rect 4388 33152 4404 33216
rect 4468 33152 4484 33216
rect 4548 33152 4564 33216
rect 4628 33152 4636 33216
rect 4316 32128 4636 33152
rect 4316 32064 4324 32128
rect 4388 32064 4404 32128
rect 4468 32064 4484 32128
rect 4548 32064 4564 32128
rect 4628 32064 4636 32128
rect 4316 31040 4636 32064
rect 4316 30976 4324 31040
rect 4388 30976 4404 31040
rect 4468 30976 4484 31040
rect 4548 30976 4564 31040
rect 4628 30976 4636 31040
rect 4316 29952 4636 30976
rect 4316 29888 4324 29952
rect 4388 29888 4404 29952
rect 4468 29888 4484 29952
rect 4548 29888 4564 29952
rect 4628 29888 4636 29952
rect 4316 28864 4636 29888
rect 4316 28800 4324 28864
rect 4388 28800 4404 28864
rect 4468 28800 4484 28864
rect 4548 28800 4564 28864
rect 4628 28800 4636 28864
rect 4316 27776 4636 28800
rect 4316 27712 4324 27776
rect 4388 27712 4404 27776
rect 4468 27712 4484 27776
rect 4548 27712 4564 27776
rect 4628 27712 4636 27776
rect 4316 26688 4636 27712
rect 4316 26624 4324 26688
rect 4388 26624 4404 26688
rect 4468 26624 4484 26688
rect 4548 26624 4564 26688
rect 4628 26624 4636 26688
rect 4316 25600 4636 26624
rect 4316 25536 4324 25600
rect 4388 25536 4404 25600
rect 4468 25536 4484 25600
rect 4548 25536 4564 25600
rect 4628 25536 4636 25600
rect 4316 24512 4636 25536
rect 4316 24448 4324 24512
rect 4388 24448 4404 24512
rect 4468 24448 4484 24512
rect 4548 24448 4564 24512
rect 4628 24448 4636 24512
rect 4316 23424 4636 24448
rect 4316 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4636 23424
rect 4316 22336 4636 23360
rect 4316 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4636 22336
rect 4316 21248 4636 22272
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 11430 35936 11750 36960
rect 11430 35872 11438 35936
rect 11502 35872 11518 35936
rect 11582 35872 11598 35936
rect 11662 35872 11678 35936
rect 11742 35872 11750 35936
rect 11430 34848 11750 35872
rect 11430 34784 11438 34848
rect 11502 34784 11518 34848
rect 11582 34784 11598 34848
rect 11662 34784 11678 34848
rect 11742 34784 11750 34848
rect 11430 33760 11750 34784
rect 11430 33696 11438 33760
rect 11502 33696 11518 33760
rect 11582 33696 11598 33760
rect 11662 33696 11678 33760
rect 11742 33696 11750 33760
rect 11430 32672 11750 33696
rect 11430 32608 11438 32672
rect 11502 32608 11518 32672
rect 11582 32608 11598 32672
rect 11662 32608 11678 32672
rect 11742 32608 11750 32672
rect 11430 31584 11750 32608
rect 11430 31520 11438 31584
rect 11502 31520 11518 31584
rect 11582 31520 11598 31584
rect 11662 31520 11678 31584
rect 11742 31520 11750 31584
rect 11430 30496 11750 31520
rect 11430 30432 11438 30496
rect 11502 30432 11518 30496
rect 11582 30432 11598 30496
rect 11662 30432 11678 30496
rect 11742 30432 11750 30496
rect 11430 29408 11750 30432
rect 11430 29344 11438 29408
rect 11502 29344 11518 29408
rect 11582 29344 11598 29408
rect 11662 29344 11678 29408
rect 11742 29344 11750 29408
rect 11430 28320 11750 29344
rect 11430 28256 11438 28320
rect 11502 28256 11518 28320
rect 11582 28256 11598 28320
rect 11662 28256 11678 28320
rect 11742 28256 11750 28320
rect 11430 27232 11750 28256
rect 11430 27168 11438 27232
rect 11502 27168 11518 27232
rect 11582 27168 11598 27232
rect 11662 27168 11678 27232
rect 11742 27168 11750 27232
rect 11430 26144 11750 27168
rect 11430 26080 11438 26144
rect 11502 26080 11518 26144
rect 11582 26080 11598 26144
rect 11662 26080 11678 26144
rect 11742 26080 11750 26144
rect 11430 25056 11750 26080
rect 11430 24992 11438 25056
rect 11502 24992 11518 25056
rect 11582 24992 11598 25056
rect 11662 24992 11678 25056
rect 11742 24992 11750 25056
rect 11430 23968 11750 24992
rect 11430 23904 11438 23968
rect 11502 23904 11518 23968
rect 11582 23904 11598 23968
rect 11662 23904 11678 23968
rect 11742 23904 11750 23968
rect 11430 22880 11750 23904
rect 11430 22816 11438 22880
rect 11502 22816 11518 22880
rect 11582 22816 11598 22880
rect 11662 22816 11678 22880
rect 11742 22816 11750 22880
rect 11430 21792 11750 22816
rect 11430 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11750 21792
rect 11430 20704 11750 21728
rect 11430 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11750 20704
rect 11430 19616 11750 20640
rect 11430 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11750 19616
rect 11430 18528 11750 19552
rect 11430 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11750 18528
rect 11430 17440 11750 18464
rect 11430 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11750 17440
rect 11430 16352 11750 17376
rect 11430 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11750 16352
rect 11430 15264 11750 16288
rect 11430 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11750 15264
rect 11430 14176 11750 15200
rect 11430 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11750 14176
rect 11430 13088 11750 14112
rect 11430 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11750 13088
rect 11430 12000 11750 13024
rect 11430 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11750 12000
rect 11430 10912 11750 11936
rect 11430 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11750 10912
rect 11430 9824 11750 10848
rect 11430 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11750 9824
rect 11430 8736 11750 9760
rect 11430 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11750 8736
rect 11430 7648 11750 8672
rect 11430 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11750 7648
rect 11430 6560 11750 7584
rect 11430 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11750 6560
rect 11430 5472 11750 6496
rect 11430 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11750 5472
rect 11430 4384 11750 5408
rect 11430 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11750 4384
rect 11430 3296 11750 4320
rect 11430 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11750 3296
rect 11430 2208 11750 3232
rect 11430 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11750 2208
rect 11430 1120 11750 2144
rect 11430 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11750 1120
rect 11430 496 11750 1056
rect 12090 44096 12410 44656
rect 12758 44573 12818 45152
rect 12755 44572 12821 44573
rect 12755 44508 12756 44572
rect 12820 44508 12821 44572
rect 12755 44507 12821 44508
rect 12090 44032 12098 44096
rect 12162 44032 12178 44096
rect 12242 44032 12258 44096
rect 12322 44032 12338 44096
rect 12402 44032 12410 44096
rect 12090 43008 12410 44032
rect 13310 44029 13370 45152
rect 13307 44028 13373 44029
rect 13307 43964 13308 44028
rect 13372 43964 13373 44028
rect 13307 43963 13373 43964
rect 13862 43757 13922 45152
rect 13859 43756 13925 43757
rect 13859 43692 13860 43756
rect 13924 43692 13925 43756
rect 13859 43691 13925 43692
rect 14414 43485 14474 45152
rect 14411 43484 14477 43485
rect 14411 43420 14412 43484
rect 14476 43420 14477 43484
rect 14411 43419 14477 43420
rect 14966 43213 15026 45152
rect 14963 43212 15029 43213
rect 14963 43148 14964 43212
rect 15028 43148 15029 43212
rect 14963 43147 15029 43148
rect 12090 42944 12098 43008
rect 12162 42944 12178 43008
rect 12242 42944 12258 43008
rect 12322 42944 12338 43008
rect 12402 42944 12410 43008
rect 12090 41920 12410 42944
rect 15518 42941 15578 45152
rect 15515 42940 15581 42941
rect 15515 42876 15516 42940
rect 15580 42876 15581 42940
rect 15515 42875 15581 42876
rect 12090 41856 12098 41920
rect 12162 41856 12178 41920
rect 12242 41856 12258 41920
rect 12322 41856 12338 41920
rect 12402 41856 12410 41920
rect 12090 40832 12410 41856
rect 13675 41852 13741 41853
rect 13675 41788 13676 41852
rect 13740 41788 13741 41852
rect 13675 41787 13741 41788
rect 12090 40768 12098 40832
rect 12162 40768 12178 40832
rect 12242 40768 12258 40832
rect 12322 40768 12338 40832
rect 12402 40768 12410 40832
rect 12090 39744 12410 40768
rect 12090 39680 12098 39744
rect 12162 39680 12178 39744
rect 12242 39680 12258 39744
rect 12322 39680 12338 39744
rect 12402 39680 12410 39744
rect 12090 38656 12410 39680
rect 12090 38592 12098 38656
rect 12162 38592 12178 38656
rect 12242 38592 12258 38656
rect 12322 38592 12338 38656
rect 12402 38592 12410 38656
rect 12090 37568 12410 38592
rect 12090 37504 12098 37568
rect 12162 37504 12178 37568
rect 12242 37504 12258 37568
rect 12322 37504 12338 37568
rect 12402 37504 12410 37568
rect 12090 36480 12410 37504
rect 12090 36416 12098 36480
rect 12162 36416 12178 36480
rect 12242 36416 12258 36480
rect 12322 36416 12338 36480
rect 12402 36416 12410 36480
rect 12090 35392 12410 36416
rect 12090 35328 12098 35392
rect 12162 35328 12178 35392
rect 12242 35328 12258 35392
rect 12322 35328 12338 35392
rect 12402 35328 12410 35392
rect 12090 34304 12410 35328
rect 12090 34240 12098 34304
rect 12162 34240 12178 34304
rect 12242 34240 12258 34304
rect 12322 34240 12338 34304
rect 12402 34240 12410 34304
rect 12090 33216 12410 34240
rect 12090 33152 12098 33216
rect 12162 33152 12178 33216
rect 12242 33152 12258 33216
rect 12322 33152 12338 33216
rect 12402 33152 12410 33216
rect 12090 32128 12410 33152
rect 12090 32064 12098 32128
rect 12162 32064 12178 32128
rect 12242 32064 12258 32128
rect 12322 32064 12338 32128
rect 12402 32064 12410 32128
rect 12090 31040 12410 32064
rect 12090 30976 12098 31040
rect 12162 30976 12178 31040
rect 12242 30976 12258 31040
rect 12322 30976 12338 31040
rect 12402 30976 12410 31040
rect 12090 29952 12410 30976
rect 12090 29888 12098 29952
rect 12162 29888 12178 29952
rect 12242 29888 12258 29952
rect 12322 29888 12338 29952
rect 12402 29888 12410 29952
rect 12090 28864 12410 29888
rect 12090 28800 12098 28864
rect 12162 28800 12178 28864
rect 12242 28800 12258 28864
rect 12322 28800 12338 28864
rect 12402 28800 12410 28864
rect 12090 27776 12410 28800
rect 13678 28797 13738 41787
rect 16070 41173 16130 45152
rect 16622 44029 16682 45152
rect 17174 44029 17234 45152
rect 16619 44028 16685 44029
rect 16619 43964 16620 44028
rect 16684 43964 16685 44028
rect 16619 43963 16685 43964
rect 17171 44028 17237 44029
rect 17171 43964 17172 44028
rect 17236 43964 17237 44028
rect 17171 43963 17237 43964
rect 17726 42941 17786 45152
rect 18278 43213 18338 45152
rect 18830 43349 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44845 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 21587 44844 21653 44845
rect 21587 44780 21588 44844
rect 21652 44780 21653 44844
rect 21587 44779 21653 44780
rect 23798 44709 23858 45152
rect 24350 44709 24410 45152
rect 24902 44709 24962 45152
rect 25454 44709 25514 45152
rect 26006 44709 26066 45152
rect 26558 44709 26618 45152
rect 27110 44845 27170 45152
rect 27662 44845 27722 45152
rect 27107 44844 27173 44845
rect 27107 44780 27108 44844
rect 27172 44780 27173 44844
rect 27107 44779 27173 44780
rect 27659 44844 27725 44845
rect 27659 44780 27660 44844
rect 27724 44780 27725 44844
rect 27659 44779 27725 44780
rect 28214 44709 28274 45152
rect 23795 44708 23861 44709
rect 19204 44640 19524 44656
rect 19204 44576 19212 44640
rect 19276 44576 19292 44640
rect 19356 44576 19372 44640
rect 19436 44576 19452 44640
rect 19516 44576 19524 44640
rect 19204 43552 19524 44576
rect 19204 43488 19212 43552
rect 19276 43488 19292 43552
rect 19356 43488 19372 43552
rect 19436 43488 19452 43552
rect 19516 43488 19524 43552
rect 18827 43348 18893 43349
rect 18827 43284 18828 43348
rect 18892 43284 18893 43348
rect 18827 43283 18893 43284
rect 18275 43212 18341 43213
rect 18275 43148 18276 43212
rect 18340 43148 18341 43212
rect 18275 43147 18341 43148
rect 17723 42940 17789 42941
rect 17723 42876 17724 42940
rect 17788 42876 17789 42940
rect 17723 42875 17789 42876
rect 19204 42464 19524 43488
rect 19204 42400 19212 42464
rect 19276 42400 19292 42464
rect 19356 42400 19372 42464
rect 19436 42400 19452 42464
rect 19516 42400 19524 42464
rect 19204 41376 19524 42400
rect 19204 41312 19212 41376
rect 19276 41312 19292 41376
rect 19356 41312 19372 41376
rect 19436 41312 19452 41376
rect 19516 41312 19524 41376
rect 16067 41172 16133 41173
rect 16067 41108 16068 41172
rect 16132 41108 16133 41172
rect 16067 41107 16133 41108
rect 19204 40288 19524 41312
rect 19204 40224 19212 40288
rect 19276 40224 19292 40288
rect 19356 40224 19372 40288
rect 19436 40224 19452 40288
rect 19516 40224 19524 40288
rect 19204 39200 19524 40224
rect 19204 39136 19212 39200
rect 19276 39136 19292 39200
rect 19356 39136 19372 39200
rect 19436 39136 19452 39200
rect 19516 39136 19524 39200
rect 19204 38112 19524 39136
rect 19204 38048 19212 38112
rect 19276 38048 19292 38112
rect 19356 38048 19372 38112
rect 19436 38048 19452 38112
rect 19516 38048 19524 38112
rect 19204 37024 19524 38048
rect 19204 36960 19212 37024
rect 19276 36960 19292 37024
rect 19356 36960 19372 37024
rect 19436 36960 19452 37024
rect 19516 36960 19524 37024
rect 18459 36004 18525 36005
rect 18459 35940 18460 36004
rect 18524 35940 18525 36004
rect 18459 35939 18525 35940
rect 18462 34101 18522 35939
rect 19204 35936 19524 36960
rect 19204 35872 19212 35936
rect 19276 35872 19292 35936
rect 19356 35872 19372 35936
rect 19436 35872 19452 35936
rect 19516 35872 19524 35936
rect 19204 34848 19524 35872
rect 19204 34784 19212 34848
rect 19276 34784 19292 34848
rect 19356 34784 19372 34848
rect 19436 34784 19452 34848
rect 19516 34784 19524 34848
rect 18459 34100 18525 34101
rect 18459 34036 18460 34100
rect 18524 34036 18525 34100
rect 18459 34035 18525 34036
rect 19204 33760 19524 34784
rect 19204 33696 19212 33760
rect 19276 33696 19292 33760
rect 19356 33696 19372 33760
rect 19436 33696 19452 33760
rect 19516 33696 19524 33760
rect 19204 32672 19524 33696
rect 19204 32608 19212 32672
rect 19276 32608 19292 32672
rect 19356 32608 19372 32672
rect 19436 32608 19452 32672
rect 19516 32608 19524 32672
rect 16987 31924 17053 31925
rect 16987 31860 16988 31924
rect 17052 31860 17053 31924
rect 16987 31859 17053 31860
rect 13675 28796 13741 28797
rect 13675 28732 13676 28796
rect 13740 28732 13741 28796
rect 13675 28731 13741 28732
rect 12090 27712 12098 27776
rect 12162 27712 12178 27776
rect 12242 27712 12258 27776
rect 12322 27712 12338 27776
rect 12402 27712 12410 27776
rect 12090 26688 12410 27712
rect 12090 26624 12098 26688
rect 12162 26624 12178 26688
rect 12242 26624 12258 26688
rect 12322 26624 12338 26688
rect 12402 26624 12410 26688
rect 12090 25600 12410 26624
rect 12090 25536 12098 25600
rect 12162 25536 12178 25600
rect 12242 25536 12258 25600
rect 12322 25536 12338 25600
rect 12402 25536 12410 25600
rect 12090 24512 12410 25536
rect 12090 24448 12098 24512
rect 12162 24448 12178 24512
rect 12242 24448 12258 24512
rect 12322 24448 12338 24512
rect 12402 24448 12410 24512
rect 12090 23424 12410 24448
rect 12090 23360 12098 23424
rect 12162 23360 12178 23424
rect 12242 23360 12258 23424
rect 12322 23360 12338 23424
rect 12402 23360 12410 23424
rect 12090 22336 12410 23360
rect 12090 22272 12098 22336
rect 12162 22272 12178 22336
rect 12242 22272 12258 22336
rect 12322 22272 12338 22336
rect 12402 22272 12410 22336
rect 12090 21248 12410 22272
rect 12090 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12410 21248
rect 12090 20160 12410 21184
rect 12090 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12410 20160
rect 12090 19072 12410 20096
rect 12090 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12410 19072
rect 12090 17984 12410 19008
rect 12090 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12410 17984
rect 12090 16896 12410 17920
rect 12090 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12410 16896
rect 12090 15808 12410 16832
rect 12090 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12410 15808
rect 12090 14720 12410 15744
rect 16990 15197 17050 31859
rect 19204 31584 19524 32608
rect 19204 31520 19212 31584
rect 19276 31520 19292 31584
rect 19356 31520 19372 31584
rect 19436 31520 19452 31584
rect 19516 31520 19524 31584
rect 19204 30496 19524 31520
rect 19204 30432 19212 30496
rect 19276 30432 19292 30496
rect 19356 30432 19372 30496
rect 19436 30432 19452 30496
rect 19516 30432 19524 30496
rect 19204 29408 19524 30432
rect 19204 29344 19212 29408
rect 19276 29344 19292 29408
rect 19356 29344 19372 29408
rect 19436 29344 19452 29408
rect 19516 29344 19524 29408
rect 19204 28320 19524 29344
rect 19204 28256 19212 28320
rect 19276 28256 19292 28320
rect 19356 28256 19372 28320
rect 19436 28256 19452 28320
rect 19516 28256 19524 28320
rect 19204 27232 19524 28256
rect 19204 27168 19212 27232
rect 19276 27168 19292 27232
rect 19356 27168 19372 27232
rect 19436 27168 19452 27232
rect 19516 27168 19524 27232
rect 19204 26144 19524 27168
rect 19204 26080 19212 26144
rect 19276 26080 19292 26144
rect 19356 26080 19372 26144
rect 19436 26080 19452 26144
rect 19516 26080 19524 26144
rect 19204 25056 19524 26080
rect 19204 24992 19212 25056
rect 19276 24992 19292 25056
rect 19356 24992 19372 25056
rect 19436 24992 19452 25056
rect 19516 24992 19524 25056
rect 19204 23968 19524 24992
rect 19204 23904 19212 23968
rect 19276 23904 19292 23968
rect 19356 23904 19372 23968
rect 19436 23904 19452 23968
rect 19516 23904 19524 23968
rect 19204 22880 19524 23904
rect 19204 22816 19212 22880
rect 19276 22816 19292 22880
rect 19356 22816 19372 22880
rect 19436 22816 19452 22880
rect 19516 22816 19524 22880
rect 19204 21792 19524 22816
rect 19204 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19524 21792
rect 19204 20704 19524 21728
rect 19204 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19524 20704
rect 19204 19616 19524 20640
rect 19204 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19524 19616
rect 19204 18528 19524 19552
rect 19204 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19524 18528
rect 19204 17440 19524 18464
rect 19204 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19524 17440
rect 19204 16352 19524 17376
rect 19204 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19524 16352
rect 19204 15264 19524 16288
rect 19204 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19524 15264
rect 16987 15196 17053 15197
rect 16987 15132 16988 15196
rect 17052 15132 17053 15196
rect 16987 15131 17053 15132
rect 12090 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12410 14720
rect 12090 13632 12410 14656
rect 12090 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12410 13632
rect 12090 12544 12410 13568
rect 12090 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12410 12544
rect 12090 11456 12410 12480
rect 12090 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12410 11456
rect 12090 10368 12410 11392
rect 12090 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12410 10368
rect 12090 9280 12410 10304
rect 12090 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12410 9280
rect 12090 8192 12410 9216
rect 12090 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12410 8192
rect 12090 7104 12410 8128
rect 12090 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12410 7104
rect 12090 6016 12410 7040
rect 12090 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12410 6016
rect 12090 4928 12410 5952
rect 12090 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12410 4928
rect 12090 3840 12410 4864
rect 12090 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12410 3840
rect 12090 2752 12410 3776
rect 12090 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12410 2752
rect 12090 1664 12410 2688
rect 12090 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12410 1664
rect 12090 576 12410 1600
rect 12090 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12410 576
rect 12090 496 12410 512
rect 19204 14176 19524 15200
rect 19204 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19524 14176
rect 19204 13088 19524 14112
rect 19204 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19524 13088
rect 19204 12000 19524 13024
rect 19204 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19524 12000
rect 19204 10912 19524 11936
rect 19204 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19524 10912
rect 19204 9824 19524 10848
rect 19204 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19524 9824
rect 19204 8736 19524 9760
rect 19204 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19524 8736
rect 19204 7648 19524 8672
rect 19204 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19524 7648
rect 19204 6560 19524 7584
rect 19204 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19524 6560
rect 19204 5472 19524 6496
rect 19204 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19524 5472
rect 19204 4384 19524 5408
rect 19204 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19524 4384
rect 19204 3296 19524 4320
rect 19204 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19524 3296
rect 19204 2208 19524 3232
rect 19204 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19524 2208
rect 19204 1120 19524 2144
rect 19204 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19524 1120
rect 19204 496 19524 1056
rect 19864 44096 20184 44656
rect 23795 44644 23796 44708
rect 23860 44644 23861 44708
rect 23795 44643 23861 44644
rect 24347 44708 24413 44709
rect 24347 44644 24348 44708
rect 24412 44644 24413 44708
rect 24347 44643 24413 44644
rect 24899 44708 24965 44709
rect 24899 44644 24900 44708
rect 24964 44644 24965 44708
rect 24899 44643 24965 44644
rect 25451 44708 25517 44709
rect 25451 44644 25452 44708
rect 25516 44644 25517 44708
rect 25451 44643 25517 44644
rect 26003 44708 26069 44709
rect 26003 44644 26004 44708
rect 26068 44644 26069 44708
rect 26003 44643 26069 44644
rect 26555 44708 26621 44709
rect 26555 44644 26556 44708
rect 26620 44644 26621 44708
rect 28211 44708 28277 44709
rect 26555 44643 26621 44644
rect 19864 44032 19872 44096
rect 19936 44032 19952 44096
rect 20016 44032 20032 44096
rect 20096 44032 20112 44096
rect 20176 44032 20184 44096
rect 19864 43008 20184 44032
rect 19864 42944 19872 43008
rect 19936 42944 19952 43008
rect 20016 42944 20032 43008
rect 20096 42944 20112 43008
rect 20176 42944 20184 43008
rect 19864 41920 20184 42944
rect 26978 44640 27298 44656
rect 26978 44576 26986 44640
rect 27050 44576 27066 44640
rect 27130 44576 27146 44640
rect 27210 44576 27226 44640
rect 27290 44576 27298 44640
rect 26978 43552 27298 44576
rect 26978 43488 26986 43552
rect 27050 43488 27066 43552
rect 27130 43488 27146 43552
rect 27210 43488 27226 43552
rect 27290 43488 27298 43552
rect 26978 42464 27298 43488
rect 26978 42400 26986 42464
rect 27050 42400 27066 42464
rect 27130 42400 27146 42464
rect 27210 42400 27226 42464
rect 27290 42400 27298 42464
rect 23611 42260 23677 42261
rect 23611 42196 23612 42260
rect 23676 42196 23677 42260
rect 23611 42195 23677 42196
rect 19864 41856 19872 41920
rect 19936 41856 19952 41920
rect 20016 41856 20032 41920
rect 20096 41856 20112 41920
rect 20176 41856 20184 41920
rect 19864 40832 20184 41856
rect 19864 40768 19872 40832
rect 19936 40768 19952 40832
rect 20016 40768 20032 40832
rect 20096 40768 20112 40832
rect 20176 40768 20184 40832
rect 19864 39744 20184 40768
rect 19864 39680 19872 39744
rect 19936 39680 19952 39744
rect 20016 39680 20032 39744
rect 20096 39680 20112 39744
rect 20176 39680 20184 39744
rect 19864 38656 20184 39680
rect 20483 39404 20549 39405
rect 20483 39340 20484 39404
rect 20548 39340 20549 39404
rect 20483 39339 20549 39340
rect 20299 38860 20365 38861
rect 20299 38796 20300 38860
rect 20364 38796 20365 38860
rect 20299 38795 20365 38796
rect 19864 38592 19872 38656
rect 19936 38592 19952 38656
rect 20016 38592 20032 38656
rect 20096 38592 20112 38656
rect 20176 38592 20184 38656
rect 19864 37568 20184 38592
rect 20302 37773 20362 38795
rect 20299 37772 20365 37773
rect 20299 37708 20300 37772
rect 20364 37708 20365 37772
rect 20299 37707 20365 37708
rect 19864 37504 19872 37568
rect 19936 37504 19952 37568
rect 20016 37504 20032 37568
rect 20096 37504 20112 37568
rect 20176 37504 20184 37568
rect 19864 36480 20184 37504
rect 20302 36821 20362 37707
rect 20299 36820 20365 36821
rect 20299 36756 20300 36820
rect 20364 36756 20365 36820
rect 20299 36755 20365 36756
rect 19864 36416 19872 36480
rect 19936 36416 19952 36480
rect 20016 36416 20032 36480
rect 20096 36416 20112 36480
rect 20176 36416 20184 36480
rect 19864 35392 20184 36416
rect 19864 35328 19872 35392
rect 19936 35328 19952 35392
rect 20016 35328 20032 35392
rect 20096 35328 20112 35392
rect 20176 35328 20184 35392
rect 19864 34304 20184 35328
rect 19864 34240 19872 34304
rect 19936 34240 19952 34304
rect 20016 34240 20032 34304
rect 20096 34240 20112 34304
rect 20176 34240 20184 34304
rect 19864 33216 20184 34240
rect 19864 33152 19872 33216
rect 19936 33152 19952 33216
rect 20016 33152 20032 33216
rect 20096 33152 20112 33216
rect 20176 33152 20184 33216
rect 19864 32128 20184 33152
rect 19864 32064 19872 32128
rect 19936 32064 19952 32128
rect 20016 32064 20032 32128
rect 20096 32064 20112 32128
rect 20176 32064 20184 32128
rect 19864 31040 20184 32064
rect 20299 31924 20365 31925
rect 20299 31860 20300 31924
rect 20364 31860 20365 31924
rect 20299 31859 20365 31860
rect 20302 31653 20362 31859
rect 20299 31652 20365 31653
rect 20299 31588 20300 31652
rect 20364 31588 20365 31652
rect 20299 31587 20365 31588
rect 19864 30976 19872 31040
rect 19936 30976 19952 31040
rect 20016 30976 20032 31040
rect 20096 30976 20112 31040
rect 20176 30976 20184 31040
rect 19864 29952 20184 30976
rect 19864 29888 19872 29952
rect 19936 29888 19952 29952
rect 20016 29888 20032 29952
rect 20096 29888 20112 29952
rect 20176 29888 20184 29952
rect 19864 28864 20184 29888
rect 19864 28800 19872 28864
rect 19936 28800 19952 28864
rect 20016 28800 20032 28864
rect 20096 28800 20112 28864
rect 20176 28800 20184 28864
rect 19864 27776 20184 28800
rect 19864 27712 19872 27776
rect 19936 27712 19952 27776
rect 20016 27712 20032 27776
rect 20096 27712 20112 27776
rect 20176 27712 20184 27776
rect 19864 26688 20184 27712
rect 19864 26624 19872 26688
rect 19936 26624 19952 26688
rect 20016 26624 20032 26688
rect 20096 26624 20112 26688
rect 20176 26624 20184 26688
rect 19864 25600 20184 26624
rect 19864 25536 19872 25600
rect 19936 25536 19952 25600
rect 20016 25536 20032 25600
rect 20096 25536 20112 25600
rect 20176 25536 20184 25600
rect 19864 24512 20184 25536
rect 19864 24448 19872 24512
rect 19936 24448 19952 24512
rect 20016 24448 20032 24512
rect 20096 24448 20112 24512
rect 20176 24448 20184 24512
rect 19864 23424 20184 24448
rect 20486 23901 20546 39339
rect 20667 37228 20733 37229
rect 20667 37164 20668 37228
rect 20732 37164 20733 37228
rect 20667 37163 20733 37164
rect 20670 29205 20730 37163
rect 21955 36684 22021 36685
rect 21955 36620 21956 36684
rect 22020 36620 22021 36684
rect 21955 36619 22021 36620
rect 20667 29204 20733 29205
rect 20667 29140 20668 29204
rect 20732 29140 20733 29204
rect 20667 29139 20733 29140
rect 21958 28661 22018 36619
rect 23614 30293 23674 42195
rect 24531 41580 24597 41581
rect 24531 41516 24532 41580
rect 24596 41516 24597 41580
rect 24531 41515 24597 41516
rect 23611 30292 23677 30293
rect 23611 30228 23612 30292
rect 23676 30228 23677 30292
rect 23611 30227 23677 30228
rect 21955 28660 22021 28661
rect 21955 28596 21956 28660
rect 22020 28596 22021 28660
rect 21955 28595 22021 28596
rect 24534 28117 24594 41515
rect 26978 41376 27298 42400
rect 26978 41312 26986 41376
rect 27050 41312 27066 41376
rect 27130 41312 27146 41376
rect 27210 41312 27226 41376
rect 27290 41312 27298 41376
rect 26978 40288 27298 41312
rect 26978 40224 26986 40288
rect 27050 40224 27066 40288
rect 27130 40224 27146 40288
rect 27210 40224 27226 40288
rect 27290 40224 27298 40288
rect 26978 39200 27298 40224
rect 26978 39136 26986 39200
rect 27050 39136 27066 39200
rect 27130 39136 27146 39200
rect 27210 39136 27226 39200
rect 27290 39136 27298 39200
rect 26978 38112 27298 39136
rect 26978 38048 26986 38112
rect 27050 38048 27066 38112
rect 27130 38048 27146 38112
rect 27210 38048 27226 38112
rect 27290 38048 27298 38112
rect 26978 37024 27298 38048
rect 26978 36960 26986 37024
rect 27050 36960 27066 37024
rect 27130 36960 27146 37024
rect 27210 36960 27226 37024
rect 27290 36960 27298 37024
rect 26978 35936 27298 36960
rect 26978 35872 26986 35936
rect 27050 35872 27066 35936
rect 27130 35872 27146 35936
rect 27210 35872 27226 35936
rect 27290 35872 27298 35936
rect 26978 34848 27298 35872
rect 26978 34784 26986 34848
rect 27050 34784 27066 34848
rect 27130 34784 27146 34848
rect 27210 34784 27226 34848
rect 27290 34784 27298 34848
rect 26978 33760 27298 34784
rect 26978 33696 26986 33760
rect 27050 33696 27066 33760
rect 27130 33696 27146 33760
rect 27210 33696 27226 33760
rect 27290 33696 27298 33760
rect 26978 32672 27298 33696
rect 26978 32608 26986 32672
rect 27050 32608 27066 32672
rect 27130 32608 27146 32672
rect 27210 32608 27226 32672
rect 27290 32608 27298 32672
rect 26978 31584 27298 32608
rect 26978 31520 26986 31584
rect 27050 31520 27066 31584
rect 27130 31520 27146 31584
rect 27210 31520 27226 31584
rect 27290 31520 27298 31584
rect 26739 30700 26805 30701
rect 26739 30636 26740 30700
rect 26804 30636 26805 30700
rect 26739 30635 26805 30636
rect 24531 28116 24597 28117
rect 24531 28052 24532 28116
rect 24596 28052 24597 28116
rect 24531 28051 24597 28052
rect 20483 23900 20549 23901
rect 20483 23836 20484 23900
rect 20548 23836 20549 23900
rect 20483 23835 20549 23836
rect 19864 23360 19872 23424
rect 19936 23360 19952 23424
rect 20016 23360 20032 23424
rect 20096 23360 20112 23424
rect 20176 23360 20184 23424
rect 19864 22336 20184 23360
rect 19864 22272 19872 22336
rect 19936 22272 19952 22336
rect 20016 22272 20032 22336
rect 20096 22272 20112 22336
rect 20176 22272 20184 22336
rect 19864 21248 20184 22272
rect 19864 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20184 21248
rect 19864 20160 20184 21184
rect 19864 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20184 20160
rect 19864 19072 20184 20096
rect 19864 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20184 19072
rect 19864 17984 20184 19008
rect 19864 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20184 17984
rect 19864 16896 20184 17920
rect 19864 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20184 16896
rect 19864 15808 20184 16832
rect 26742 16693 26802 30635
rect 26978 30496 27298 31520
rect 26978 30432 26986 30496
rect 27050 30432 27066 30496
rect 27130 30432 27146 30496
rect 27210 30432 27226 30496
rect 27290 30432 27298 30496
rect 26978 29408 27298 30432
rect 26978 29344 26986 29408
rect 27050 29344 27066 29408
rect 27130 29344 27146 29408
rect 27210 29344 27226 29408
rect 27290 29344 27298 29408
rect 26978 28320 27298 29344
rect 26978 28256 26986 28320
rect 27050 28256 27066 28320
rect 27130 28256 27146 28320
rect 27210 28256 27226 28320
rect 27290 28256 27298 28320
rect 26978 27232 27298 28256
rect 26978 27168 26986 27232
rect 27050 27168 27066 27232
rect 27130 27168 27146 27232
rect 27210 27168 27226 27232
rect 27290 27168 27298 27232
rect 26978 26144 27298 27168
rect 26978 26080 26986 26144
rect 27050 26080 27066 26144
rect 27130 26080 27146 26144
rect 27210 26080 27226 26144
rect 27290 26080 27298 26144
rect 26978 25056 27298 26080
rect 26978 24992 26986 25056
rect 27050 24992 27066 25056
rect 27130 24992 27146 25056
rect 27210 24992 27226 25056
rect 27290 24992 27298 25056
rect 26978 23968 27298 24992
rect 26978 23904 26986 23968
rect 27050 23904 27066 23968
rect 27130 23904 27146 23968
rect 27210 23904 27226 23968
rect 27290 23904 27298 23968
rect 26978 22880 27298 23904
rect 26978 22816 26986 22880
rect 27050 22816 27066 22880
rect 27130 22816 27146 22880
rect 27210 22816 27226 22880
rect 27290 22816 27298 22880
rect 26978 21792 27298 22816
rect 26978 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27298 21792
rect 26978 20704 27298 21728
rect 26978 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27298 20704
rect 26978 19616 27298 20640
rect 26978 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27298 19616
rect 26978 18528 27298 19552
rect 26978 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27298 18528
rect 26978 17440 27298 18464
rect 26978 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27298 17440
rect 26739 16692 26805 16693
rect 26739 16628 26740 16692
rect 26804 16628 26805 16692
rect 26739 16627 26805 16628
rect 19864 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20184 15808
rect 19864 14720 20184 15744
rect 19864 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20184 14720
rect 19864 13632 20184 14656
rect 19864 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20184 13632
rect 19864 12544 20184 13568
rect 19864 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20184 12544
rect 19864 11456 20184 12480
rect 19864 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20184 11456
rect 19864 10368 20184 11392
rect 19864 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20184 10368
rect 19864 9280 20184 10304
rect 19864 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20184 9280
rect 19864 8192 20184 9216
rect 19864 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20184 8192
rect 19864 7104 20184 8128
rect 19864 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20184 7104
rect 19864 6016 20184 7040
rect 19864 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20184 6016
rect 19864 4928 20184 5952
rect 19864 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20184 4928
rect 19864 3840 20184 4864
rect 19864 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20184 3840
rect 19864 2752 20184 3776
rect 19864 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20184 2752
rect 19864 1664 20184 2688
rect 19864 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20184 1664
rect 19864 576 20184 1600
rect 19864 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20184 576
rect 19864 496 20184 512
rect 26978 16352 27298 17376
rect 26978 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27298 16352
rect 26978 15264 27298 16288
rect 26978 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27298 15264
rect 26978 14176 27298 15200
rect 26978 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27298 14176
rect 26978 13088 27298 14112
rect 26978 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27298 13088
rect 26978 12000 27298 13024
rect 26978 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27298 12000
rect 26978 10912 27298 11936
rect 26978 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27298 10912
rect 26978 9824 27298 10848
rect 26978 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27298 9824
rect 26978 8736 27298 9760
rect 26978 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27298 8736
rect 26978 7648 27298 8672
rect 26978 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27298 7648
rect 26978 6560 27298 7584
rect 26978 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27298 6560
rect 26978 5472 27298 6496
rect 26978 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27298 5472
rect 26978 4384 27298 5408
rect 26978 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27298 4384
rect 26978 3296 27298 4320
rect 26978 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27298 3296
rect 26978 2208 27298 3232
rect 26978 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27298 2208
rect 26978 1120 27298 2144
rect 26978 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27298 1120
rect 26978 496 27298 1056
rect 27638 44096 27958 44656
rect 28211 44644 28212 44708
rect 28276 44644 28277 44708
rect 28211 44643 28277 44644
rect 27638 44032 27646 44096
rect 27710 44032 27726 44096
rect 27790 44032 27806 44096
rect 27870 44032 27886 44096
rect 27950 44032 27958 44096
rect 27638 43008 27958 44032
rect 27638 42944 27646 43008
rect 27710 42944 27726 43008
rect 27790 42944 27806 43008
rect 27870 42944 27886 43008
rect 27950 42944 27958 43008
rect 27638 41920 27958 42944
rect 27638 41856 27646 41920
rect 27710 41856 27726 41920
rect 27790 41856 27806 41920
rect 27870 41856 27886 41920
rect 27950 41856 27958 41920
rect 27638 40832 27958 41856
rect 27638 40768 27646 40832
rect 27710 40768 27726 40832
rect 27790 40768 27806 40832
rect 27870 40768 27886 40832
rect 27950 40768 27958 40832
rect 27638 39744 27958 40768
rect 27638 39680 27646 39744
rect 27710 39680 27726 39744
rect 27790 39680 27806 39744
rect 27870 39680 27886 39744
rect 27950 39680 27958 39744
rect 27638 38656 27958 39680
rect 27638 38592 27646 38656
rect 27710 38592 27726 38656
rect 27790 38592 27806 38656
rect 27870 38592 27886 38656
rect 27950 38592 27958 38656
rect 27638 37568 27958 38592
rect 27638 37504 27646 37568
rect 27710 37504 27726 37568
rect 27790 37504 27806 37568
rect 27870 37504 27886 37568
rect 27950 37504 27958 37568
rect 27638 36480 27958 37504
rect 27638 36416 27646 36480
rect 27710 36416 27726 36480
rect 27790 36416 27806 36480
rect 27870 36416 27886 36480
rect 27950 36416 27958 36480
rect 27638 35392 27958 36416
rect 27638 35328 27646 35392
rect 27710 35328 27726 35392
rect 27790 35328 27806 35392
rect 27870 35328 27886 35392
rect 27950 35328 27958 35392
rect 27638 34304 27958 35328
rect 27638 34240 27646 34304
rect 27710 34240 27726 34304
rect 27790 34240 27806 34304
rect 27870 34240 27886 34304
rect 27950 34240 27958 34304
rect 27638 33216 27958 34240
rect 27638 33152 27646 33216
rect 27710 33152 27726 33216
rect 27790 33152 27806 33216
rect 27870 33152 27886 33216
rect 27950 33152 27958 33216
rect 27638 32128 27958 33152
rect 27638 32064 27646 32128
rect 27710 32064 27726 32128
rect 27790 32064 27806 32128
rect 27870 32064 27886 32128
rect 27950 32064 27958 32128
rect 27638 31040 27958 32064
rect 27638 30976 27646 31040
rect 27710 30976 27726 31040
rect 27790 30976 27806 31040
rect 27870 30976 27886 31040
rect 27950 30976 27958 31040
rect 27638 29952 27958 30976
rect 27638 29888 27646 29952
rect 27710 29888 27726 29952
rect 27790 29888 27806 29952
rect 27870 29888 27886 29952
rect 27950 29888 27958 29952
rect 27638 28864 27958 29888
rect 27638 28800 27646 28864
rect 27710 28800 27726 28864
rect 27790 28800 27806 28864
rect 27870 28800 27886 28864
rect 27950 28800 27958 28864
rect 27638 27776 27958 28800
rect 28766 28525 28826 45152
rect 29318 44952 29378 45152
rect 28763 28524 28829 28525
rect 28763 28460 28764 28524
rect 28828 28460 28829 28524
rect 28763 28459 28829 28460
rect 27638 27712 27646 27776
rect 27710 27712 27726 27776
rect 27790 27712 27806 27776
rect 27870 27712 27886 27776
rect 27950 27712 27958 27776
rect 27638 26688 27958 27712
rect 27638 26624 27646 26688
rect 27710 26624 27726 26688
rect 27790 26624 27806 26688
rect 27870 26624 27886 26688
rect 27950 26624 27958 26688
rect 27638 25600 27958 26624
rect 27638 25536 27646 25600
rect 27710 25536 27726 25600
rect 27790 25536 27806 25600
rect 27870 25536 27886 25600
rect 27950 25536 27958 25600
rect 27638 24512 27958 25536
rect 27638 24448 27646 24512
rect 27710 24448 27726 24512
rect 27790 24448 27806 24512
rect 27870 24448 27886 24512
rect 27950 24448 27958 24512
rect 27638 23424 27958 24448
rect 27638 23360 27646 23424
rect 27710 23360 27726 23424
rect 27790 23360 27806 23424
rect 27870 23360 27886 23424
rect 27950 23360 27958 23424
rect 27638 22336 27958 23360
rect 27638 22272 27646 22336
rect 27710 22272 27726 22336
rect 27790 22272 27806 22336
rect 27870 22272 27886 22336
rect 27950 22272 27958 22336
rect 27638 21248 27958 22272
rect 27638 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27958 21248
rect 27638 20160 27958 21184
rect 27638 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27958 20160
rect 27638 19072 27958 20096
rect 27638 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27958 19072
rect 27638 17984 27958 19008
rect 27638 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27958 17984
rect 27638 16896 27958 17920
rect 27638 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27958 16896
rect 27638 15808 27958 16832
rect 27638 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27958 15808
rect 27638 14720 27958 15744
rect 27638 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27958 14720
rect 27638 13632 27958 14656
rect 27638 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27958 13632
rect 27638 12544 27958 13568
rect 27638 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27958 12544
rect 27638 11456 27958 12480
rect 27638 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27958 11456
rect 27638 10368 27958 11392
rect 27638 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27958 10368
rect 27638 9280 27958 10304
rect 27638 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27958 9280
rect 27638 8192 27958 9216
rect 27638 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27958 8192
rect 27638 7104 27958 8128
rect 27638 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27958 7104
rect 27638 6016 27958 7040
rect 27638 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27958 6016
rect 27638 4928 27958 5952
rect 27638 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27958 4928
rect 27638 3840 27958 4864
rect 27638 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27958 3840
rect 27638 2752 27958 3776
rect 27638 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27958 2752
rect 27638 1664 27958 2688
rect 27638 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27958 1664
rect 27638 576 27958 1600
rect 27638 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27958 576
rect 27638 496 27958 512
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1
transform 1 0 9752 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1
transform -1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1
transform -1 0 26680 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1
transform 1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1
transform -1 0 27324 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1
transform -1 0 27140 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1
transform -1 0 26312 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1
transform 1 0 26036 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1
transform -1 0 26680 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1
transform 1 0 22724 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1
transform 1 0 19780 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1
transform 1 0 20240 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1
transform -1 0 17112 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1
transform -1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1
transform -1 0 16560 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1
transform -1 0 17940 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1
transform -1 0 18584 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1
transform 1 0 13248 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1
transform 1 0 21252 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1
transform 1 0 21988 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1
transform 1 0 26956 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1
transform 1 0 24656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1
transform 1 0 25208 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1
transform -1 0 21436 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1
transform 1 0 26956 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1
transform 1 0 25300 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1
transform 1 0 26864 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1
transform 1 0 24472 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753__1
timestamp 1
transform -1 0 12420 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753__2
timestamp 1
transform 1 0 13984 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0754_
timestamp 1
transform -1 0 14536 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _0755_
timestamp 1
transform -1 0 18308 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _0756_
timestamp 1
transform -1 0 20148 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__mux4_1  _0757_
timestamp 1
transform -1 0 29532 0 -1 39712
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0758_
timestamp 1
transform -1 0 27692 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0759_
timestamp 1
transform 1 0 25208 0 1 38624
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _0760_
timestamp 1
transform 1 0 26404 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _0761_
timestamp 1
transform -1 0 29440 0 -1 35360
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0762_
timestamp 1
transform -1 0 30084 0 -1 37536
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1
transform 1 0 27324 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _0764_
timestamp 1
transform 1 0 25668 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0765_
timestamp 1
transform 1 0 25760 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0766_
timestamp 1
transform 1 0 24472 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0767_
timestamp 1
transform 1 0 25576 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0768_
timestamp 1
transform 1 0 25852 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0769_
timestamp 1
transform -1 0 27416 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0770_
timestamp 1
transform 1 0 27416 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1
transform 1 0 26496 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 1
transform 1 0 26404 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0773_
timestamp 1
transform 1 0 25116 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0774_
timestamp 1
transform -1 0 26956 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0775_
timestamp 1
transform 1 0 25484 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0776_
timestamp 1
transform 1 0 25208 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0777_
timestamp 1
transform 1 0 25116 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0778_
timestamp 1
transform -1 0 26312 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0779_
timestamp 1
transform 1 0 24748 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0780_
timestamp 1
transform 1 0 25024 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0781_
timestamp 1
transform 1 0 24104 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0782_
timestamp 1
transform 1 0 25852 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_1  _0783_
timestamp 1
transform 1 0 25392 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0784_
timestamp 1
transform -1 0 26864 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_1  _0785_
timestamp 1
transform 1 0 25576 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0786_
timestamp 1
transform -1 0 27232 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0787_
timestamp 1
transform 1 0 26404 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0788_
timestamp 1
transform 1 0 26404 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0789_
timestamp 1
transform 1 0 26680 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0790_
timestamp 1
transform 1 0 26404 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _0791_
timestamp 1
transform -1 0 24380 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0792_
timestamp 1
transform 1 0 21620 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0793_
timestamp 1
transform 1 0 21252 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0794_
timestamp 1
transform -1 0 20792 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0795_
timestamp 1
transform 1 0 22356 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0796_
timestamp 1
transform -1 0 22448 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0797_
timestamp 1
transform -1 0 23828 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0798_
timestamp 1
transform -1 0 24288 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0799_
timestamp 1
transform -1 0 20424 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1
transform -1 0 20240 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0801_
timestamp 1
transform 1 0 21712 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1
transform -1 0 20884 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0803_
timestamp 1
transform 1 0 21344 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0804_
timestamp 1
transform -1 0 25300 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0805_
timestamp 1
transform 1 0 23276 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0806_
timestamp 1
transform 1 0 23828 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0807_
timestamp 1
transform -1 0 24288 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0808_
timestamp 1
transform 1 0 23828 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0809_
timestamp 1
transform 1 0 23736 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0810_
timestamp 1
transform -1 0 24196 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0811_
timestamp 1
transform 1 0 23828 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_4  _0812_
timestamp 1
transform 1 0 19044 0 1 25568
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_2  _0813_
timestamp 1
transform 1 0 20700 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0814_
timestamp 1
transform 1 0 20240 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1
transform -1 0 20700 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0816_
timestamp 1
transform 1 0 21252 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1
transform -1 0 20976 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0818_
timestamp 1
transform -1 0 22816 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0819_
timestamp 1
transform -1 0 22540 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0820_
timestamp 1
transform 1 0 22632 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0821_
timestamp 1
transform 1 0 22356 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1
transform 1 0 21988 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0823_
timestamp 1
transform 1 0 21436 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0824_
timestamp 1
transform 1 0 21068 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0825_
timestamp 1
transform 1 0 19964 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1
transform -1 0 19228 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0827_
timestamp 1
transform 1 0 22448 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0828_
timestamp 1
transform 1 0 22172 0 -1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1
transform 1 0 26036 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0830_
timestamp 1
transform 1 0 24564 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0831_
timestamp 1
transform 1 0 25024 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0832_
timestamp 1
transform -1 0 26128 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0833_
timestamp 1
transform 1 0 24656 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0834_
timestamp 1
transform 1 0 23644 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0835_
timestamp 1
transform 1 0 25024 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0836_
timestamp 1
transform -1 0 26036 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0837_
timestamp 1
transform 1 0 26312 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0838_
timestamp 1
transform -1 0 27140 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0839_
timestamp 1
transform 1 0 25576 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0840_
timestamp 1
transform 1 0 27232 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0841_
timestamp 1
transform -1 0 27692 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1
transform 1 0 24748 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0843_
timestamp 1
transform 1 0 26404 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0844_
timestamp 1
transform 1 0 26404 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0845_
timestamp 1
transform -1 0 27876 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0846_
timestamp 1
transform -1 0 27232 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0847_
timestamp 1
transform 1 0 25392 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0848_
timestamp 1
transform 1 0 25484 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_1  _0849_
timestamp 1
transform 1 0 26312 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0850_
timestamp 1
transform -1 0 26588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0851_
timestamp 1
transform 1 0 25392 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0852_
timestamp 1
transform -1 0 25116 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0853_
timestamp 1
transform 1 0 24748 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0854_
timestamp 1
transform 1 0 17940 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _0855_
timestamp 1
transform 1 0 19504 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0856_
timestamp 1
transform 1 0 17940 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1
transform 1 0 15088 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0858_
timestamp 1
transform -1 0 15088 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0859_
timestamp 1
transform 1 0 18216 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0860_
timestamp 1
transform 1 0 18400 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0861_
timestamp 1
transform 1 0 19320 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0862_
timestamp 1
transform -1 0 19872 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0863_
timestamp 1
transform -1 0 13432 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _0864_
timestamp 1
transform -1 0 14168 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0865_
timestamp 1
transform 1 0 13248 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1
transform -1 0 19136 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0867_
timestamp 1
transform -1 0 18492 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0868_
timestamp 1
transform 1 0 18676 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _0869_
timestamp 1
transform -1 0 19136 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0870_
timestamp 1
transform 1 0 18676 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0871_
timestamp 1
transform 1 0 24564 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0872_
timestamp 1
transform -1 0 22908 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0873_
timestamp 1
transform 1 0 21620 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0874_
timestamp 1
transform -1 0 23184 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1
transform -1 0 23368 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0876_
timestamp 1
transform 1 0 22264 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1
transform 1 0 21712 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0878_
timestamp 1
transform 1 0 23828 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0879_
timestamp 1
transform 1 0 23828 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1
transform 1 0 23460 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0881_
timestamp 1
transform -1 0 25300 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0882_
timestamp 1
transform -1 0 26128 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0883_
timestamp 1
transform 1 0 23552 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1
transform 1 0 23276 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0885_
timestamp 1
transform -1 0 25300 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0886_
timestamp 1
transform -1 0 23644 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1
transform -1 0 19412 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0888_
timestamp 1
transform 1 0 18860 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0889_
timestamp 1
transform -1 0 21068 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0890_
timestamp 1
transform 1 0 20148 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1
transform -1 0 19872 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0892_
timestamp 1
transform 1 0 21252 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0893_
timestamp 1
transform 1 0 20700 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0894_
timestamp 1
transform 1 0 19688 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1
transform -1 0 19688 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0896_
timestamp 1
transform 1 0 21528 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0897_
timestamp 1
transform 1 0 21252 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1
transform -1 0 20976 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0899_
timestamp 1
transform 1 0 20240 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1
transform -1 0 19872 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0901_
timestamp 1
transform 1 0 21252 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0902_
timestamp 1
transform -1 0 21068 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0903_
timestamp 1
transform -1 0 21528 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0904_
timestamp 1
transform -1 0 20148 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0905_
timestamp 1
transform -1 0 19320 0 -1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0906_
timestamp 1
transform 1 0 19044 0 -1 37536
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1
transform -1 0 24104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0908_
timestamp 1
transform -1 0 24748 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1
transform 1 0 23920 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0910_
timestamp 1
transform -1 0 24840 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1
transform 1 0 24748 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0912_
timestamp 1
transform -1 0 23920 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1
transform -1 0 24012 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0914_
timestamp 1
transform -1 0 23736 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0915_
timestamp 1
transform -1 0 23828 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _0916_
timestamp 1
transform 1 0 26404 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0917_
timestamp 1
transform 1 0 27324 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0918_
timestamp 1
transform 1 0 27416 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0919_
timestamp 1
transform 1 0 27784 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1
transform -1 0 28336 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0921_
timestamp 1
transform -1 0 28060 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1
transform 1 0 27140 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1
transform 1 0 27140 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0924_
timestamp 1
transform -1 0 26680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0925_
timestamp 1
transform -1 0 27140 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1
transform -1 0 26312 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1
transform 1 0 25760 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0928_
timestamp 1
transform -1 0 25392 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1
transform -1 0 24288 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1
transform -1 0 24840 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0931_
timestamp 1
transform -1 0 24196 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0932_
timestamp 1
transform 1 0 23276 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1
transform 1 0 25300 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0934_
timestamp 1
transform 1 0 24288 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0935_
timestamp 1
transform -1 0 26312 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0936_
timestamp 1
transform -1 0 25668 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 1
transform -1 0 27416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0938_
timestamp 1
transform 1 0 26680 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0939_
timestamp 1
transform -1 0 27968 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0940_
timestamp 1
transform -1 0 28796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 1
transform -1 0 28704 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0942_
timestamp 1
transform 1 0 27600 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0943_
timestamp 1
transform 1 0 27508 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1
transform -1 0 28428 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1
transform -1 0 28244 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0946_
timestamp 1
transform 1 0 28060 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0947_
timestamp 1
transform -1 0 28796 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1
transform 1 0 29624 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0949_
timestamp 1
transform 1 0 28980 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0950_
timestamp 1
transform -1 0 27784 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 1
transform -1 0 27416 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0952_
timestamp 1
transform 1 0 28152 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0953_
timestamp 1
transform 1 0 27968 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0954_
timestamp 1
transform 1 0 27692 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0955_
timestamp 1
transform -1 0 28152 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0956_
timestamp 1
transform 1 0 28060 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0957_
timestamp 1
transform -1 0 27692 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0958_
timestamp 1
transform -1 0 28244 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0959_
timestamp 1
transform 1 0 27692 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1
transform -1 0 28152 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0961_
timestamp 1
transform -1 0 28244 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0962_
timestamp 1
transform 1 0 27140 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0963_
timestamp 1
transform -1 0 27048 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0964_
timestamp 1
transform 1 0 26680 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0965_
timestamp 1
transform 1 0 29440 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1
transform 1 0 29440 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0967_
timestamp 1
transform -1 0 30728 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1
transform -1 0 31004 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0969_
timestamp 1
transform 1 0 29348 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0970_
timestamp 1
transform 1 0 28244 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1
transform -1 0 28888 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0972_
timestamp 1
transform -1 0 26864 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1
transform -1 0 25392 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0974_
timestamp 1
transform 1 0 25208 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0975_
timestamp 1
transform 1 0 24656 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0976_
timestamp 1
transform 1 0 26404 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0977_
timestamp 1
transform 1 0 25668 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0978_
timestamp 1
transform -1 0 25208 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0979_
timestamp 1
transform 1 0 26220 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0980_
timestamp 1
transform -1 0 26956 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 1
transform -1 0 26128 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0982_
timestamp 1
transform 1 0 27784 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0983_
timestamp 1
transform 1 0 27048 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0984_
timestamp 1
transform -1 0 28612 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0985_
timestamp 1
transform -1 0 28244 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0986_
timestamp 1
transform -1 0 29348 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1
transform -1 0 28888 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0988_
timestamp 1
transform 1 0 30360 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1
transform 1 0 30728 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0990_
timestamp 1
transform -1 0 29900 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0991_
timestamp 1
transform 1 0 30176 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0992_
timestamp 1
transform -1 0 31096 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0993_
timestamp 1
transform 1 0 31096 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0994_
timestamp 1
transform 1 0 30636 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0995_
timestamp 1
transform -1 0 30636 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0996_
timestamp 1
transform -1 0 31188 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0997_
timestamp 1
transform -1 0 30820 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0998_
timestamp 1
transform 1 0 29256 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0999_
timestamp 1
transform 1 0 28612 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1000_
timestamp 1
transform 1 0 27600 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1001_
timestamp 1
transform 1 0 27048 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1002_
timestamp 1
transform -1 0 28796 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1003_
timestamp 1
transform -1 0 28428 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1004_
timestamp 1
transform -1 0 28060 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1005_
timestamp 1
transform -1 0 16376 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1
transform -1 0 16836 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1007_
timestamp 1
transform 1 0 13524 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1
transform 1 0 14628 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1009_
timestamp 1
transform -1 0 14628 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1010_
timestamp 1
transform 1 0 17020 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1011_
timestamp 1
transform -1 0 17020 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1
transform -1 0 18584 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1013_
timestamp 1
transform -1 0 17664 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1014_
timestamp 1
transform -1 0 18860 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1015_
timestamp 1
transform -1 0 18216 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1
transform 1 0 19964 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1
transform 1 0 19780 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1
transform 1 0 20608 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1019_
timestamp 1
transform 1 0 20424 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1
transform 1 0 19504 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1021_
timestamp 1
transform -1 0 20700 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1
transform 1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _1023_
timestamp 1
transform 1 0 19320 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1
transform 1 0 20056 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1025_
timestamp 1
transform -1 0 21068 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1
transform 1 0 19412 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1027_
timestamp 1
transform -1 0 20884 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1028_
timestamp 1
transform 1 0 20148 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1029_
timestamp 1
transform -1 0 21160 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1
transform 1 0 21252 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1
transform -1 0 21988 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1032_
timestamp 1
transform -1 0 18216 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1033_
timestamp 1
transform -1 0 18676 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1034_
timestamp 1
transform 1 0 15548 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1035_
timestamp 1
transform 1 0 15364 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1
transform -1 0 15272 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1037_
timestamp 1
transform 1 0 14352 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1038_
timestamp 1
transform -1 0 16284 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1
transform 1 0 14536 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1040_
timestamp 1
transform -1 0 16284 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1041_
timestamp 1
transform -1 0 16008 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1
transform -1 0 17756 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1
transform 1 0 16468 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1
transform 1 0 17296 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1
transform 1 0 17848 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1
transform 1 0 17756 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1047_
timestamp 1
transform 1 0 17572 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1
transform -1 0 18032 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1049_
timestamp 1
transform 1 0 17020 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1050_
timestamp 1
transform 1 0 18124 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1051_
timestamp 1
transform -1 0 18124 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1052_
timestamp 1
transform -1 0 14904 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1053_
timestamp 1
transform 1 0 13064 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1
transform -1 0 14812 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1055_
timestamp 1
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1
transform 1 0 12972 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1057_
timestamp 1
transform 1 0 13708 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1058_
timestamp 1
transform 1 0 12972 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1059_
timestamp 1
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1060_
timestamp 1
transform -1 0 16652 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1061_
timestamp 1
transform -1 0 16928 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1062_
timestamp 1
transform 1 0 14812 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1063_
timestamp 1
transform 1 0 15088 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1064_
timestamp 1
transform -1 0 14444 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1
transform -1 0 14536 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1
transform 1 0 15456 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1
transform 1 0 15456 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1
transform -1 0 9292 0 1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1069_
timestamp 1
transform 1 0 20424 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1
transform -1 0 17388 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1071_
timestamp 1
transform -1 0 19504 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1072_
timestamp 1
transform -1 0 20148 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1073_
timestamp 1
transform 1 0 22632 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1074_
timestamp 1
transform 1 0 17296 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1075_
timestamp 1
transform 1 0 23276 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1076_
timestamp 1
transform 1 0 16376 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1077_
timestamp 1
transform -1 0 19688 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1078_
timestamp 1
transform -1 0 18492 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _1079_
timestamp 1
transform -1 0 18124 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _1080_
timestamp 1
transform 1 0 17756 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1081_
timestamp 1
transform -1 0 15456 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1082_
timestamp 1
transform -1 0 15916 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1083_
timestamp 1
transform 1 0 17020 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1084_
timestamp 1
transform 1 0 16284 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1085_
timestamp 1
transform -1 0 16008 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1
transform 1 0 15272 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1087_
timestamp 1
transform -1 0 16744 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1088_
timestamp 1
transform 1 0 15364 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1089_
timestamp 1
transform 1 0 14812 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1090_
timestamp 1
transform -1 0 17020 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1091_
timestamp 1
transform -1 0 16560 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1
transform 1 0 16008 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1093_
timestamp 1
transform 1 0 15272 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1094_
timestamp 1
transform -1 0 15824 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1095_
timestamp 1
transform -1 0 18124 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1096_
timestamp 1
transform 1 0 17204 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1097_
timestamp 1
transform 1 0 15548 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1098_
timestamp 1
transform 1 0 16376 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1
transform -1 0 16008 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1100_
timestamp 1
transform -1 0 16836 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1101_
timestamp 1
transform 1 0 16560 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1102_
timestamp 1
transform 1 0 16100 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1103_
timestamp 1
transform 1 0 15548 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1104_
timestamp 1
transform 1 0 15272 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1105_
timestamp 1
transform 1 0 17848 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1106_
timestamp 1
transform -1 0 17480 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1
transform -1 0 16560 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1108_
timestamp 1
transform -1 0 15364 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1109_
timestamp 1
transform 1 0 15364 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1110_
timestamp 1
transform -1 0 16008 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 1
transform -1 0 15180 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1112_
timestamp 1
transform -1 0 14720 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1113_
timestamp 1
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1115_
timestamp 1
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1116_
timestamp 1
transform -1 0 17296 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1117_
timestamp 1
transform 1 0 17664 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1118_
timestamp 1
transform 1 0 18768 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1119_
timestamp 1
transform 1 0 18676 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1120_
timestamp 1
transform 1 0 19228 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1121_
timestamp 1
transform -1 0 17388 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1122_
timestamp 1
transform -1 0 16008 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1
transform 1 0 15732 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_4  _1124_
timestamp 1
transform 1 0 14168 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1
transform -1 0 17940 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1
transform 1 0 17848 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1127_
timestamp 1
transform 1 0 17848 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1128_
timestamp 1
transform 1 0 17020 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1129_
timestamp 1
transform -1 0 18676 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1130_
timestamp 1
transform 1 0 18676 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 1
transform -1 0 16008 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1132_
timestamp 1
transform 1 0 17296 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1133_
timestamp 1
transform -1 0 16928 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1134_
timestamp 1
transform -1 0 18032 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _1135_
timestamp 1
transform -1 0 17480 0 1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1136_
timestamp 1
transform 1 0 15916 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1
transform -1 0 15364 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1138_
timestamp 1
transform -1 0 13984 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1139_
timestamp 1
transform 1 0 14260 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1140_
timestamp 1
transform -1 0 12144 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1141_
timestamp 1
transform 1 0 12052 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 1
transform 1 0 11500 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1
transform 1 0 11408 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1144_
timestamp 1
transform 1 0 11316 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 1
transform -1 0 13432 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1146_
timestamp 1
transform 1 0 12604 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1147_
timestamp 1
transform 1 0 15272 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1148_
timestamp 1
transform 1 0 12880 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1149_
timestamp 1
transform 1 0 15824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1150_
timestamp 1
transform 1 0 15272 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1151_
timestamp 1
transform 1 0 16192 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1152_
timestamp 1
transform -1 0 17388 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1153_
timestamp 1
transform 1 0 15272 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1154_
timestamp 1
transform 1 0 18492 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1155_
timestamp 1
transform 1 0 17940 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1156_
timestamp 1
transform 1 0 18032 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1157_
timestamp 1
transform 1 0 18676 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1158_
timestamp 1
transform 1 0 17388 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1159_
timestamp 1
transform -1 0 17388 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1160_
timestamp 1
transform 1 0 16928 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1161_
timestamp 1
transform -1 0 16744 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1162_
timestamp 1
transform -1 0 15824 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1163_
timestamp 1
transform 1 0 15180 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1164_
timestamp 1
transform 1 0 15824 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1165_
timestamp 1
transform -1 0 18400 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1166_
timestamp 1
transform 1 0 16836 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1167_
timestamp 1
transform -1 0 17020 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 1
transform -1 0 16928 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1169_
timestamp 1
transform -1 0 19136 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1170_
timestamp 1
transform 1 0 17388 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1171_
timestamp 1
transform 1 0 15916 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1172_
timestamp 1
transform 1 0 14904 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1173_
timestamp 1
transform 1 0 17204 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1174_
timestamp 1
transform 1 0 17020 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1
transform 1 0 15364 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1176_
timestamp 1
transform 1 0 16100 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1177_
timestamp 1
transform 1 0 14720 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1178_
timestamp 1
transform -1 0 15732 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1179_
timestamp 1
transform 1 0 16192 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1180_
timestamp 1
transform -1 0 16836 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1181_
timestamp 1
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1182_
timestamp 1
transform 1 0 16928 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1183_
timestamp 1
transform 1 0 17480 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1184_
timestamp 1
transform -1 0 16376 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1185_
timestamp 1
transform 1 0 17572 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1186_
timestamp 1
transform 1 0 13524 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1187_
timestamp 1
transform -1 0 24748 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1188_
timestamp 1
transform 1 0 23828 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1189_
timestamp 1
transform 1 0 24564 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 1
transform 1 0 24472 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1191_
timestamp 1
transform 1 0 25024 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1192_
timestamp 1
transform -1 0 24472 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1193_
timestamp 1
transform 1 0 23828 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1194_
timestamp 1
transform -1 0 22632 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1195_
timestamp 1
transform 1 0 22448 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1196_
timestamp 1
transform 1 0 21804 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1197_
timestamp 1
transform 1 0 14720 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1198_
timestamp 1
transform 1 0 12604 0 -1 26656
box -38 -48 1970 592
use sky130_fd_sc_hd__nand3_1  _1199_
timestamp 1
transform -1 0 13892 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1200_
timestamp 1
transform 1 0 14444 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1201_
timestamp 1
transform -1 0 14720 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1202_
timestamp 1
transform 1 0 14536 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1203_
timestamp 1
transform 1 0 13708 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1204_
timestamp 1
transform 1 0 14260 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1205_
timestamp 1
transform 1 0 13524 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1206_
timestamp 1
transform -1 0 23552 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1207_
timestamp 1
transform 1 0 19136 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1208_
timestamp 1
transform 1 0 23368 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1209_
timestamp 1
transform -1 0 24472 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1210_
timestamp 1
transform 1 0 22724 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1211_
timestamp 1
transform 1 0 24012 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1212_
timestamp 1
transform 1 0 22816 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1213_
timestamp 1
transform 1 0 18492 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1
transform -1 0 15916 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1215_
timestamp 1
transform -1 0 17020 0 1 34272
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1216_
timestamp 1
transform -1 0 16652 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1217_
timestamp 1
transform 1 0 15916 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1218_
timestamp 1
transform -1 0 14168 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1219_
timestamp 1
transform 1 0 14168 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1
transform 1 0 12144 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1221_
timestamp 1
transform 1 0 13432 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1222_
timestamp 1
transform 1 0 12604 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1223_
timestamp 1
transform -1 0 13248 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1224_
timestamp 1
transform -1 0 13524 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1225_
timestamp 1
transform 1 0 12788 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1226_
timestamp 1
transform 1 0 12604 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1227_
timestamp 1
transform 1 0 12604 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1228_
timestamp 1
transform 1 0 12144 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1229_
timestamp 1
transform 1 0 11132 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1230_
timestamp 1
transform -1 0 12512 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1231_
timestamp 1
transform 1 0 11224 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1232_
timestamp 1
transform 1 0 11224 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1233_
timestamp 1
transform -1 0 11224 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1234_
timestamp 1
transform 1 0 11776 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1
transform 1 0 9660 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1236_
timestamp 1
transform -1 0 10856 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp 1
transform 1 0 10948 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1238_
timestamp 1
transform -1 0 10672 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1
transform 1 0 9660 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1
transform -1 0 8832 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1241_
timestamp 1
transform -1 0 10304 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1
transform 1 0 9660 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1243_
timestamp 1
transform 1 0 8648 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1244_
timestamp 1
transform 1 0 8832 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1
transform -1 0 9660 0 1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1246_
timestamp 1
transform 1 0 8832 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1247_
timestamp 1
transform 1 0 9660 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1248_
timestamp 1
transform -1 0 9660 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1249_
timestamp 1
transform 1 0 9568 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1250_
timestamp 1
transform 1 0 10304 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1251_
timestamp 1
transform 1 0 10028 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1252_
timestamp 1
transform -1 0 10948 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1253_
timestamp 1
transform 1 0 10948 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1254_
timestamp 1
transform 1 0 9016 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1255_
timestamp 1
transform -1 0 10028 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1256_
timestamp 1
transform -1 0 10212 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1257_
timestamp 1
transform -1 0 10396 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1258_
timestamp 1
transform 1 0 9844 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1
transform 1 0 8832 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1260_
timestamp 1
transform 1 0 9200 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1261_
timestamp 1
transform 1 0 9292 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1262_
timestamp 1
transform 1 0 9384 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1263_
timestamp 1
transform 1 0 8648 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1264_
timestamp 1
transform 1 0 8648 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1265_
timestamp 1
transform 1 0 10396 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1266_
timestamp 1
transform 1 0 10304 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1267_
timestamp 1
transform 1 0 10028 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1268_
timestamp 1
transform 1 0 10212 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1269_
timestamp 1
transform 1 0 9384 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1270_
timestamp 1
transform 1 0 11132 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1271_
timestamp 1
transform 1 0 11040 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1272_
timestamp 1
transform 1 0 11132 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1273_
timestamp 1
transform -1 0 11592 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1
transform -1 0 11500 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1
transform 1 0 11776 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1
transform -1 0 12972 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1277_
timestamp 1
transform -1 0 13156 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1278_
timestamp 1
transform 1 0 13156 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1279_
timestamp 1
transform -1 0 13064 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1280_
timestamp 1
transform 1 0 13524 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1281_
timestamp 1
transform 1 0 12696 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1282_
timestamp 1
transform 1 0 12144 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1283_
timestamp 1
transform 1 0 11776 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1284_
timestamp 1
transform 1 0 11408 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1285_
timestamp 1
transform -1 0 13432 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1286_
timestamp 1
transform -1 0 14536 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1287_
timestamp 1
transform 1 0 14076 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1288_
timestamp 1
transform -1 0 14076 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1
transform 1 0 19596 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1290_
timestamp 1
transform 1 0 21252 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _1291_
timestamp 1
transform -1 0 19596 0 1 37536
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _1292_
timestamp 1
transform -1 0 18584 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1293_
timestamp 1
transform 1 0 17204 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1294_
timestamp 1
transform -1 0 17572 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1295_
timestamp 1
transform 1 0 18308 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1296_
timestamp 1
transform -1 0 17940 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1297_
timestamp 1
transform -1 0 19412 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1298_
timestamp 1
transform -1 0 19504 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1299_
timestamp 1
transform 1 0 18676 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1300_
timestamp 1
transform -1 0 19228 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1301_
timestamp 1
transform 1 0 19412 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1302_
timestamp 1
transform -1 0 20240 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1303_
timestamp 1
transform 1 0 19688 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1304_
timestamp 1
transform 1 0 10948 0 -1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1305_
timestamp 1
transform 1 0 12604 0 -1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1306_
timestamp 1
transform -1 0 13984 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1307_
timestamp 1
transform 1 0 11684 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1308_
timestamp 1
transform 1 0 14812 0 1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1309__3
timestamp 1
transform 1 0 19320 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1310__4
timestamp 1
transform 1 0 18308 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1311__5
timestamp 1
transform 1 0 18676 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1312__6
timestamp 1
transform -1 0 17112 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1313__7
timestamp 1
transform -1 0 20240 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1314__8
timestamp 1
transform 1 0 12420 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1315__9
timestamp 1
transform 1 0 10948 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1316__10
timestamp 1
transform 1 0 13156 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1317__11
timestamp 1
transform 1 0 10764 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1318__12
timestamp 1
transform 1 0 9016 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1319__13
timestamp 1
transform -1 0 9200 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1320__14
timestamp 1
transform -1 0 8280 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1321__15
timestamp 1
transform 1 0 8004 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1322__16
timestamp 1
transform -1 0 8648 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1323__17
timestamp 1
transform -1 0 8648 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1324__18
timestamp 1
transform -1 0 9752 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1325__19
timestamp 1
transform 1 0 11040 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1326__20
timestamp 1
transform 1 0 10856 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1327__21
timestamp 1
transform -1 0 13892 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1328__22
timestamp 1
transform -1 0 17112 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1329__23
timestamp 1
transform 1 0 12420 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1330__24
timestamp 1
transform -1 0 22172 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1331__25
timestamp 1
transform -1 0 12328 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1332__26
timestamp 1
transform -1 0 19228 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1333__27
timestamp 1
transform 1 0 16560 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1334__28
timestamp 1
transform -1 0 14444 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1335__29
timestamp 1
transform -1 0 14444 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1336__30
timestamp 1
transform 1 0 12328 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1337__31
timestamp 1
transform -1 0 11316 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1338__32
timestamp 1
transform -1 0 11132 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339__33
timestamp 1
transform -1 0 18952 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1340__34
timestamp 1
transform -1 0 19044 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1341__35
timestamp 1
transform 1 0 16192 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1342__36
timestamp 1
transform -1 0 16836 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1343__37
timestamp 1
transform 1 0 19872 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1344__38
timestamp 1
transform -1 0 20332 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1345__39
timestamp 1
transform -1 0 18952 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1346__40
timestamp 1
transform -1 0 17204 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1347__41
timestamp 1
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1348__42
timestamp 1
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1349__43
timestamp 1
transform -1 0 14996 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1350__44
timestamp 1
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1351__45
timestamp 1
transform -1 0 14628 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1352__46
timestamp 1
transform -1 0 16376 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1353__47
timestamp 1
transform 1 0 14628 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1354__48
timestamp 1
transform -1 0 14444 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1355__49
timestamp 1
transform 1 0 8004 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1356__50
timestamp 1
transform -1 0 14904 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1357__51
timestamp 1
transform 1 0 13524 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1358__52
timestamp 1
transform 1 0 14352 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1359__53
timestamp 1
transform 1 0 17112 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1360__54
timestamp 1
transform 1 0 12604 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1361__55
timestamp 1
transform -1 0 12604 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1362__56
timestamp 1
transform 1 0 11316 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1363__57
timestamp 1
transform -1 0 12236 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1364__58
timestamp 1
transform 1 0 16560 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1365__59
timestamp 1
transform -1 0 18492 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1366__60
timestamp 1
transform -1 0 18124 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1367__61
timestamp 1
transform 1 0 17204 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1368__62
timestamp 1
transform -1 0 16468 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1369__63
timestamp 1
transform 1 0 14076 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1370__64
timestamp 1
transform 1 0 13616 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1371__65
timestamp 1
transform 1 0 14536 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1372__66
timestamp 1
transform -1 0 22264 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1373__67
timestamp 1
transform -1 0 22264 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1374__68
timestamp 1
transform -1 0 22448 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1375__69
timestamp 1
transform -1 0 21620 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1376__70
timestamp 1
transform -1 0 19320 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1377__71
timestamp 1
transform 1 0 20056 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1378__72
timestamp 1
transform -1 0 22080 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1379__73
timestamp 1
transform -1 0 20056 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1380__74
timestamp 1
transform -1 0 13800 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1381__75
timestamp 1
transform 1 0 27140 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1382__76
timestamp 1
transform 1 0 28980 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1383__77
timestamp 1
transform 1 0 26680 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1384__78
timestamp 1
transform 1 0 28612 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1385__79
timestamp 1
transform 1 0 30084 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1386__80
timestamp 1
transform 1 0 29164 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1387__81
timestamp 1
transform -1 0 29440 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1388__82
timestamp 1
transform 1 0 31004 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1389__83
timestamp 1
transform 1 0 31004 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1390__84
timestamp 1
transform -1 0 29716 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1391__85
timestamp 1
transform -1 0 28244 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1392__86
timestamp 1
transform -1 0 27416 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1393__87
timestamp 1
transform -1 0 26772 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1394__88
timestamp 1
transform -1 0 24288 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1395__89
timestamp 1
transform -1 0 28888 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1396__90
timestamp 1
transform 1 0 24288 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1397__91
timestamp 1
transform -1 0 26312 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1398__92
timestamp 1
transform 1 0 27140 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1399__93
timestamp 1
transform -1 0 28520 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1400__94
timestamp 1
transform 1 0 28980 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1401__95
timestamp 1
transform -1 0 27784 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1402__96
timestamp 1
transform 1 0 28612 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1403__97
timestamp 1
transform 1 0 27048 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1404__98
timestamp 1
transform 1 0 29072 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1405__99
timestamp 1
transform 1 0 28980 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1406__100
timestamp 1
transform -1 0 28796 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1407__101
timestamp 1
transform 1 0 28980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1408__102
timestamp 1
transform 1 0 27968 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1409__103
timestamp 1
transform -1 0 26036 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1410__104
timestamp 1
transform -1 0 26772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1411__105
timestamp 1
transform -1 0 26128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1412__106
timestamp 1
transform -1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1413__107
timestamp 1
transform -1 0 22540 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1414__108
timestamp 1
transform 1 0 22356 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1415__109
timestamp 1
transform -1 0 26220 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1416__110
timestamp 1
transform -1 0 25484 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1417__111
timestamp 1
transform 1 0 19596 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1418__112
timestamp 1
transform -1 0 20332 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1419__113
timestamp 1
transform -1 0 19596 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1420__114
timestamp 1
transform -1 0 20424 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1421__115
timestamp 1
transform -1 0 21620 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1422__116
timestamp 1
transform -1 0 19688 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1423__117
timestamp 1
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1424__118
timestamp 1
transform -1 0 19688 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1425__119
timestamp 1
transform -1 0 23552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1426__120
timestamp 1
transform -1 0 24564 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1427__121
timestamp 1
transform -1 0 24564 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1428__122
timestamp 1
transform 1 0 23460 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1429__123
timestamp 1
transform -1 0 22080 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1430__124
timestamp 1
transform 1 0 21436 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1431__125
timestamp 1
transform 1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1432__126
timestamp 1
transform -1 0 22448 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1433__127
timestamp 1
transform 1 0 18308 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1434__128
timestamp 1
transform -1 0 24748 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1435__129
timestamp 1
transform -1 0 23736 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1436__130
timestamp 1
transform 1 0 19596 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1437__131
timestamp 1
transform -1 0 21804 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1438__132
timestamp 1
transform -1 0 23460 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1439__133
timestamp 1
transform -1 0 22356 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1440__134
timestamp 1
transform -1 0 22816 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1441__135
timestamp 1
transform -1 0 20792 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1442__136
timestamp 1
transform -1 0 19688 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1443__137
timestamp 1
transform 1 0 23460 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1444__138
timestamp 1
transform 1 0 23920 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1445__139
timestamp 1
transform -1 0 23920 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1446__140
timestamp 1
transform 1 0 23460 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1447__141
timestamp 1
transform -1 0 21528 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1448__142
timestamp 1
transform 1 0 23368 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1449__143
timestamp 1
transform -1 0 22264 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1450__144
timestamp 1
transform -1 0 20608 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1
transform -1 0 12420 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1
transform 1 0 19228 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1
transform 1 0 18676 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1
transform -1 0 19688 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1
transform 1 0 16744 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1
transform 1 0 20240 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1
transform 1 0 13616 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1
transform 1 0 11224 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1
transform 1 0 13524 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1
transform 1 0 11040 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1461_
timestamp 1
transform 1 0 9292 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1
transform 1 0 8832 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1
transform 1 0 8372 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1
transform 1 0 8372 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1
transform 1 0 8096 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1
transform 1 0 8096 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1
transform 1 0 9384 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1
transform 1 0 11316 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1
transform 1 0 11132 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1
transform 1 0 13524 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1471_
timestamp 1
transform 1 0 16744 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1472_
timestamp 1
transform 1 0 12512 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1473_
timestamp 1
transform 1 0 21804 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1474_
timestamp 1
transform 1 0 11960 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1475_
timestamp 1
transform -1 0 22724 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1476_
timestamp 1
transform -1 0 29348 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1477_
timestamp 1
transform -1 0 28244 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1478_
timestamp 1
transform -1 0 27876 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1479_
timestamp 1
transform -1 0 27876 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1480_
timestamp 1
transform -1 0 26772 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1481_
timestamp 1
transform -1 0 25484 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1482_
timestamp 1
transform -1 0 25300 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1483_
timestamp 1
transform 1 0 21712 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1484_
timestamp 1
transform 1 0 18676 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1485_
timestamp 1
transform 1 0 16836 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1486_
timestamp 1
transform 1 0 14076 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1487_
timestamp 1
transform 1 0 14444 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1488_
timestamp 1
transform 1 0 12512 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1489_
timestamp 1
transform 1 0 10948 0 -1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1490_
timestamp 1
transform 1 0 11132 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1491_
timestamp 1
transform 1 0 18308 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1492_
timestamp 1
transform 1 0 18676 0 -1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1493_
timestamp 1
transform 1 0 16468 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1494_
timestamp 1
transform 1 0 16468 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1495_
timestamp 1
transform 1 0 19596 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1496_
timestamp 1
transform -1 0 20056 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1497_
timestamp 1
transform 1 0 18216 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1498_
timestamp 1
transform 1 0 16836 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1499_
timestamp 1
transform 1 0 15180 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1500_
timestamp 1
transform 1 0 13892 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1501_
timestamp 1
transform 1 0 14168 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1502_
timestamp 1
transform 1 0 16100 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1503_
timestamp 1
transform 1 0 14260 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1504_
timestamp 1
transform 1 0 16100 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1505_
timestamp 1
transform 1 0 14260 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1506_
timestamp 1
transform 1 0 14076 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1507_
timestamp 1
transform 1 0 8280 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1508_
timestamp 1
transform 1 0 14536 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1509_
timestamp 1
transform 1 0 13984 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1510_
timestamp 1
transform 1 0 14628 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1511_
timestamp 1
transform -1 0 17664 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1512_
timestamp 1
transform -1 0 13984 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1513_
timestamp 1
transform 1 0 12236 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1514_
timestamp 1
transform 1 0 11592 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1515_
timestamp 1
transform 1 0 11868 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1516_
timestamp 1
transform 1 0 16836 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1517_
timestamp 1
transform 1 0 17664 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1518_
timestamp 1
transform 1 0 17756 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1519_
timestamp 1
transform 1 0 16468 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1520_
timestamp 1
transform 1 0 16100 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1521_
timestamp 1
transform 1 0 14352 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1522_
timestamp 1
transform 1 0 13892 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1
transform 1 0 15364 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1
transform 1 0 21896 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1
transform 1 0 21252 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1
transform 1 0 21252 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1
transform 1 0 21252 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1
transform 1 0 18952 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1
transform 1 0 20332 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1530_
timestamp 1
transform 1 0 21252 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1
transform 1 0 19688 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1
transform 1 0 13800 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1
transform 1 0 27416 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1534_
timestamp 1
transform -1 0 29440 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1535_
timestamp 1
transform 1 0 26956 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1536_
timestamp 1
transform 1 0 28980 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1537_
timestamp 1
transform 1 0 29900 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1538_
timestamp 1
transform 1 0 29900 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1539_
timestamp 1
transform 1 0 29072 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1540_
timestamp 1
transform -1 0 31372 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1541_
timestamp 1
transform -1 0 30912 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1542_
timestamp 1
transform 1 0 29348 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1543_
timestamp 1
transform 1 0 27876 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1544_
timestamp 1
transform 1 0 27048 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1545_
timestamp 1
transform 1 0 26404 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1546_
timestamp 1
transform 1 0 23920 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1547_
timestamp 1
transform -1 0 28612 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1548_
timestamp 1
transform 1 0 24196 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1549_
timestamp 1
transform 1 0 25944 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1550_
timestamp 1
transform 1 0 27416 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1551_
timestamp 1
transform -1 0 29164 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1552_
timestamp 1
transform -1 0 28888 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1553_
timestamp 1
transform 1 0 27416 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1554_
timestamp 1
transform 1 0 28980 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1555_
timestamp 1
transform 1 0 27324 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1556_
timestamp 1
transform 1 0 28980 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1557_
timestamp 1
transform 1 0 28796 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1558_
timestamp 1
transform 1 0 28428 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1559_
timestamp 1
transform -1 0 28888 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1560_
timestamp 1
transform -1 0 28796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1561_
timestamp 1
transform 1 0 25668 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1562_
timestamp 1
transform 1 0 26404 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1563_
timestamp 1
transform -1 0 25760 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1564_
timestamp 1
transform 1 0 23828 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1565_
timestamp 1
transform 1 0 22172 0 1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1566_
timestamp 1
transform 1 0 22724 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1567_
timestamp 1
transform 1 0 25852 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1568_
timestamp 1
transform 1 0 24380 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1569_
timestamp 1
transform 1 0 19320 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1570_
timestamp 1
transform 1 0 20332 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1571_
timestamp 1
transform 1 0 18768 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1572_
timestamp 1
transform 1 0 20424 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1573_
timestamp 1
transform 1 0 21252 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1574_
timestamp 1
transform 1 0 19136 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1575_
timestamp 1
transform 1 0 21252 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1576_
timestamp 1
transform 1 0 19320 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1577_
timestamp 1
transform 1 0 23092 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1578_
timestamp 1
transform 1 0 23828 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1579_
timestamp 1
transform 1 0 24196 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1580_
timestamp 1
transform 1 0 23828 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1
transform 1 0 21712 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1
transform 1 0 21804 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1
transform 1 0 22172 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1
transform 1 0 22080 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1
transform 1 0 19044 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1
transform 1 0 24564 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1
transform 1 0 22448 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1
transform 1 0 19504 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1
transform 1 0 21252 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1
transform 1 0 22724 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1
transform 1 0 21712 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1
transform 1 0 21896 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1
transform 1 0 20424 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1
transform 1 0 19688 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1
transform 1 0 23828 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1
transform 1 0 24196 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1
transform 1 0 23092 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1
transform 1 0 24196 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1
transform 1 0 21160 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1
transform -1 0 24104 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1
transform 1 0 21896 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1
transform 1 0 20240 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1609_
timestamp 1
transform 1 0 10488 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1610_
timestamp 1
transform 1 0 9108 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1611_
timestamp 1
transform 1 0 8556 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1612_
timestamp 1
transform -1 0 7176 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1613_
timestamp 1
transform -1 0 6808 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1614_
timestamp 1
transform -1 0 13892 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1615_
timestamp 1
transform -1 0 12972 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1616_
timestamp 1
transform -1 0 13524 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1617_
timestamp 1
transform 1 0 11408 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1618_
timestamp 1
transform -1 0 22724 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 21068 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 20976 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1
transform -1 0 17848 0 1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1
transform 1 0 18032 0 -1 19040
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1
transform -1 0 15456 0 1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1
transform 1 0 17112 0 1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1
transform -1 0 23184 0 -1 20128
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1
transform 1 0 25300 0 1 19040
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1
transform 1 0 22264 0 -1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1
transform 1 0 25024 0 -1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1
transform -1 0 15088 0 -1 33184
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1
transform 1 0 16836 0 -1 34272
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1
transform -1 0 15180 0 -1 37536
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1
transform 1 0 16100 0 -1 37536
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1
transform 1 0 22632 0 1 33184
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1
transform 1 0 25116 0 1 34272
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1
transform -1 0 23552 0 -1 38624
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1
transform 1 0 24840 0 -1 37536
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_12  clkload0
timestamp 1
transform 1 0 16100 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_16  clkload1
timestamp 1
transform 1 0 18676 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_12  clkload2
timestamp 1
transform 1 0 14444 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload3
timestamp 1
transform 1 0 17664 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload4
timestamp 1
transform 1 0 22172 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload5
timestamp 1
transform 1 0 24932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload6
timestamp 1
transform 1 0 22264 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_16  clkload7
timestamp 1
transform 1 0 25024 0 1 22304
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_8  clkload8
timestamp 1
transform 1 0 14076 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_16  clkload9
timestamp 1
transform 1 0 16836 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__clkinv_8  clkload10
timestamp 1
transform 1 0 16008 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload11
timestamp 1
transform 1 0 22632 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload12
timestamp 1
transform 1 0 25116 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload13
timestamp 1
transform 1 0 22724 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  clkload14
timestamp 1
transform 1 0 24840 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1
transform 1 0 28428 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1
transform 1 0 27600 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 1
transform 1 0 14720 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1
transform -1 0 14076 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1
transform -1 0 26496 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1
transform 1 0 28152 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1
transform 1 0 21068 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1
transform 1 0 20240 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1
transform -1 0 13064 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1
transform -1 0 19228 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1
transform -1 0 13340 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1
transform 1 0 17204 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1
transform -1 0 14904 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1
transform -1 0 16560 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1
transform -1 0 13432 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1
transform 1 0 12880 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1
transform 1 0 20240 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1
transform -1 0 21068 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1
transform 1 0 20700 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout34
timestamp 1
transform 1 0 20884 0 1 34272
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1
transform -1 0 20608 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 1
transform -1 0 21068 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1
transform -1 0 22172 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1
transform -1 0 21804 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1
transform -1 0 21804 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1
transform -1 0 21620 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1
transform 1 0 18492 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1
transform 1 0 18216 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1
transform 1 0 23184 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1
transform 1 0 17848 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1
transform -1 0 24012 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 1
transform 1 0 22724 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1
transform 1 0 23368 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1
transform -1 0 23552 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1
transform 1 0 23092 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1
transform -1 0 15548 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 1
transform -1 0 16468 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 1
transform 1 0 19872 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 1
transform -1 0 23644 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 1
transform 1 0 23368 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 1
transform -1 0 23644 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1
transform 1 0 16836 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 1
transform -1 0 15272 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp 1
transform -1 0 16468 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1
transform -1 0 22172 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1
transform -1 0 20608 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout61
timestamp 1
transform -1 0 21344 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout62
timestamp 1
transform 1 0 21252 0 1 41888
box -38 -48 958 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636968456
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636968456
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636968456
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1636968456
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636968456
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636968456
transform 1 0 30084 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333
timestamp 1
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636968456
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636968456
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636968456
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636968456
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1
transform 1 0 30820 0 -1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636968456
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636968456
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636968456
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636968456
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636968456
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636968456
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636968456
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636968456
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636968456
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636968456
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636968456
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636968456
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636968456
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636968456
transform 1 0 30084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 1
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636968456
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636968456
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636968456
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636968456
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1636968456
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1636968456
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1636968456
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1636968456
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636968456
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636968456
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636968456
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636968456
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636968456
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1636968456
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1636968456
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1636968456
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1
transform 1 0 30820 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636968456
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636968456
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636968456
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1636968456
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1636968456
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1636968456
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1636968456
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636968456
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1636968456
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1636968456
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1636968456
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636968456
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636968456
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1636968456
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1636968456
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636968456
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636968456
transform 1 0 30084 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_333
timestamp 1
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636968456
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636968456
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636968456
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636968456
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636968456
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636968456
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1636968456
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1636968456
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1636968456
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636968456
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1636968456
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1636968456
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1636968456
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636968456
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1636968456
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1636968456
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636968456
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1636968456
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1636968456
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1636968456
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1
transform 1 0 30820 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636968456
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636968456
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636968456
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636968456
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636968456
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1636968456
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1636968456
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1636968456
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1636968456
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1636968456
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1636968456
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1636968456
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1636968456
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1636968456
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1636968456
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1636968456
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636968456
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636968456
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1636968456
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636968456
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1636968456
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1636968456
transform 1 0 30084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 1
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636968456
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636968456
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636968456
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636968456
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636968456
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1636968456
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1636968456
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1636968456
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1636968456
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1636968456
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1636968456
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1636968456
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1636968456
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1636968456
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1636968456
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1636968456
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1636968456
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1636968456
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1636968456
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1636968456
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636968456
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1636968456
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1636968456
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1
transform 1 0 30820 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636968456
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1636968456
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1636968456
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1636968456
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1636968456
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1636968456
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1636968456
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1636968456
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1636968456
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1636968456
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1636968456
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1636968456
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1636968456
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1636968456
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1636968456
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1636968456
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636968456
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1636968456
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1636968456
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1636968456
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1636968456
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1636968456
transform 1 0 30084 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_333
timestamp 1
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636968456
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636968456
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636968456
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1636968456
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1636968456
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1636968456
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1636968456
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1636968456
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1636968456
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1636968456
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636968456
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1636968456
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1636968456
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1636968456
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1636968456
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1636968456
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1636968456
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1636968456
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636968456
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636968456
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1636968456
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1636968456
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1
transform 1 0 30820 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636968456
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636968456
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636968456
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1636968456
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1636968456
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1636968456
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1636968456
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1636968456
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1636968456
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636968456
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1636968456
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1636968456
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1636968456
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636968456
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636968456
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1636968456
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1636968456
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1636968456
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1636968456
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1636968456
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1636968456
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1636968456
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1636968456
transform 1 0 30084 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_333
timestamp 1
transform 1 0 31188 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636968456
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636968456
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636968456
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1636968456
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636968456
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1636968456
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1636968456
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1636968456
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1636968456
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1636968456
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1636968456
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1636968456
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1636968456
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1636968456
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1636968456
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1636968456
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636968456
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1636968456
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1636968456
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1636968456
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1636968456
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1636968456
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1636968456
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1636968456
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1
transform 1 0 30820 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636968456
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636968456
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636968456
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636968456
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1636968456
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1636968456
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636968456
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1636968456
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1636968456
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1636968456
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636968456
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636968456
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1636968456
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1636968456
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636968456
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1636968456
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1636968456
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1636968456
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1
transform 1 0 23092 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636968456
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1636968456
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1636968456
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1636968456
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636968456
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1636968456
transform 1 0 30084 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 1
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636968456
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636968456
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636968456
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1636968456
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1636968456
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1636968456
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1636968456
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1636968456
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1636968456
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1636968456
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1636968456
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636968456
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1636968456
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1636968456
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1636968456
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1
transform 1 0 20516 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1636968456
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1636968456
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1636968456
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1636968456
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1636968456
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1636968456
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1636968456
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1636968456
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1
transform 1 0 30820 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636968456
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636968456
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636968456
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1636968456
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1636968456
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1636968456
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1636968456
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1636968456
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1636968456
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1636968456
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1636968456
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1636968456
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1636968456
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1636968456
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1636968456
transform 1 0 19780 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1636968456
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1636968456
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1636968456
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1636968456
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1636968456
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1636968456
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1636968456
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1636968456
transform 1 0 30084 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_333
timestamp 1
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636968456
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1636968456
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1636968456
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636968456
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1636968456
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1636968456
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1636968456
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636968456
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1636968456
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1636968456
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1636968456
transform 1 0 14260 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1
transform 1 0 15364 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1636968456
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1636968456
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1636968456
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1636968456
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1
transform 1 0 20516 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1636968456
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1636968456
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1636968456
transform 1 0 23460 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1636968456
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1
transform 1 0 25668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1636968456
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1636968456
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1636968456
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1636968456
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1
transform 1 0 30820 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636968456
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636968456
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636968456
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636968456
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1636968456
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1636968456
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1636968456
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1636968456
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1636968456
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1636968456
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1
transform 1 0 12788 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1636968456
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1636968456
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1636968456
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1636968456
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1
transform 1 0 17940 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1636968456
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1636968456
transform 1 0 19780 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1636968456
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1636968456
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1
transform 1 0 23092 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1636968456
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1636968456
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1636968456
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1636968456
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1636968456
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1636968456
transform 1 0 30084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_333
timestamp 1
transform 1 0 31188 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636968456
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1636968456
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1636968456
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1636968456
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636968456
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1636968456
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1636968456
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1636968456
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1
transform 1 0 10212 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636968456
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1636968456
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1636968456
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1636968456
transform 1 0 14260 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1636968456
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1636968456
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1636968456
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1636968456
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1
transform 1 0 20516 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636968456
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1636968456
transform 1 0 22356 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1636968456
transform 1 0 23460 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1636968456
transform 1 0 24564 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1
transform 1 0 25668 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1636968456
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1636968456
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1636968456
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1636968456
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1
transform 1 0 30820 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636968456
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1636968456
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1636968456
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1636968456
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1636968456
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1636968456
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636968456
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636968456
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1636968456
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1636968456
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1636968456
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1636968456
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1636968456
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1636968456
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1
transform 1 0 17940 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1636968456
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1636968456
transform 1 0 19780 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1636968456
transform 1 0 20884 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1636968456
transform 1 0 21988 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1
transform 1 0 23092 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1636968456
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1636968456
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1636968456
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1636968456
transform 1 0 27140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1
transform 1 0 28244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1636968456
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1636968456
transform 1 0 30084 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_333
timestamp 1
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636968456
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1636968456
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1636968456
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1636968456
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1636968456
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1636968456
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1636968456
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1636968456
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636968456
transform 1 0 10948 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636968456
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1636968456
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1636968456
transform 1 0 14260 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_161
timestamp 1
transform 1 0 15364 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_169
timestamp 1
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_177
timestamp 1
transform 1 0 16836 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1636968456
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1636968456
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1636968456
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1
transform 1 0 20516 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1636968456
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1636968456
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1636968456
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1636968456
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1636968456
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1636968456
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1636968456
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1636968456
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1
transform 1 0 30820 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636968456
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1636968456
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1636968456
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1636968456
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1636968456
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1636968456
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1636968456
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1636968456
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1636968456
transform 1 0 10580 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1636968456
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1636968456
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_153
timestamp 1
transform 1 0 14628 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_175
timestamp 1
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1636968456
transform 1 0 18676 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1636968456
transform 1 0 19780 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1636968456
transform 1 0 20884 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1636968456
transform 1 0 21988 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1
transform 1 0 23092 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1636968456
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1636968456
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1636968456
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1636968456
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1
transform 1 0 28244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1636968456
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1636968456
transform 1 0 30084 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_333
timestamp 1
transform 1 0 31188 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636968456
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1636968456
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1636968456
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1636968456
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1636968456
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1636968456
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1636968456
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1636968456
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1636968456
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1636968456
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1636968456
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1636968456
transform 1 0 14260 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_161
timestamp 1
transform 1 0 15364 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_208
timestamp 1636968456
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp 1
transform 1 0 20792 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1636968456
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1636968456
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1636968456
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1636968456
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1636968456
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1636968456
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1636968456
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1636968456
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1
transform 1 0 30820 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636968456
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1636968456
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636968456
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1636968456
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1636968456
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1636968456
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1636968456
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1636968456
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1636968456
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1636968456
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1636968456
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_153
timestamp 1
transform 1 0 14628 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_159
timestamp 1
transform 1 0 15180 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_167
timestamp 1
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_177
timestamp 1
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_200
timestamp 1636968456
transform 1 0 18952 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_212
timestamp 1636968456
transform 1 0 20056 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_224
timestamp 1636968456
transform 1 0 21160 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_236
timestamp 1636968456
transform 1 0 22264 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_248
timestamp 1
transform 1 0 23368 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1636968456
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_265
timestamp 1
transform 1 0 24932 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_271
timestamp 1
transform 1 0 25484 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_280
timestamp 1636968456
transform 1 0 26312 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_292
timestamp 1636968456
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_304
timestamp 1
transform 1 0 28520 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1636968456
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1636968456
transform 1 0 30084 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_333
timestamp 1
transform 1 0 31188 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636968456
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1636968456
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1636968456
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1636968456
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1636968456
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1636968456
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1636968456
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1636968456
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636968456
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1636968456
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_137
timestamp 1
transform 1 0 13156 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_145
timestamp 1
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_180
timestamp 1
transform 1 0 17112 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_196
timestamp 1
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_208
timestamp 1636968456
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 1
transform 1 0 20792 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1636968456
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1636968456
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_249
timestamp 1
transform 1 0 23460 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1
transform 1 0 26036 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_298
timestamp 1636968456
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_310
timestamp 1636968456
transform 1 0 29072 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_322
timestamp 1636968456
transform 1 0 30176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_334
timestamp 1
transform 1 0 31280 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636968456
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636968456
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1636968456
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1636968456
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1636968456
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1636968456
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636968456
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1636968456
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1636968456
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1636968456
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_203
timestamp 1636968456
transform 1 0 19228 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_215
timestamp 1636968456
transform 1 0 20332 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_227
timestamp 1636968456
transform 1 0 21436 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_239
timestamp 1
transform 1 0 22540 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_243
timestamp 1
transform 1 0 22908 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_278
timestamp 1
transform 1 0 26128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_285
timestamp 1
transform 1 0 26772 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_294
timestamp 1636968456
transform 1 0 27600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1
transform 1 0 28704 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1636968456
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1636968456
transform 1 0 30084 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_333
timestamp 1
transform 1 0 31188 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636968456
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1636968456
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1636968456
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1636968456
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1636968456
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1636968456
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1636968456
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1636968456
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1636968456
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1636968456
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_137
timestamp 1
transform 1 0 13156 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_145
timestamp 1
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_154
timestamp 1
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_183
timestamp 1
transform 1 0 17388 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_187
timestamp 1
transform 1 0 17756 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_194
timestamp 1
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_215
timestamp 1
transform 1 0 20332 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1
transform 1 0 21252 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_233
timestamp 1
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_238
timestamp 1636968456
transform 1 0 22448 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_250
timestamp 1
transform 1 0 23552 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_257
timestamp 1
transform 1 0 24196 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_270
timestamp 1
transform 1 0 25392 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1636968456
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1636968456
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1636968456
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1636968456
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1
transform 1 0 30820 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636968456
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1636968456
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1636968456
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1636968456
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1636968456
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1636968456
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1636968456
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1636968456
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1636968456
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1636968456
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636968456
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_153
timestamp 1
transform 1 0 14628 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_157
timestamp 1
transform 1 0 14996 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_168
timestamp 1
transform 1 0 16008 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_179
timestamp 1
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_187
timestamp 1
transform 1 0 17756 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_197
timestamp 1
transform 1 0 18676 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_205
timestamp 1
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_223
timestamp 1
transform 1 0 21068 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1
transform 1 0 23552 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1636968456
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_292
timestamp 1636968456
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_304
timestamp 1
transform 1 0 28520 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1636968456
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1636968456
transform 1 0 30084 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_333
timestamp 1
transform 1 0 31188 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1636968456
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1636968456
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1636968456
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1636968456
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1636968456
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1636968456
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1636968456
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1636968456
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1636968456
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1636968456
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_149
timestamp 1
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_157
timestamp 1
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_169
timestamp 1
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_174
timestamp 1636968456
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_189
timestamp 1636968456
transform 1 0 17940 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_201
timestamp 1
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_213
timestamp 1
transform 1 0 20148 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_222
timestamp 1
transform 1 0 20976 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_241
timestamp 1636968456
transform 1 0 22724 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_253
timestamp 1636968456
transform 1 0 23828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_265
timestamp 1636968456
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 1
transform 1 0 26036 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_307
timestamp 1636968456
transform 1 0 28796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_319
timestamp 1636968456
transform 1 0 29900 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_331
timestamp 1
transform 1 0 31004 0 -1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636968456
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636968456
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1636968456
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1636968456
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1636968456
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1636968456
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1636968456
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1636968456
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1636968456
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1636968456
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1636968456
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_153
timestamp 1
transform 1 0 14628 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_174
timestamp 1
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_208
timestamp 1
transform 1 0 19688 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_216
timestamp 1
transform 1 0 20424 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_224
timestamp 1
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_229
timestamp 1636968456
transform 1 0 21620 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_241
timestamp 1
transform 1 0 22724 0 1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_269
timestamp 1636968456
transform 1 0 25300 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_281
timestamp 1
transform 1 0 26404 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_312
timestamp 1636968456
transform 1 0 29256 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_324
timestamp 1
transform 1 0 30360 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_332
timestamp 1
transform 1 0 31096 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1636968456
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1636968456
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1636968456
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1636968456
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1636968456
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1636968456
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1636968456
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1636968456
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636968456
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1636968456
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1636968456
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_149
timestamp 1
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_157
timestamp 1
transform 1 0 14996 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1
transform 1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_176
timestamp 1
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_184
timestamp 1
transform 1 0 17480 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_188
timestamp 1
transform 1 0 17848 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_200
timestamp 1636968456
transform 1 0 18952 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_212
timestamp 1
transform 1 0 20056 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_216
timestamp 1
transform 1 0 20424 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1
transform 1 0 20976 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_233
timestamp 1
transform 1 0 21988 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_237
timestamp 1
transform 1 0 22356 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_246
timestamp 1
transform 1 0 23184 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_254
timestamp 1
transform 1 0 23920 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_281
timestamp 1
transform 1 0 26404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_285
timestamp 1
transform 1 0 26772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_289
timestamp 1
transform 1 0 27140 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_301
timestamp 1636968456
transform 1 0 28244 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_313
timestamp 1636968456
transform 1 0 29348 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_325
timestamp 1
transform 1 0 30452 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_333
timestamp 1
transform 1 0 31188 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1636968456
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1636968456
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1636968456
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1636968456
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1636968456
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1636968456
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1636968456
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1636968456
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1636968456
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1636968456
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1
transform 1 0 13524 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_169
timestamp 1636968456
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_181
timestamp 1
transform 1 0 17204 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_187
timestamp 1
transform 1 0 17756 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_191
timestamp 1
transform 1 0 18124 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_197
timestamp 1
transform 1 0 18676 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_210
timestamp 1
transform 1 0 19872 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_269
timestamp 1
transform 1 0 25300 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_291
timestamp 1636968456
transform 1 0 27324 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_303
timestamp 1
transform 1 0 28428 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1636968456
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1636968456
transform 1 0 30084 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_333
timestamp 1
transform 1 0 31188 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636968456
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1636968456
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1636968456
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1636968456
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1636968456
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1636968456
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1636968456
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1636968456
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1636968456
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1636968456
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1636968456
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_149
timestamp 1
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_158
timestamp 1
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_203
timestamp 1
transform 1 0 19228 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 1
transform 1 0 20792 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_233
timestamp 1
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_248
timestamp 1
transform 1 0 23368 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_256
timestamp 1
transform 1 0 24104 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_261
timestamp 1
transform 1 0 24564 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_265
timestamp 1
transform 1 0 24932 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 1
transform 1 0 26128 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1636968456
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1636968456
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_305
timestamp 1
transform 1 0 28612 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_309
timestamp 1
transform 1 0 28980 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_313
timestamp 1636968456
transform 1 0 29348 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_325
timestamp 1
transform 1 0 30452 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_333
timestamp 1
transform 1 0 31188 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1636968456
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1636968456
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1636968456
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1636968456
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1636968456
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1636968456
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1636968456
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1636968456
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1636968456
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1636968456
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_141
timestamp 1
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_149
timestamp 1
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_160
timestamp 1
transform 1 0 15272 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1636968456
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1636968456
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1636968456
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1636968456
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_277
timestamp 1
transform 1 0 26036 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_285
timestamp 1
transform 1 0 26772 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_325
timestamp 1
transform 1 0 30452 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_333
timestamp 1
transform 1 0 31188 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636968456
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1636968456
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1636968456
transform 1 0 3036 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1636968456
transform 1 0 4140 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1
transform 1 0 5244 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1636968456
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1636968456
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1636968456
transform 1 0 8004 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1636968456
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1
transform 1 0 10212 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1
transform 1 0 10764 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1636968456
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1636968456
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1636968456
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1636968456
transform 1 0 14260 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_161
timestamp 1
transform 1 0 15364 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_169
timestamp 1
transform 1 0 16100 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_189
timestamp 1
transform 1 0 17940 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_201
timestamp 1
transform 1 0 19044 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_208
timestamp 1636968456
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 1
transform 1 0 20792 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_225
timestamp 1
transform 1 0 21252 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_248
timestamp 1
transform 1 0 23368 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_261
timestamp 1
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_288
timestamp 1
transform 1 0 27048 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_321
timestamp 1636968456
transform 1 0 30084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_333
timestamp 1
transform 1 0 31188 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1636968456
transform 1 0 828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1636968456
transform 1 0 1932 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1636968456
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1636968456
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1636968456
transform 1 0 5428 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1636968456
transform 1 0 6532 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1
transform 1 0 7636 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1
transform 1 0 8188 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1636968456
transform 1 0 8372 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1636968456
transform 1 0 9476 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1636968456
transform 1 0 10580 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1636968456
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1
transform 1 0 12788 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1
transform 1 0 13340 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_141
timestamp 1
transform 1 0 13524 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_171
timestamp 1
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_184
timestamp 1
transform 1 0 17480 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1
transform 1 0 18308 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_197
timestamp 1
transform 1 0 18676 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_208
timestamp 1
transform 1 0 19688 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_285
timestamp 1
transform 1 0 26772 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_290
timestamp 1
transform 1 0 27232 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_298
timestamp 1
transform 1 0 27968 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_304
timestamp 1
transform 1 0 28520 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1636968456
transform 1 0 28980 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1636968456
transform 1 0 30084 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_333
timestamp 1
transform 1 0 31188 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1636968456
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1636968456
transform 1 0 1932 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1636968456
transform 1 0 3036 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1636968456
transform 1 0 4140 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1
transform 1 0 5244 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1636968456
transform 1 0 5796 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1636968456
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1636968456
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1636968456
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1
transform 1 0 10212 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1
transform 1 0 10764 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1636968456
transform 1 0 10948 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1636968456
transform 1 0 12052 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1636968456
transform 1 0 13156 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_149
timestamp 1
transform 1 0 14260 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_160
timestamp 1
transform 1 0 15272 0 -1 20128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1636968456
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_181
timestamp 1
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_185
timestamp 1
transform 1 0 17572 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_233
timestamp 1
transform 1 0 21988 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_246
timestamp 1
transform 1 0 23184 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_250
timestamp 1
transform 1 0 23552 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_258
timestamp 1
transform 1 0 24288 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_262
timestamp 1
transform 1 0 24656 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_270
timestamp 1
transform 1 0 25392 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_297
timestamp 1636968456
transform 1 0 27876 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_309
timestamp 1636968456
transform 1 0 28980 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_321
timestamp 1636968456
transform 1 0 30084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_333
timestamp 1
transform 1 0 31188 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1636968456
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1636968456
transform 1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1636968456
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1636968456
transform 1 0 4324 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1636968456
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1636968456
transform 1 0 6532 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1
transform 1 0 7636 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1636968456
transform 1 0 8372 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1636968456
transform 1 0 9476 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1636968456
transform 1 0 10580 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1636968456
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1
transform 1 0 12788 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1
transform 1 0 13340 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1636968456
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1636968456
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_165
timestamp 1
transform 1 0 15732 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_171
timestamp 1636968456
transform 1 0 16284 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_183
timestamp 1
transform 1 0 17388 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1
transform 1 0 18492 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_216
timestamp 1636968456
transform 1 0 20424 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_228
timestamp 1
transform 1 0 21528 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_232
timestamp 1
transform 1 0 21896 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_244
timestamp 1
transform 1 0 23000 0 1 20128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1636968456
transform 1 0 23828 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_265
timestamp 1
transform 1 0 24932 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_274
timestamp 1
transform 1 0 25760 0 1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_280
timestamp 1636968456
transform 1 0 26312 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_292
timestamp 1
transform 1 0 27416 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_298
timestamp 1
transform 1 0 27968 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_302
timestamp 1
transform 1 0 28336 0 1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1636968456
transform 1 0 28980 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1636968456
transform 1 0 30084 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_333
timestamp 1
transform 1 0 31188 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1636968456
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1636968456
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1636968456
transform 1 0 3036 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1636968456
transform 1 0 4140 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1
transform 1 0 5244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1636968456
transform 1 0 5796 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1636968456
transform 1 0 6900 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1636968456
transform 1 0 8004 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1636968456
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1
transform 1 0 10212 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1636968456
transform 1 0 10948 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1636968456
transform 1 0 12052 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1636968456
transform 1 0 13156 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_149
timestamp 1
transform 1 0 14260 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_157
timestamp 1
transform 1 0 14996 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_190
timestamp 1636968456
transform 1 0 18032 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_202
timestamp 1636968456
transform 1 0 19136 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_214
timestamp 1
transform 1 0 20240 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1
transform 1 0 20976 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_225
timestamp 1
transform 1 0 21252 0 -1 21216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_234
timestamp 1636968456
transform 1 0 22080 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_246
timestamp 1636968456
transform 1 0 23184 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_258
timestamp 1
transform 1 0 24288 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_268
timestamp 1636968456
transform 1 0 25208 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_281
timestamp 1
transform 1 0 26404 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_289
timestamp 1
transform 1 0 27140 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_323
timestamp 1636968456
transform 1 0 30268 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636968456
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1636968456
transform 1 0 1932 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1636968456
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1636968456
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1636968456
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1636968456
transform 1 0 6532 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1
transform 1 0 7636 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1
transform 1 0 8188 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1636968456
transform 1 0 8372 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1636968456
transform 1 0 9476 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1636968456
transform 1 0 10580 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1636968456
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1
transform 1 0 12788 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1
transform 1 0 13340 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_149
timestamp 1
transform 1 0 14260 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_156
timestamp 1636968456
transform 1 0 14904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_168
timestamp 1
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_173
timestamp 1
transform 1 0 16468 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1
transform 1 0 18308 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_218
timestamp 1
transform 1 0 20608 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_229
timestamp 1
transform 1 0 21620 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1
transform 1 0 23644 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_269
timestamp 1
transform 1 0 25300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_283
timestamp 1
transform 1 0 26588 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1
transform 1 0 28796 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_312
timestamp 1636968456
transform 1 0 29256 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_324
timestamp 1
transform 1 0 30360 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_332
timestamp 1
transform 1 0 31096 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1636968456
transform 1 0 828 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1636968456
transform 1 0 1932 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1636968456
transform 1 0 3036 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1636968456
transform 1 0 4140 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1
transform 1 0 5244 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1
transform 1 0 5612 0 -1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1636968456
transform 1 0 5796 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1636968456
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1636968456
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1636968456
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1
transform 1 0 10212 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1
transform 1 0 10764 0 -1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1636968456
transform 1 0 10948 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_125
timestamp 1
transform 1 0 12052 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_129
timestamp 1
transform 1 0 12420 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1
transform 1 0 15916 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_177
timestamp 1
transform 1 0 16836 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_197
timestamp 1
transform 1 0 18676 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1
transform 1 0 20976 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_241
timestamp 1
transform 1 0 22724 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_261
timestamp 1
transform 1 0 24564 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_295
timestamp 1
transform 1 0 27692 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_301
timestamp 1
transform 1 0 28244 0 -1 22304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_319
timestamp 1636968456
transform 1 0 29900 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_331
timestamp 1
transform 1 0 31004 0 -1 22304
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1636968456
transform 1 0 828 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1636968456
transform 1 0 1932 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1636968456
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1636968456
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1636968456
transform 1 0 5428 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1636968456
transform 1 0 6532 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1
transform 1 0 7636 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1
transform 1 0 8188 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1636968456
transform 1 0 8372 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1636968456
transform 1 0 9476 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1636968456
transform 1 0 10580 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_121
timestamp 1
transform 1 0 11684 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_129
timestamp 1
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_134
timestamp 1
transform 1 0 12880 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_168
timestamp 1
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_178
timestamp 1
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 1
transform 1 0 18400 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_202
timestamp 1
transform 1 0 19136 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_245
timestamp 1
transform 1 0 23092 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1
transform 1 0 23644 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_298
timestamp 1
transform 1 0 27968 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1
transform 1 0 28796 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1636968456
transform 1 0 28980 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1636968456
transform 1 0 30084 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_333
timestamp 1
transform 1 0 31188 0 1 22304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1636968456
transform 1 0 828 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1636968456
transform 1 0 1932 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1636968456
transform 1 0 3036 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1636968456
transform 1 0 4140 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1
transform 1 0 5244 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1
transform 1 0 5612 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1636968456
transform 1 0 5796 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1636968456
transform 1 0 6900 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1636968456
transform 1 0 8004 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1636968456
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1
transform 1 0 10212 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1
transform 1 0 10764 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1636968456
transform 1 0 10948 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_125
timestamp 1
transform 1 0 12052 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_164
timestamp 1
transform 1 0 15640 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_169
timestamp 1
transform 1 0 16100 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_213
timestamp 1
transform 1 0 20148 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_217
timestamp 1
transform 1 0 20516 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1
transform 1 0 21068 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_228
timestamp 1
transform 1 0 21528 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_235
timestamp 1
transform 1 0 22172 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_250
timestamp 1
transform 1 0 23552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_261
timestamp 1
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_265
timestamp 1
transform 1 0 24932 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1
transform 1 0 26036 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_284
timestamp 1
transform 1 0 26680 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_290
timestamp 1
transform 1 0 27232 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_307
timestamp 1636968456
transform 1 0 28796 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_319
timestamp 1636968456
transform 1 0 29900 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_331
timestamp 1
transform 1 0 31004 0 -1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1636968456
transform 1 0 828 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1636968456
transform 1 0 1932 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1
transform 1 0 3036 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1636968456
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1636968456
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1636968456
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1636968456
transform 1 0 6532 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1
transform 1 0 7636 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1
transform 1 0 8188 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1636968456
transform 1 0 8372 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1636968456
transform 1 0 9476 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1636968456
transform 1 0 10580 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_121
timestamp 1
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_127
timestamp 1
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_131
timestamp 1
transform 1 0 12604 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_141
timestamp 1
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_170
timestamp 1
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_183
timestamp 1
transform 1 0 17388 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_191
timestamp 1
transform 1 0 18124 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1
transform 1 0 18492 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_205
timestamp 1
transform 1 0 19412 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_213
timestamp 1
transform 1 0 20148 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_217
timestamp 1636968456
transform 1 0 20516 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_229
timestamp 1636968456
transform 1 0 21620 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_241
timestamp 1
transform 1 0 22724 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_249
timestamp 1
transform 1 0 23460 0 1 23392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1636968456
transform 1 0 23828 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1636968456
transform 1 0 24932 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_277
timestamp 1
transform 1 0 26036 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_285
timestamp 1
transform 1 0 26772 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_289
timestamp 1
transform 1 0 27140 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_325
timestamp 1
transform 1 0 30452 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_333
timestamp 1
transform 1 0 31188 0 1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1636968456
transform 1 0 828 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1636968456
transform 1 0 1932 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1636968456
transform 1 0 3036 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1636968456
transform 1 0 4140 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1
transform 1 0 5244 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1
transform 1 0 5612 0 -1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1636968456
transform 1 0 5796 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1636968456
transform 1 0 6900 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1636968456
transform 1 0 8004 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1636968456
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1
transform 1 0 10212 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1
transform 1 0 10764 0 -1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1636968456
transform 1 0 10948 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_125
timestamp 1
transform 1 0 12052 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_133
timestamp 1
transform 1 0 12788 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_144
timestamp 1
transform 1 0 13800 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_156
timestamp 1
transform 1 0 14904 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_169
timestamp 1
transform 1 0 16100 0 -1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_175
timestamp 1636968456
transform 1 0 16652 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_187
timestamp 1636968456
transform 1 0 17756 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_199
timestamp 1636968456
transform 1 0 18860 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_211
timestamp 1
transform 1 0 19964 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_220
timestamp 1
transform 1 0 20792 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_238
timestamp 1
transform 1 0 22448 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_284
timestamp 1
transform 1 0 26680 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_292
timestamp 1
transform 1 0 27416 0 -1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1636968456
transform 1 0 28612 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1636968456
transform 1 0 29716 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1
transform 1 0 30820 0 -1 24480
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1636968456
transform 1 0 828 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1636968456
transform 1 0 1932 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1
transform 1 0 3036 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1636968456
transform 1 0 3220 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1636968456
transform 1 0 4324 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1636968456
transform 1 0 5428 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1636968456
transform 1 0 6532 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1
transform 1 0 7636 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1
transform 1 0 8188 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1636968456
transform 1 0 8372 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1636968456
transform 1 0 9476 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_109
timestamp 1
transform 1 0 10580 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_136
timestamp 1
transform 1 0 13064 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_149
timestamp 1
transform 1 0 14260 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_169
timestamp 1636968456
transform 1 0 16100 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_181
timestamp 1
transform 1 0 17204 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1
transform 1 0 18308 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_197
timestamp 1
transform 1 0 18676 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_213
timestamp 1
transform 1 0 20148 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_230
timestamp 1
transform 1 0 21712 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1
transform 1 0 23644 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_258
timestamp 1
transform 1 0 24288 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_291
timestamp 1
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1636968456
transform 1 0 28980 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1636968456
transform 1 0 30084 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_333
timestamp 1
transform 1 0 31188 0 1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1636968456
transform 1 0 828 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1636968456
transform 1 0 1932 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1636968456
transform 1 0 3036 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1636968456
transform 1 0 4140 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1
transform 1 0 5244 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1
transform 1 0 5612 0 -1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1636968456
transform 1 0 5796 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1636968456
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1636968456
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1636968456
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1
transform 1 0 10212 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1
transform 1 0 10764 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_113
timestamp 1
transform 1 0 10948 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_121
timestamp 1
transform 1 0 11684 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_139
timestamp 1
transform 1 0 13340 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_189
timestamp 1
transform 1 0 17940 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_209
timestamp 1
transform 1 0 19780 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_218
timestamp 1
transform 1 0 20608 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_225
timestamp 1
transform 1 0 21252 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_236
timestamp 1
transform 1 0 22264 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_258
timestamp 1
transform 1 0 24288 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_263
timestamp 1
transform 1 0 24748 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_274
timestamp 1
transform 1 0 25760 0 -1 25568
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1636968456
transform 1 0 26404 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_296
timestamp 1636968456
transform 1 0 27784 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_308
timestamp 1636968456
transform 1 0 28888 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_320
timestamp 1636968456
transform 1 0 29992 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_332
timestamp 1
transform 1 0 31096 0 -1 25568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1636968456
transform 1 0 828 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1636968456
transform 1 0 1932 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1
transform 1 0 3036 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1636968456
transform 1 0 3220 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1636968456
transform 1 0 4324 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1636968456
transform 1 0 5428 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1636968456
transform 1 0 6532 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1
transform 1 0 7636 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1
transform 1 0 8188 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1636968456
transform 1 0 8372 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1636968456
transform 1 0 9476 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1636968456
transform 1 0 10580 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_121
timestamp 1
transform 1 0 11684 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_127
timestamp 1
transform 1 0 12236 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_133
timestamp 1
transform 1 0 12788 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_149
timestamp 1
transform 1 0 14260 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_169
timestamp 1
transform 1 0 16100 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_200
timestamp 1
transform 1 0 18952 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_216
timestamp 1636968456
transform 1 0 20424 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_228
timestamp 1636968456
transform 1 0 21528 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_240
timestamp 1636968456
transform 1 0 22632 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1636968456
transform 1 0 23828 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1636968456
transform 1 0 24932 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1636968456
transform 1 0 26036 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_289
timestamp 1
transform 1 0 27140 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1
transform 1 0 28244 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1
transform 1 0 28796 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1636968456
transform 1 0 28980 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1636968456
transform 1 0 30084 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_333
timestamp 1
transform 1 0 31188 0 1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636968456
transform 1 0 828 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1636968456
transform 1 0 1932 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1636968456
transform 1 0 3036 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1636968456
transform 1 0 4140 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1
transform 1 0 5244 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1
transform 1 0 5612 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1636968456
transform 1 0 5796 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1636968456
transform 1 0 6900 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1636968456
transform 1 0 8004 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1636968456
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1
transform 1 0 10212 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1
transform 1 0 10764 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1636968456
transform 1 0 10948 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_125
timestamp 1
transform 1 0 12052 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_152
timestamp 1
transform 1 0 14536 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 1
transform 1 0 15548 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1
transform 1 0 15916 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_169
timestamp 1
transform 1 0 16100 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_173
timestamp 1
transform 1 0 16468 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_177
timestamp 1
transform 1 0 16836 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_213
timestamp 1
transform 1 0 20148 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1
transform 1 0 20976 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_228
timestamp 1
transform 1 0 21528 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_246
timestamp 1
transform 1 0 23184 0 -1 26656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_257
timestamp 1636968456
transform 1 0 24196 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_269
timestamp 1
transform 1 0 25300 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_277
timestamp 1
transform 1 0 26036 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_289
timestamp 1
transform 1 0 27140 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_293
timestamp 1
transform 1 0 27508 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_303
timestamp 1636968456
transform 1 0 28428 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_315
timestamp 1636968456
transform 1 0 29532 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_327
timestamp 1
transform 1 0 30636 0 -1 26656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1636968456
transform 1 0 828 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1636968456
transform 1 0 1932 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1
transform 1 0 3036 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1636968456
transform 1 0 3220 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1636968456
transform 1 0 4324 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1636968456
transform 1 0 5428 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1636968456
transform 1 0 6532 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1
transform 1 0 7636 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1
transform 1 0 8188 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1636968456
transform 1 0 8372 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1636968456
transform 1 0 9476 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_109
timestamp 1
transform 1 0 10580 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_132
timestamp 1
transform 1 0 12696 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_141
timestamp 1
transform 1 0 13524 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_147
timestamp 1
transform 1 0 14076 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_155
timestamp 1636968456
transform 1 0 14812 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_167
timestamp 1
transform 1 0 15916 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_175
timestamp 1
transform 1 0 16652 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1
transform 1 0 18400 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_248
timestamp 1
transform 1 0 23368 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_269
timestamp 1
transform 1 0 25300 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_289
timestamp 1
transform 1 0 27140 0 1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_312
timestamp 1636968456
transform 1 0 29256 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_324
timestamp 1
transform 1 0 30360 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_332
timestamp 1
transform 1 0 31096 0 1 26656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1636968456
transform 1 0 828 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1636968456
transform 1 0 1932 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1636968456
transform 1 0 3036 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1636968456
transform 1 0 4140 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1
transform 1 0 5244 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1
transform 1 0 5612 0 -1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1636968456
transform 1 0 5796 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1636968456
transform 1 0 6900 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1636968456
transform 1 0 8004 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1636968456
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1
transform 1 0 10212 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1
transform 1 0 10764 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_113
timestamp 1
transform 1 0 10948 0 -1 27744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_129
timestamp 1636968456
transform 1 0 12420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_141
timestamp 1
transform 1 0 13524 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_154
timestamp 1
transform 1 0 14720 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_160
timestamp 1
transform 1 0 15272 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1
transform 1 0 15916 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_169
timestamp 1
transform 1 0 16100 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_178
timestamp 1
transform 1 0 16928 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_186
timestamp 1
transform 1 0 17664 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1
transform 1 0 21068 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_225
timestamp 1
transform 1 0 21252 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_234
timestamp 1
transform 1 0 22080 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_243
timestamp 1
transform 1 0 22908 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_258
timestamp 1
transform 1 0 24288 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_270
timestamp 1
transform 1 0 25392 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_290
timestamp 1
transform 1 0 27232 0 -1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_311
timestamp 1636968456
transform 1 0 29164 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_323
timestamp 1636968456
transform 1 0 30268 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1636968456
transform 1 0 828 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1636968456
transform 1 0 1932 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1
transform 1 0 3036 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1636968456
transform 1 0 3220 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1636968456
transform 1 0 4324 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1636968456
transform 1 0 5428 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1636968456
transform 1 0 6532 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1
transform 1 0 7636 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1
transform 1 0 8188 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1636968456
transform 1 0 8372 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1636968456
transform 1 0 9476 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_109
timestamp 1
transform 1 0 10580 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_120
timestamp 1
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_126
timestamp 1636968456
transform 1 0 12144 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1
transform 1 0 13248 0 1 27744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_145
timestamp 1636968456
transform 1 0 13892 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_157
timestamp 1
transform 1 0 14996 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_190
timestamp 1
transform 1 0 18032 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_197
timestamp 1
transform 1 0 18676 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_201
timestamp 1
transform 1 0 19044 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_222
timestamp 1636968456
transform 1 0 20976 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_237
timestamp 1636968456
transform 1 0 22356 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_249
timestamp 1
transform 1 0 23460 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_267
timestamp 1
transform 1 0 25116 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_271
timestamp 1
transform 1 0 25484 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1636968456
transform 1 0 26036 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_289
timestamp 1
transform 1 0 27140 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_302
timestamp 1
transform 1 0 28336 0 1 27744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1636968456
transform 1 0 28980 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1636968456
transform 1 0 30084 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_333
timestamp 1
transform 1 0 31188 0 1 27744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1636968456
transform 1 0 828 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1636968456
transform 1 0 1932 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1636968456
transform 1 0 3036 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1636968456
transform 1 0 4140 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1
transform 1 0 5244 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1
transform 1 0 5612 0 -1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1636968456
transform 1 0 5796 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1636968456
transform 1 0 6900 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1636968456
transform 1 0 8004 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1636968456
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1
transform 1 0 10212 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1
transform 1 0 10764 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_161
timestamp 1
transform 1 0 15364 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_169
timestamp 1
transform 1 0 16100 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_175
timestamp 1
transform 1 0 16652 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_179
timestamp 1
transform 1 0 17020 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_185
timestamp 1
transform 1 0 17572 0 -1 28832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_191
timestamp 1636968456
transform 1 0 18124 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_203
timestamp 1
transform 1 0 19228 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_209
timestamp 1
transform 1 0 19780 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_216
timestamp 1
transform 1 0 20424 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_222
timestamp 1
transform 1 0 20976 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_233
timestamp 1
transform 1 0 21988 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_242
timestamp 1
transform 1 0 22816 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_261
timestamp 1
transform 1 0 24564 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_290
timestamp 1
transform 1 0 27232 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_294
timestamp 1
transform 1 0 27600 0 -1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_311
timestamp 1636968456
transform 1 0 29164 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_323
timestamp 1636968456
transform 1 0 30268 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1636968456
transform 1 0 828 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1636968456
transform 1 0 1932 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1
transform 1 0 3036 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1636968456
transform 1 0 3220 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1636968456
transform 1 0 4324 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1636968456
transform 1 0 5428 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1636968456
transform 1 0 6532 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1
transform 1 0 7636 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1
transform 1 0 8188 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1636968456
transform 1 0 8372 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1636968456
transform 1 0 9476 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_109
timestamp 1
transform 1 0 10580 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_113
timestamp 1
transform 1 0 10948 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_117
timestamp 1
transform 1 0 11316 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_122
timestamp 1
transform 1 0 11776 0 1 28832
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_162
timestamp 1636968456
transform 1 0 15456 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_174
timestamp 1
transform 1 0 16560 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_178
timestamp 1
transform 1 0 16928 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_185
timestamp 1
transform 1 0 17572 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_197
timestamp 1
transform 1 0 18676 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_203
timestamp 1
transform 1 0 19228 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_214
timestamp 1
transform 1 0 20240 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_258
timestamp 1
transform 1 0 24288 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_266
timestamp 1
transform 1 0 25024 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_279
timestamp 1636968456
transform 1 0 26220 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_291
timestamp 1
transform 1 0 27324 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_295
timestamp 1
transform 1 0 27692 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_304
timestamp 1
transform 1 0 28520 0 1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1636968456
transform 1 0 28980 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1636968456
transform 1 0 30084 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_333
timestamp 1
transform 1 0 31188 0 1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1636968456
transform 1 0 828 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1636968456
transform 1 0 1932 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1636968456
transform 1 0 3036 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1636968456
transform 1 0 4140 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1
transform 1 0 5244 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1
transform 1 0 5612 0 -1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1636968456
transform 1 0 5796 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1636968456
transform 1 0 6900 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1636968456
transform 1 0 8004 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1636968456
transform 1 0 9108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1
transform 1 0 10212 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1
transform 1 0 10764 0 -1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1636968456
transform 1 0 10948 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1636968456
transform 1 0 12052 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_137
timestamp 1
transform 1 0 13156 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_145
timestamp 1
transform 1 0 13892 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_164
timestamp 1
transform 1 0 15640 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_178
timestamp 1
transform 1 0 16928 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_199
timestamp 1
transform 1 0 18860 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_216
timestamp 1
transform 1 0 20424 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_220
timestamp 1
transform 1 0 20792 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_225
timestamp 1
transform 1 0 21252 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_242
timestamp 1
transform 1 0 22816 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_246
timestamp 1
transform 1 0 23184 0 -1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_254
timestamp 1636968456
transform 1 0 23920 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_266
timestamp 1
transform 1 0 25024 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1
transform 1 0 25668 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1
transform 1 0 26220 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_288
timestamp 1
transform 1 0 27048 0 -1 29920
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_306
timestamp 1636968456
transform 1 0 28704 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_318
timestamp 1636968456
transform 1 0 29808 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_330
timestamp 1
transform 1 0 30912 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_334
timestamp 1
transform 1 0 31280 0 -1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1636968456
transform 1 0 828 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1636968456
transform 1 0 1932 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1
transform 1 0 3036 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1636968456
transform 1 0 3220 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1636968456
transform 1 0 4324 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1636968456
transform 1 0 5428 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1636968456
transform 1 0 6532 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1
transform 1 0 7636 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1
transform 1 0 8188 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_85
timestamp 1
transform 1 0 8372 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_91
timestamp 1
transform 1 0 8924 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_130
timestamp 1
transform 1 0 12512 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_138
timestamp 1
transform 1 0 13248 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_141
timestamp 1
transform 1 0 13524 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_147
timestamp 1
transform 1 0 14076 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_151
timestamp 1
transform 1 0 14444 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_159
timestamp 1
transform 1 0 15180 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_168
timestamp 1
transform 1 0 16008 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1
transform 1 0 17940 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1
transform 1 0 18492 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_197
timestamp 1
transform 1 0 18676 0 1 29920
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_204
timestamp 1636968456
transform 1 0 19320 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_216
timestamp 1636968456
transform 1 0 20424 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_228
timestamp 1636968456
transform 1 0 21528 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_240
timestamp 1636968456
transform 1 0 22632 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_269
timestamp 1636968456
transform 1 0 25300 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_281
timestamp 1
transform 1 0 26404 0 1 29920
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1636968456
transform 1 0 28980 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1636968456
transform 1 0 30084 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_333
timestamp 1
transform 1 0 31188 0 1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1636968456
transform 1 0 828 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1636968456
transform 1 0 1932 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1636968456
transform 1 0 3036 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1636968456
transform 1 0 4140 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1
transform 1 0 5244 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1
transform 1 0 5612 0 -1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1636968456
transform 1 0 5796 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1636968456
transform 1 0 6900 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_81
timestamp 1
transform 1 0 8004 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_89
timestamp 1
transform 1 0 8740 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_106
timestamp 1
transform 1 0 10304 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_134
timestamp 1
transform 1 0 12880 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_146
timestamp 1
transform 1 0 13984 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_169
timestamp 1
transform 1 0 16100 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_179
timestamp 1
transform 1 0 17020 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_186
timestamp 1
transform 1 0 17664 0 -1 31008
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_203
timestamp 1636968456
transform 1 0 19228 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_215
timestamp 1
transform 1 0 20332 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1
transform 1 0 21068 0 -1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1636968456
transform 1 0 21252 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_237
timestamp 1
transform 1 0 22356 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_245
timestamp 1
transform 1 0 23092 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1
transform 1 0 25668 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1
transform 1 0 26220 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_289
timestamp 1
transform 1 0 27140 0 -1 31008
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_300
timestamp 1636968456
transform 1 0 28152 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_312
timestamp 1636968456
transform 1 0 29256 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_324
timestamp 1
transform 1 0 30360 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_332
timestamp 1
transform 1 0 31096 0 -1 31008
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1636968456
transform 1 0 828 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1636968456
transform 1 0 1932 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1
transform 1 0 3036 0 1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1636968456
transform 1 0 3220 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1636968456
transform 1 0 4324 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1636968456
transform 1 0 5428 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1636968456
transform 1 0 6532 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1
transform 1 0 7636 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1
transform 1 0 8188 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_85
timestamp 1
transform 1 0 8372 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_104
timestamp 1
transform 1 0 10120 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_110
timestamp 1
transform 1 0 10672 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_119
timestamp 1
transform 1 0 11500 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_129
timestamp 1
transform 1 0 12420 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_157
timestamp 1
transform 1 0 14996 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_172
timestamp 1
transform 1 0 16376 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_176
timestamp 1
transform 1 0 16744 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_183
timestamp 1
transform 1 0 17388 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_194
timestamp 1
transform 1 0 18400 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_213
timestamp 1
transform 1 0 20148 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_235
timestamp 1
transform 1 0 22172 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_245
timestamp 1
transform 1 0 23092 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_253
timestamp 1
transform 1 0 23828 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_273
timestamp 1
transform 1 0 25668 0 1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_295
timestamp 1636968456
transform 1 0 27692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1
transform 1 0 28796 0 1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1636968456
transform 1 0 28980 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1636968456
transform 1 0 30084 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_333
timestamp 1
transform 1 0 31188 0 1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1636968456
transform 1 0 828 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1636968456
transform 1 0 1932 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1636968456
transform 1 0 3036 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1636968456
transform 1 0 4140 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1
transform 1 0 5244 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1
transform 1 0 5612 0 -1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1636968456
transform 1 0 5796 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1636968456
transform 1 0 6900 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_81
timestamp 1
transform 1 0 8004 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_89
timestamp 1
transform 1 0 8740 0 -1 32096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_94
timestamp 1636968456
transform 1 0 9200 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_106
timestamp 1
transform 1 0 10304 0 -1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1636968456
transform 1 0 10948 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_125
timestamp 1
transform 1 0 12052 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_152
timestamp 1
transform 1 0 14536 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1
transform 1 0 15916 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_169
timestamp 1
transform 1 0 16100 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_183
timestamp 1
transform 1 0 17388 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_190
timestamp 1
transform 1 0 18032 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_198
timestamp 1
transform 1 0 18768 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_203
timestamp 1
transform 1 0 19228 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_222
timestamp 1
transform 1 0 20976 0 -1 32096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_263
timestamp 1636968456
transform 1 0 24748 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_275
timestamp 1
transform 1 0 25852 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1
transform 1 0 26220 0 -1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_284
timestamp 1636968456
transform 1 0 26680 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_296
timestamp 1
transform 1 0 27784 0 -1 32096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_314
timestamp 1636968456
transform 1 0 29440 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_326
timestamp 1
transform 1 0 30544 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_334
timestamp 1
transform 1 0 31280 0 -1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1636968456
transform 1 0 828 0 1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1636968456
transform 1 0 1932 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1
transform 1 0 3036 0 1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1636968456
transform 1 0 3220 0 1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1636968456
transform 1 0 4324 0 1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1636968456
transform 1 0 5428 0 1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1636968456
transform 1 0 6532 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1
transform 1 0 7636 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1
transform 1 0 8188 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_85
timestamp 1
transform 1 0 8372 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_93
timestamp 1
transform 1 0 9108 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_112
timestamp 1
transform 1 0 10856 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_120
timestamp 1
transform 1 0 11592 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_136
timestamp 1
transform 1 0 13064 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_141
timestamp 1
transform 1 0 13524 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_147
timestamp 1
transform 1 0 14076 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_174
timestamp 1
transform 1 0 16560 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1
transform 1 0 17940 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1
transform 1 0 18492 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_197
timestamp 1
transform 1 0 18676 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_205
timestamp 1
transform 1 0 19412 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_210
timestamp 1
transform 1 0 19872 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_231
timestamp 1
transform 1 0 21804 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_249
timestamp 1
transform 1 0 23460 0 1 32096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1636968456
transform 1 0 23828 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_265
timestamp 1
transform 1 0 24932 0 1 32096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_271
timestamp 1636968456
transform 1 0 25484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_283
timestamp 1
transform 1 0 26588 0 1 32096
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_312
timestamp 1636968456
transform 1 0 29256 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_324
timestamp 1
transform 1 0 30360 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_332
timestamp 1
transform 1 0 31096 0 1 32096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1636968456
transform 1 0 828 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1636968456
transform 1 0 1932 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1636968456
transform 1 0 3036 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1636968456
transform 1 0 4140 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1
transform 1 0 5244 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1
transform 1 0 5612 0 -1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1636968456
transform 1 0 5796 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1636968456
transform 1 0 6900 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_81
timestamp 1
transform 1 0 8004 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_87
timestamp 1
transform 1 0 8556 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_113
timestamp 1
transform 1 0 10948 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_124
timestamp 1
transform 1 0 11960 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_144
timestamp 1
transform 1 0 13800 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_158
timestamp 1
transform 1 0 15088 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_163
timestamp 1
transform 1 0 15548 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1
transform 1 0 15916 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_169
timestamp 1
transform 1 0 16100 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_193
timestamp 1
transform 1 0 18308 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_204
timestamp 1
transform 1 0 19320 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_213
timestamp 1
transform 1 0 20148 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_221
timestamp 1
transform 1 0 20884 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_225
timestamp 1
transform 1 0 21252 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_233
timestamp 1
transform 1 0 21988 0 -1 33184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_240
timestamp 1636968456
transform 1 0 22632 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_252
timestamp 1
transform 1 0 23736 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_256
timestamp 1
transform 1 0 24104 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_260
timestamp 1
transform 1 0 24472 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_269
timestamp 1
transform 1 0 25300 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1
transform 1 0 26220 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_288
timestamp 1
transform 1 0 27048 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_292
timestamp 1
transform 1 0 27416 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_299
timestamp 1
transform 1 0 28060 0 -1 33184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_318
timestamp 1636968456
transform 1 0 29808 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_330
timestamp 1
transform 1 0 30912 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_334
timestamp 1
transform 1 0 31280 0 -1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1636968456
transform 1 0 828 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1636968456
transform 1 0 1932 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1
transform 1 0 3036 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1636968456
transform 1 0 3220 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1636968456
transform 1 0 4324 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1636968456
transform 1 0 5428 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1636968456
transform 1 0 6532 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1
transform 1 0 7636 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1
transform 1 0 8188 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_85
timestamp 1
transform 1 0 8372 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_93
timestamp 1
transform 1 0 9108 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_99
timestamp 1
transform 1 0 9660 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_105
timestamp 1
transform 1 0 10212 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_135
timestamp 1
transform 1 0 12972 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1
transform 1 0 13340 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_141
timestamp 1
transform 1 0 13524 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_160
timestamp 1
transform 1 0 15272 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_168
timestamp 1
transform 1 0 16008 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_194
timestamp 1
transform 1 0 18400 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_202
timestamp 1
transform 1 0 19136 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_210
timestamp 1
transform 1 0 19872 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_238
timestamp 1
transform 1 0 22448 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1
transform 1 0 23644 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_262
timestamp 1
transform 1 0 24656 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_266
timestamp 1
transform 1 0 25024 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_292
timestamp 1
transform 1 0 27416 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_298
timestamp 1
transform 1 0 27968 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1
transform 1 0 28796 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1636968456
transform 1 0 28980 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1636968456
transform 1 0 30084 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_333
timestamp 1
transform 1 0 31188 0 1 33184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1636968456
transform 1 0 828 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1636968456
transform 1 0 1932 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1636968456
transform 1 0 3036 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1636968456
transform 1 0 4140 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1
transform 1 0 5244 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1
transform 1 0 5612 0 -1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1636968456
transform 1 0 5796 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1636968456
transform 1 0 6900 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_81
timestamp 1
transform 1 0 8004 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_89
timestamp 1
transform 1 0 8740 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_103
timestamp 1
transform 1 0 10028 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1
transform 1 0 10764 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_113
timestamp 1
transform 1 0 10948 0 -1 34272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_120
timestamp 1636968456
transform 1 0 11592 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_132
timestamp 1
transform 1 0 12696 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1
transform 1 0 15916 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_169
timestamp 1
transform 1 0 16100 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_188
timestamp 1
transform 1 0 17848 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_202
timestamp 1
transform 1 0 19136 0 -1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_210
timestamp 1636968456
transform 1 0 19872 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_222
timestamp 1
transform 1 0 20976 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_234
timestamp 1
transform 1 0 22080 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_254
timestamp 1
transform 1 0 23920 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_260
timestamp 1
transform 1 0 24472 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_298
timestamp 1
transform 1 0 27968 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_304
timestamp 1
transform 1 0 28520 0 -1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1636968456
transform 1 0 828 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1636968456
transform 1 0 1932 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1
transform 1 0 3036 0 1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1636968456
transform 1 0 3220 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1636968456
transform 1 0 4324 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1636968456
transform 1 0 5428 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1636968456
transform 1 0 6532 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_77
timestamp 1
transform 1 0 7636 0 1 34272
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_108
timestamp 1636968456
transform 1 0 10488 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_120
timestamp 1
transform 1 0 11592 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_128
timestamp 1
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_141
timestamp 1
transform 1 0 13524 0 1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_179
timestamp 1636968456
transform 1 0 17020 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_191
timestamp 1
transform 1 0 18124 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_217
timestamp 1
transform 1 0 20516 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_235
timestamp 1
transform 1 0 22172 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_259
timestamp 1
transform 1 0 24380 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_278
timestamp 1
transform 1 0 26128 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_303
timestamp 1
transform 1 0 28428 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_325
timestamp 1
transform 1 0 30452 0 1 34272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1636968456
transform 1 0 828 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1636968456
transform 1 0 1932 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1636968456
transform 1 0 3036 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1636968456
transform 1 0 4140 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1
transform 1 0 5244 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1
transform 1 0 5612 0 -1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1636968456
transform 1 0 5796 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1636968456
transform 1 0 6900 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1636968456
transform 1 0 8004 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_93
timestamp 1
transform 1 0 9108 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_97
timestamp 1
transform 1 0 9476 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_107
timestamp 1
transform 1 0 10396 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1
transform 1 0 10764 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_113
timestamp 1
transform 1 0 10948 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_117
timestamp 1
transform 1 0 11316 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_158
timestamp 1
transform 1 0 15088 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_166
timestamp 1
transform 1 0 15824 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_175
timestamp 1
transform 1 0 16652 0 -1 35360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_180
timestamp 1636968456
transform 1 0 17112 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_192
timestamp 1
transform 1 0 18216 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_202
timestamp 1
transform 1 0 19136 0 -1 35360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_211
timestamp 1636968456
transform 1 0 19964 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1
transform 1 0 21068 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_225
timestamp 1
transform 1 0 21252 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_236
timestamp 1
transform 1 0 22264 0 -1 35360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_247
timestamp 1636968456
transform 1 0 23276 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_259
timestamp 1
transform 1 0 24380 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_264
timestamp 1
transform 1 0 24840 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_271
timestamp 1
transform 1 0 25484 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1
transform 1 0 26220 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_281
timestamp 1
transform 1 0 26404 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_324
timestamp 1
transform 1 0 30360 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_333
timestamp 1
transform 1 0 31188 0 -1 35360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1636968456
transform 1 0 828 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1636968456
transform 1 0 1932 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1
transform 1 0 3036 0 1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1636968456
transform 1 0 3220 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1636968456
transform 1 0 4324 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1636968456
transform 1 0 5428 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1636968456
transform 1 0 6532 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1
transform 1 0 7636 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1
transform 1 0 8188 0 1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1636968456
transform 1 0 8372 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_105
timestamp 1
transform 1 0 10212 0 1 35360
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_146
timestamp 1636968456
transform 1 0 13984 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_158
timestamp 1
transform 1 0 15088 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_192
timestamp 1
transform 1 0 18216 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_197
timestamp 1
transform 1 0 18676 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_203
timestamp 1
transform 1 0 19228 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_211
timestamp 1
transform 1 0 19964 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_247
timestamp 1
transform 1 0 23276 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1
transform 1 0 23644 0 1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_256
timestamp 1636968456
transform 1 0 24104 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_268
timestamp 1636968456
transform 1 0 25208 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_280
timestamp 1636968456
transform 1 0 26312 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_292
timestamp 1
transform 1 0 27416 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_304
timestamp 1
transform 1 0 28520 0 1 35360
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1636968456
transform 1 0 28980 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1636968456
transform 1 0 30084 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_333
timestamp 1
transform 1 0 31188 0 1 35360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1636968456
transform 1 0 828 0 -1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1636968456
transform 1 0 1932 0 -1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1636968456
transform 1 0 3036 0 -1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1636968456
transform 1 0 4140 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1
transform 1 0 5244 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1
transform 1 0 5612 0 -1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1636968456
transform 1 0 5796 0 -1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1636968456
transform 1 0 6900 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_81
timestamp 1
transform 1 0 8004 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_89
timestamp 1
transform 1 0 8740 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_100
timestamp 1
transform 1 0 9752 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1
transform 1 0 10764 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_113
timestamp 1
transform 1 0 10948 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_121
timestamp 1
transform 1 0 11684 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_129
timestamp 1
transform 1 0 12420 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_140
timestamp 1
transform 1 0 13432 0 -1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_154
timestamp 1636968456
transform 1 0 14720 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_166
timestamp 1
transform 1 0 15824 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_181
timestamp 1
transform 1 0 17204 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_197
timestamp 1
transform 1 0 18676 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_205
timestamp 1
transform 1 0 19412 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_219
timestamp 1
transform 1 0 20700 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1
transform 1 0 21068 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_229
timestamp 1
transform 1 0 21620 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_241
timestamp 1
transform 1 0 22724 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_245
timestamp 1
transform 1 0 23092 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_254
timestamp 1
transform 1 0 23920 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_271
timestamp 1
transform 1 0 25484 0 -1 36448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_290
timestamp 1636968456
transform 1 0 27232 0 -1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_302
timestamp 1636968456
transform 1 0 28336 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_314
timestamp 1
transform 1 0 29440 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_333
timestamp 1
transform 1 0 31188 0 -1 36448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1636968456
transform 1 0 828 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1636968456
transform 1 0 1932 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1
transform 1 0 3036 0 1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1636968456
transform 1 0 3220 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1636968456
transform 1 0 4324 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1636968456
transform 1 0 5428 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1636968456
transform 1 0 6532 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_77
timestamp 1
transform 1 0 7636 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_101
timestamp 1
transform 1 0 9844 0 1 36448
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_120
timestamp 1636968456
transform 1 0 11592 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_132
timestamp 1
transform 1 0 12696 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_148
timestamp 1
transform 1 0 14168 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_161
timestamp 1
transform 1 0 15364 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_176
timestamp 1
transform 1 0 16744 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_184
timestamp 1
transform 1 0 17480 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_206
timestamp 1
transform 1 0 19504 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_235
timestamp 1
transform 1 0 22172 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_243
timestamp 1
transform 1 0 22908 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_253
timestamp 1
transform 1 0 23828 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_300
timestamp 1
transform 1 0 28152 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_309
timestamp 1
transform 1 0 28980 0 1 36448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1636968456
transform 1 0 828 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1636968456
transform 1 0 1932 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1636968456
transform 1 0 3036 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1636968456
transform 1 0 4140 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1
transform 1 0 5244 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1
transform 1 0 5612 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1636968456
transform 1 0 5796 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1636968456
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_81
timestamp 1
transform 1 0 8004 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_89
timestamp 1
transform 1 0 8740 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1
transform 1 0 10764 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1636968456
transform 1 0 10948 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1636968456
transform 1 0 12052 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_137
timestamp 1
transform 1 0 13156 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_159
timestamp 1
transform 1 0 15180 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_180
timestamp 1636968456
transform 1 0 17112 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_197
timestamp 1
transform 1 0 18676 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_253
timestamp 1
transform 1 0 23828 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_275
timestamp 1
transform 1 0 25852 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1
transform 1 0 26220 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_295
timestamp 1
transform 1 0 27692 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_299
timestamp 1
transform 1 0 28060 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1636968456
transform 1 0 828 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1636968456
transform 1 0 1932 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1
transform 1 0 3036 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1636968456
transform 1 0 3220 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1636968456
transform 1 0 4324 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1636968456
transform 1 0 5428 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1636968456
transform 1 0 6532 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1
transform 1 0 7636 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1
transform 1 0 8188 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_85
timestamp 1
transform 1 0 8372 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_93
timestamp 1
transform 1 0 9108 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_108
timestamp 1
transform 1 0 10488 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_138
timestamp 1
transform 1 0 13248 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_190
timestamp 1
transform 1 0 18032 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_207
timestamp 1
transform 1 0 19596 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_223
timestamp 1
transform 1 0 21068 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_234
timestamp 1
transform 1 0 22080 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_253
timestamp 1
transform 1 0 23828 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_261
timestamp 1
transform 1 0 24564 0 1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_270
timestamp 1636968456
transform 1 0 25392 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_282
timestamp 1636968456
transform 1 0 26496 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_294
timestamp 1636968456
transform 1 0 27600 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_306
timestamp 1
transform 1 0 28704 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_309
timestamp 1
transform 1 0 28980 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_326
timestamp 1
transform 1 0 30544 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1636968456
transform 1 0 828 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1636968456
transform 1 0 1932 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1636968456
transform 1 0 3036 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1636968456
transform 1 0 4140 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1
transform 1 0 5244 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1
transform 1 0 5612 0 -1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1636968456
transform 1 0 5796 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1636968456
transform 1 0 6900 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_81
timestamp 1
transform 1 0 8004 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_106
timestamp 1
transform 1 0 10304 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_113
timestamp 1
transform 1 0 10948 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_159
timestamp 1
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_166
timestamp 1
transform 1 0 15824 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_191
timestamp 1
transform 1 0 18124 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_205
timestamp 1
transform 1 0 19412 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_225
timestamp 1
transform 1 0 21252 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_233
timestamp 1
transform 1 0 21988 0 -1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_255
timestamp 1636968456
transform 1 0 24012 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_267
timestamp 1636968456
transform 1 0 25116 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1
transform 1 0 26220 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_281
timestamp 1
transform 1 0 26404 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_287
timestamp 1
transform 1 0 26956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_304
timestamp 1
transform 1 0 28520 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_310
timestamp 1
transform 1 0 29072 0 -1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_314
timestamp 1636968456
transform 1 0 29440 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_326
timestamp 1
transform 1 0 30544 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_334
timestamp 1
transform 1 0 31280 0 -1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1636968456
transform 1 0 828 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1636968456
transform 1 0 1932 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1
transform 1 0 3036 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1636968456
transform 1 0 3220 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1636968456
transform 1 0 4324 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1636968456
transform 1 0 5428 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1636968456
transform 1 0 6532 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1
transform 1 0 7636 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1
transform 1 0 8188 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_88
timestamp 1
transform 1 0 8648 0 1 38624
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_107
timestamp 1636968456
transform 1 0 10396 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_119
timestamp 1
transform 1 0 11500 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_125
timestamp 1
transform 1 0 12052 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_131
timestamp 1
transform 1 0 12604 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1
transform 1 0 13340 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1636968456
transform 1 0 13524 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_153
timestamp 1
transform 1 0 14628 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_161
timestamp 1
transform 1 0 15364 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_168
timestamp 1
transform 1 0 16008 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_185
timestamp 1
transform 1 0 17572 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_193
timestamp 1
transform 1 0 18308 0 1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1636968456
transform 1 0 18676 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_218
timestamp 1636968456
transform 1 0 20608 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_230
timestamp 1636968456
transform 1 0 21712 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_242
timestamp 1
transform 1 0 22816 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_250
timestamp 1
transform 1 0 23552 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_253
timestamp 1
transform 1 0 23828 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_261
timestamp 1
transform 1 0 24564 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_309
timestamp 1
transform 1 0 28980 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_318
timestamp 1
transform 1 0 29808 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_325
timestamp 1
transform 1 0 30452 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_333
timestamp 1
transform 1 0 31188 0 1 38624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1636968456
transform 1 0 828 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1636968456
transform 1 0 1932 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1636968456
transform 1 0 3036 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1636968456
transform 1 0 4140 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1
transform 1 0 5244 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1
transform 1 0 5612 0 -1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1636968456
transform 1 0 5796 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1636968456
transform 1 0 6900 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1636968456
transform 1 0 8004 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_93
timestamp 1
transform 1 0 9108 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_97
timestamp 1
transform 1 0 9476 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_106
timestamp 1
transform 1 0 10304 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_113
timestamp 1
transform 1 0 10948 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_124
timestamp 1
transform 1 0 11960 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_141
timestamp 1
transform 1 0 13524 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_145
timestamp 1
transform 1 0 13892 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_154
timestamp 1
transform 1 0 14720 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_166
timestamp 1
transform 1 0 15824 0 -1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1636968456
transform 1 0 16100 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1636968456
transform 1 0 17204 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_193
timestamp 1
transform 1 0 18308 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_206
timestamp 1
transform 1 0 19504 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_212
timestamp 1
transform 1 0 20056 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_288
timestamp 1
transform 1 0 27048 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_292
timestamp 1
transform 1 0 27416 0 -1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1636968456
transform 1 0 828 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1636968456
transform 1 0 1932 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1
transform 1 0 3036 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1636968456
transform 1 0 3220 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1636968456
transform 1 0 4324 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1636968456
transform 1 0 5428 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1636968456
transform 1 0 6532 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1
transform 1 0 7636 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1
transform 1 0 8188 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_98
timestamp 1
transform 1 0 9568 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_108
timestamp 1
transform 1 0 10488 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_130
timestamp 1
transform 1 0 12512 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_157
timestamp 1
transform 1 0 14996 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_168
timestamp 1
transform 1 0 16008 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_177
timestamp 1
transform 1 0 16836 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_183
timestamp 1
transform 1 0 17388 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_191
timestamp 1
transform 1 0 18124 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_221
timestamp 1
transform 1 0 20884 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_236
timestamp 1
transform 1 0 22264 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_253
timestamp 1
transform 1 0 23828 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_257
timestamp 1
transform 1 0 24196 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_261
timestamp 1
transform 1 0 24564 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_282
timestamp 1
transform 1 0 26496 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_295
timestamp 1
transform 1 0 27692 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_309
timestamp 1
transform 1 0 28980 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_317
timestamp 1
transform 1 0 29716 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_334
timestamp 1
transform 1 0 31280 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1636968456
transform 1 0 828 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1636968456
transform 1 0 1932 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1636968456
transform 1 0 3036 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1636968456
transform 1 0 4140 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1
transform 1 0 5244 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1
transform 1 0 5612 0 -1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1636968456
transform 1 0 5796 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1636968456
transform 1 0 6900 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_81
timestamp 1
transform 1 0 8004 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_98
timestamp 1
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_130
timestamp 1
transform 1 0 12512 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_139
timestamp 1
transform 1 0 13340 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_166
timestamp 1
transform 1 0 15824 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_169
timestamp 1
transform 1 0 16100 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_191
timestamp 1
transform 1 0 18124 0 -1 40800
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_203
timestamp 1636968456
transform 1 0 19228 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_215
timestamp 1
transform 1 0 20332 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1
transform 1 0 21068 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_230
timestamp 1
transform 1 0 21712 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_254
timestamp 1
transform 1 0 23920 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_258
timestamp 1
transform 1 0 24288 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_268
timestamp 1
transform 1 0 25208 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_274
timestamp 1
transform 1 0 25760 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_278
timestamp 1
transform 1 0 26128 0 -1 40800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_286
timestamp 1636968456
transform 1 0 26864 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_298
timestamp 1
transform 1 0 27968 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_306
timestamp 1
transform 1 0 28704 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_314
timestamp 1
transform 1 0 29440 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_334
timestamp 1
transform 1 0 31280 0 -1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1636968456
transform 1 0 828 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1636968456
transform 1 0 1932 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1
transform 1 0 3036 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1636968456
transform 1 0 3220 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1636968456
transform 1 0 4324 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1636968456
transform 1 0 5428 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1636968456
transform 1 0 6532 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1
transform 1 0 7636 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1
transform 1 0 8188 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_110
timestamp 1
transform 1 0 10672 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_138
timestamp 1
transform 1 0 13248 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_141
timestamp 1
transform 1 0 13524 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_147
timestamp 1
transform 1 0 14076 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_151
timestamp 1
transform 1 0 14444 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_177
timestamp 1
transform 1 0 16836 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_181
timestamp 1
transform 1 0 17204 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_197
timestamp 1
transform 1 0 18676 0 1 40800
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 1636968456
transform 1 0 20884 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_236
timestamp 1
transform 1 0 22264 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_240
timestamp 1
transform 1 0 22632 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_250
timestamp 1
transform 1 0 23552 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_253
timestamp 1
transform 1 0 23828 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_270
timestamp 1
transform 1 0 25392 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_287
timestamp 1
transform 1 0 26956 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_313
timestamp 1
transform 1 0 29348 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_330
timestamp 1
transform 1 0 30912 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_334
timestamp 1
transform 1 0 31280 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1636968456
transform 1 0 828 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1636968456
transform 1 0 1932 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1636968456
transform 1 0 3036 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1636968456
transform 1 0 4140 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1
transform 1 0 5244 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1
transform 1 0 5612 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1636968456
transform 1 0 5796 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1636968456
transform 1 0 6900 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1636968456
transform 1 0 8004 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_93
timestamp 1
transform 1 0 9108 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_107
timestamp 1
transform 1 0 10396 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1
transform 1 0 10764 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1636968456
transform 1 0 10948 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_125
timestamp 1
transform 1 0 12052 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_137
timestamp 1
transform 1 0 13156 0 -1 41888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_146
timestamp 1636968456
transform 1 0 13984 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_158
timestamp 1
transform 1 0 15088 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_166
timestamp 1
transform 1 0 15824 0 -1 41888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1636968456
transform 1 0 16100 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_181
timestamp 1
transform 1 0 17204 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_187
timestamp 1
transform 1 0 17756 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_192
timestamp 1636968456
transform 1 0 18216 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_204
timestamp 1636968456
transform 1 0 19320 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_216
timestamp 1
transform 1 0 20424 0 -1 41888
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_255
timestamp 1636968456
transform 1 0 24012 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_267
timestamp 1636968456
transform 1 0 25116 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1
transform 1 0 26220 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 1
transform 1 0 30820 0 -1 41888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1636968456
transform 1 0 828 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1636968456
transform 1 0 1932 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1
transform 1 0 3036 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1636968456
transform 1 0 3220 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1636968456
transform 1 0 4324 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1636968456
transform 1 0 5428 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1636968456
transform 1 0 6532 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1
transform 1 0 7636 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1
transform 1 0 8188 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1636968456
transform 1 0 8372 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1636968456
transform 1 0 9476 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1636968456
transform 1 0 10580 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1636968456
transform 1 0 11684 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1
transform 1 0 12788 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1
transform 1 0 13340 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_149
timestamp 1
transform 1 0 14260 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_156
timestamp 1
transform 1 0 14904 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_166
timestamp 1
transform 1 0 15824 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_179
timestamp 1
transform 1 0 17020 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_185
timestamp 1
transform 1 0 17572 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_208
timestamp 1
transform 1 0 19688 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_238
timestamp 1
transform 1 0 22448 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_249
timestamp 1
transform 1 0 23460 0 1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_260
timestamp 1636968456
transform 1 0 24472 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_272
timestamp 1
transform 1 0 25576 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_280
timestamp 1
transform 1 0 26312 0 1 41888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_285
timestamp 1636968456
transform 1 0 26772 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_297
timestamp 1
transform 1 0 27876 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 1
transform 1 0 28244 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 1
transform 1 0 28796 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_325
timestamp 1
transform 1 0 30452 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_333
timestamp 1
transform 1 0 31188 0 1 41888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1636968456
transform 1 0 828 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1636968456
transform 1 0 1932 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1636968456
transform 1 0 3036 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1636968456
transform 1 0 4140 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1
transform 1 0 5244 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1
transform 1 0 5612 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1636968456
transform 1 0 5796 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1636968456
transform 1 0 6900 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1636968456
transform 1 0 8004 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_93
timestamp 1
transform 1 0 9108 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_121
timestamp 1
transform 1 0 11684 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_128
timestamp 1
transform 1 0 12328 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_169
timestamp 1
transform 1 0 16100 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_180
timestamp 1
transform 1 0 17112 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_216
timestamp 1
transform 1 0 20424 0 -1 42976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_262
timestamp 1636968456
transform 1 0 24656 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_274
timestamp 1
transform 1 0 25760 0 -1 42976
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1636968456
transform 1 0 26404 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1636968456
transform 1 0 27508 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_305
timestamp 1
transform 1 0 28612 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_313
timestamp 1
transform 1 0 29348 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1636968456
transform 1 0 29716 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 1
transform 1 0 30820 0 -1 42976
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1636968456
transform 1 0 828 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1636968456
transform 1 0 1932 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1
transform 1 0 3036 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1636968456
transform 1 0 3220 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1636968456
transform 1 0 4324 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1636968456
transform 1 0 5428 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1636968456
transform 1 0 6532 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1
transform 1 0 7636 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1
transform 1 0 8188 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_85
timestamp 1
transform 1 0 8372 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_89
timestamp 1
transform 1 0 8740 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_95
timestamp 1
transform 1 0 9292 0 1 42976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_103
timestamp 1636968456
transform 1 0 10028 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_115
timestamp 1
transform 1 0 11132 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_122
timestamp 1
transform 1 0 11776 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_145
timestamp 1
transform 1 0 13892 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_180
timestamp 1
transform 1 0 17112 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 1
transform 1 0 18492 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_200
timestamp 1
transform 1 0 18952 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_218
timestamp 1
transform 1 0 20608 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_222
timestamp 1
transform 1 0 20976 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_229
timestamp 1
transform 1 0 21620 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 1
transform 1 0 28244 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 1
transform 1 0 28796 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1636968456
transform 1 0 28980 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1636968456
transform 1 0 30084 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_333
timestamp 1
transform 1 0 31188 0 1 42976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1636968456
transform 1 0 828 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1636968456
transform 1 0 1932 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1636968456
transform 1 0 3036 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1636968456
transform 1 0 4140 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 1
transform 1 0 5244 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1
transform 1 0 5612 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_57
timestamp 1
transform 1 0 5796 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_63
timestamp 1
transform 1 0 6348 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_72
timestamp 1636968456
transform 1 0 7176 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_173
timestamp 1
transform 1 0 16468 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_195
timestamp 1
transform 1 0 18492 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_222
timestamp 1
transform 1 0 20976 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_241
timestamp 1
transform 1 0 22724 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_250
timestamp 1
transform 1 0 23552 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_254
timestamp 1
transform 1 0 23920 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_271
timestamp 1
transform 1 0 25484 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 1
transform 1 0 26220 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_313
timestamp 1636968456
transform 1 0 29348 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_325
timestamp 1
transform 1 0 30452 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_333
timestamp 1
transform 1 0 31188 0 -1 44064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 1636968456
transform 1 0 828 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 1636968456
transform 1 0 1932 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 1
transform 1 0 3036 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1636968456
transform 1 0 3220 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1636968456
transform 1 0 4324 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_53
timestamp 1
transform 1 0 5428 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_57
timestamp 1636968456
transform 1 0 5796 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_69
timestamp 1
transform 1 0 6900 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_85
timestamp 1
transform 1 0 8372 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_91
timestamp 1
transform 1 0 8924 0 1 44064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1636968456
transform 1 0 9476 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_109
timestamp 1
transform 1 0 10580 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_113
timestamp 1
transform 1 0 10948 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_124
timestamp 1
transform 1 0 11960 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_132
timestamp 1
transform 1 0 12696 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 1
transform 1 0 13340 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_148
timestamp 1
transform 1 0 14168 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_153
timestamp 1
transform 1 0 14628 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_160
timestamp 1
transform 1 0 15272 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_169
timestamp 1
transform 1 0 16100 0 1 44064
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_180
timestamp 1636968456
transform 1 0 17112 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_192
timestamp 1
transform 1 0 18216 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_197
timestamp 1
transform 1 0 18676 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_203
timestamp 1
transform 1 0 19228 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_207
timestamp 1636968456
transform 1 0 19596 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_219
timestamp 1
transform 1 0 20700 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_223
timestamp 1
transform 1 0 21068 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_225
timestamp 1
transform 1 0 21252 0 1 44064
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_232
timestamp 1636968456
transform 1 0 21896 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_244
timestamp 1
transform 1 0 23000 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_256
timestamp 1
transform 1 0 24104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_262
timestamp 1
transform 1 0 24656 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_268
timestamp 1
transform 1 0 25208 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_303
timestamp 1
transform 1 0 28428 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 1
transform 1 0 28796 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_319
timestamp 1636968456
transform 1 0 29900 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_331
timestamp 1
transform 1 0 31004 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 26128 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 14076 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 19412 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 18400 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 17664 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 26220 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 29716 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform 1 0 29624 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 14260 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform 1 0 30636 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 31372 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 28428 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform 1 0 28428 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 24564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 18308 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 10488 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform 1 0 17480 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 18032 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 22448 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform 1 0 23828 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform 1 0 15364 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 16836 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 30544 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 17020 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 20976 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 22908 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 29808 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform 1 0 28336 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 27876 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 30452 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 16836 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 14720 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 12604 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform -1 0 10304 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 13156 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 18952 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 19688 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 19412 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 27140 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 10028 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform -1 0 11684 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 10396 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform -1 0 14260 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 15916 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform 1 0 13616 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 23828 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 16008 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 27600 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 14444 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform -1 0 28980 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 19412 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 16836 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform -1 0 17112 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1
transform 1 0 28980 0 1 44064
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 28428 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 28152 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 26036 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 26312 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 25760 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 25208 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 24656 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform 1 0 23828 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform -1 0 21896 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap18
timestamp 1
transform -1 0 15916 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap19
timestamp 1
transform 1 0 16284 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap20
timestamp 1
transform 1 0 17664 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_81
timestamp 1
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_82
timestamp 1
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_83
timestamp 1
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_84
timestamp 1
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_85
timestamp 1
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_86
timestamp 1
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_87
timestamp 1
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_88
timestamp 1
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_89
timestamp 1
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_90
timestamp 1
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_91
timestamp 1
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_92
timestamp 1
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_93
timestamp 1
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_94
timestamp 1
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_95
timestamp 1
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_96
timestamp 1
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_97
timestamp 1
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_98
timestamp 1
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_99
timestamp 1
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_100
timestamp 1
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_101
timestamp 1
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_102
timestamp 1
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_103
timestamp 1
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_104
timestamp 1
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_105
timestamp 1
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_106
timestamp 1
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_107
timestamp 1
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_108
timestamp 1
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_109
timestamp 1
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_110
timestamp 1
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_111
timestamp 1
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_112
timestamp 1
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_113
timestamp 1
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_114
timestamp 1
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_115
timestamp 1
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_116
timestamp 1
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_117
timestamp 1
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_118
timestamp 1
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_119
timestamp 1
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_120
timestamp 1
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 31648 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_121
timestamp 1
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 31648 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_122
timestamp 1
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 31648 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_123
timestamp 1
transform 1 0 552 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 31648 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_124
timestamp 1
transform 1 0 552 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 31648 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_125
timestamp 1
transform 1 0 552 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 31648 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_126
timestamp 1
transform 1 0 552 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 31648 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_127
timestamp 1
transform 1 0 552 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 31648 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_128
timestamp 1
transform 1 0 552 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 31648 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_129
timestamp 1
transform 1 0 552 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 31648 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_130
timestamp 1
transform 1 0 552 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 31648 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_131
timestamp 1
transform 1 0 552 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 31648 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_132
timestamp 1
transform 1 0 552 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 31648 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_133
timestamp 1
transform 1 0 552 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 31648 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_134
timestamp 1
transform 1 0 552 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 31648 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_135
timestamp 1
transform 1 0 552 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1
transform -1 0 31648 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_136
timestamp 1
transform 1 0 552 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1
transform -1 0 31648 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_137
timestamp 1
transform 1 0 552 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1
transform -1 0 31648 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_138
timestamp 1
transform 1 0 552 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1
transform -1 0 31648 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_139
timestamp 1
transform 1 0 552 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1
transform -1 0 31648 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_140
timestamp 1
transform 1 0 552 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1
transform -1 0 31648 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_141
timestamp 1
transform 1 0 552 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1
transform -1 0 31648 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_142
timestamp 1
transform 1 0 552 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1
transform -1 0 31648 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_143
timestamp 1
transform 1 0 552 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1
transform -1 0 31648 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_144
timestamp 1
transform 1 0 552 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1
transform -1 0 31648 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_145
timestamp 1
transform 1 0 552 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1
transform -1 0 31648 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_146
timestamp 1
transform 1 0 552 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1
transform -1 0 31648 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_147
timestamp 1
transform 1 0 552 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1
transform -1 0 31648 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_148
timestamp 1
transform 1 0 552 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1
transform -1 0 31648 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_149
timestamp 1
transform 1 0 552 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1
transform -1 0 31648 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_150
timestamp 1
transform 1 0 552 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1
transform -1 0 31648 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_151
timestamp 1
transform 1 0 552 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1
transform -1 0 31648 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_152
timestamp 1
transform 1 0 552 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1
transform -1 0 31648 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_153
timestamp 1
transform 1 0 552 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1
transform -1 0 31648 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_154
timestamp 1
transform 1 0 552 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1
transform -1 0 31648 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_155
timestamp 1
transform 1 0 552 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1
transform -1 0 31648 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_156
timestamp 1
transform 1 0 552 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1
transform -1 0 31648 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_157
timestamp 1
transform 1 0 552 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1
transform -1 0 31648 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_158
timestamp 1
transform 1 0 552 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1
transform -1 0 31648 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_159
timestamp 1
transform 1 0 552 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 1
transform -1 0 31648 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_160
timestamp 1
transform 1 0 552 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 1
transform -1 0 31648 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_161
timestamp 1
transform 1 0 552 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 1
transform -1 0 31648 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_162
timestamp 1
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_163
timestamp 1
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_164
timestamp 1
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_165
timestamp 1
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_166
timestamp 1
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_167
timestamp 1
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_168
timestamp 1
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_169
timestamp 1
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_170
timestamp 1
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_171
timestamp 1
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_172
timestamp 1
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_173
timestamp 1
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_174
timestamp 1
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_175
timestamp 1
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_176
timestamp 1
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_177
timestamp 1
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_178
timestamp 1
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_179
timestamp 1
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_180
timestamp 1
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 1
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_182
timestamp 1
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_183
timestamp 1
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_184
timestamp 1
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_185
timestamp 1
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_186
timestamp 1
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_187
timestamp 1
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_188
timestamp 1
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_189
timestamp 1
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_190
timestamp 1
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_191
timestamp 1
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_192
timestamp 1
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_193
timestamp 1
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_194
timestamp 1
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_195
timestamp 1
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_196
timestamp 1
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_197
timestamp 1
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_198
timestamp 1
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_199
timestamp 1
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_200
timestamp 1
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_201
timestamp 1
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_202
timestamp 1
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_203
timestamp 1
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_204
timestamp 1
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_205
timestamp 1
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_206
timestamp 1
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_207
timestamp 1
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_208
timestamp 1
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_209
timestamp 1
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_210
timestamp 1
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_211
timestamp 1
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_212
timestamp 1
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_213
timestamp 1
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_214
timestamp 1
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_215
timestamp 1
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_216
timestamp 1
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_217
timestamp 1
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_218
timestamp 1
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_219
timestamp 1
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_220
timestamp 1
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_221
timestamp 1
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_222
timestamp 1
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_223
timestamp 1
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_224
timestamp 1
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_225
timestamp 1
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_226
timestamp 1
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_227
timestamp 1
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_228
timestamp 1
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_229
timestamp 1
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_230
timestamp 1
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_231
timestamp 1
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_232
timestamp 1
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_233
timestamp 1
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_234
timestamp 1
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_235
timestamp 1
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_236
timestamp 1
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_237
timestamp 1
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_238
timestamp 1
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_239
timestamp 1
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_240
timestamp 1
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_241
timestamp 1
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_242
timestamp 1
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_243
timestamp 1
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_244
timestamp 1
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_245
timestamp 1
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_246
timestamp 1
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_247
timestamp 1
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_248
timestamp 1
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_249
timestamp 1
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_250
timestamp 1
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_251
timestamp 1
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_252
timestamp 1
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_253
timestamp 1
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_254
timestamp 1
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_255
timestamp 1
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_256
timestamp 1
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_257
timestamp 1
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_258
timestamp 1
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_259
timestamp 1
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_260
timestamp 1
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_261
timestamp 1
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_262
timestamp 1
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_263
timestamp 1
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_264
timestamp 1
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_265
timestamp 1
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_266
timestamp 1
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_267
timestamp 1
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_268
timestamp 1
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_269
timestamp 1
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_270
timestamp 1
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_271
timestamp 1
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_272
timestamp 1
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_273
timestamp 1
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_274
timestamp 1
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_275
timestamp 1
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_276
timestamp 1
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_277
timestamp 1
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_278
timestamp 1
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_279
timestamp 1
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_280
timestamp 1
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_281
timestamp 1
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_282
timestamp 1
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_283
timestamp 1
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_284
timestamp 1
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_285
timestamp 1
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_286
timestamp 1
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_287
timestamp 1
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_288
timestamp 1
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_289
timestamp 1
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_290
timestamp 1
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_291
timestamp 1
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_292
timestamp 1
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_293
timestamp 1
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_294
timestamp 1
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_295
timestamp 1
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_296
timestamp 1
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_297
timestamp 1
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_298
timestamp 1
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_299
timestamp 1
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_300
timestamp 1
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_301
timestamp 1
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_302
timestamp 1
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_303
timestamp 1
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_304
timestamp 1
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_305
timestamp 1
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_306
timestamp 1
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_307
timestamp 1
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_308
timestamp 1
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_309
timestamp 1
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_310
timestamp 1
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_311
timestamp 1
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_312
timestamp 1
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_313
timestamp 1
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_314
timestamp 1
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_315
timestamp 1
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_316
timestamp 1
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_317
timestamp 1
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_318
timestamp 1
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_319
timestamp 1
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_320
timestamp 1
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_321
timestamp 1
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_322
timestamp 1
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_323
timestamp 1
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_324
timestamp 1
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_325
timestamp 1
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_326
timestamp 1
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_327
timestamp 1
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_328
timestamp 1
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_329
timestamp 1
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_330
timestamp 1
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_331
timestamp 1
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_332
timestamp 1
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_333
timestamp 1
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_334
timestamp 1
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_335
timestamp 1
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_336
timestamp 1
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_337
timestamp 1
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_338
timestamp 1
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_339
timestamp 1
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_340
timestamp 1
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_341
timestamp 1
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_342
timestamp 1
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_343
timestamp 1
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_344
timestamp 1
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_345
timestamp 1
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_346
timestamp 1
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_347
timestamp 1
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_348
timestamp 1
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_349
timestamp 1
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_350
timestamp 1
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_351
timestamp 1
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_352
timestamp 1
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_353
timestamp 1
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_354
timestamp 1
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_355
timestamp 1
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_356
timestamp 1
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_357
timestamp 1
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_358
timestamp 1
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_359
timestamp 1
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_360
timestamp 1
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_361
timestamp 1
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_362
timestamp 1
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_363
timestamp 1
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_364
timestamp 1
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_365
timestamp 1
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_366
timestamp 1
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_367
timestamp 1
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_368
timestamp 1
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_369
timestamp 1
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_370
timestamp 1
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_371
timestamp 1
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_372
timestamp 1
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_373
timestamp 1
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_374
timestamp 1
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_375
timestamp 1
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_376
timestamp 1
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_377
timestamp 1
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_378
timestamp 1
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_379
timestamp 1
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_380
timestamp 1
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_381
timestamp 1
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_382
timestamp 1
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_383
timestamp 1
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_384
timestamp 1
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_385
timestamp 1
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_386
timestamp 1
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_387
timestamp 1
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_388
timestamp 1
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_389
timestamp 1
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_390
timestamp 1
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_391
timestamp 1
transform 1 0 23736 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_392
timestamp 1
transform 1 0 28888 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_393
timestamp 1
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_394
timestamp 1
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_395
timestamp 1
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_396
timestamp 1
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_397
timestamp 1
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_398
timestamp 1
transform 1 0 3128 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_399
timestamp 1
transform 1 0 8280 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_400
timestamp 1
transform 1 0 13432 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_401
timestamp 1
transform 1 0 18584 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_402
timestamp 1
transform 1 0 23736 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_403
timestamp 1
transform 1 0 28888 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_404
timestamp 1
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_405
timestamp 1
transform 1 0 10856 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_406
timestamp 1
transform 1 0 16008 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_407
timestamp 1
transform 1 0 21160 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_408
timestamp 1
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_409
timestamp 1
transform 1 0 3128 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_410
timestamp 1
transform 1 0 8280 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_411
timestamp 1
transform 1 0 13432 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_412
timestamp 1
transform 1 0 18584 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_413
timestamp 1
transform 1 0 23736 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_414
timestamp 1
transform 1 0 28888 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_415
timestamp 1
transform 1 0 5704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_416
timestamp 1
transform 1 0 10856 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_417
timestamp 1
transform 1 0 16008 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_418
timestamp 1
transform 1 0 21160 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_419
timestamp 1
transform 1 0 26312 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_420
timestamp 1
transform 1 0 3128 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_421
timestamp 1
transform 1 0 8280 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_422
timestamp 1
transform 1 0 13432 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_423
timestamp 1
transform 1 0 18584 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_424
timestamp 1
transform 1 0 23736 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_425
timestamp 1
transform 1 0 28888 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_426
timestamp 1
transform 1 0 5704 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_427
timestamp 1
transform 1 0 10856 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_428
timestamp 1
transform 1 0 16008 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_429
timestamp 1
transform 1 0 21160 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_430
timestamp 1
transform 1 0 26312 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_431
timestamp 1
transform 1 0 3128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_432
timestamp 1
transform 1 0 8280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_433
timestamp 1
transform 1 0 13432 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_434
timestamp 1
transform 1 0 18584 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_435
timestamp 1
transform 1 0 23736 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_436
timestamp 1
transform 1 0 28888 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_437
timestamp 1
transform 1 0 5704 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_438
timestamp 1
transform 1 0 10856 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_439
timestamp 1
transform 1 0 16008 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_440
timestamp 1
transform 1 0 21160 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_441
timestamp 1
transform 1 0 26312 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_442
timestamp 1
transform 1 0 3128 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_443
timestamp 1
transform 1 0 8280 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_444
timestamp 1
transform 1 0 13432 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_445
timestamp 1
transform 1 0 18584 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_446
timestamp 1
transform 1 0 23736 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_447
timestamp 1
transform 1 0 28888 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_448
timestamp 1
transform 1 0 5704 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_449
timestamp 1
transform 1 0 10856 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_450
timestamp 1
transform 1 0 16008 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_451
timestamp 1
transform 1 0 21160 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_452
timestamp 1
transform 1 0 26312 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_453
timestamp 1
transform 1 0 3128 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_454
timestamp 1
transform 1 0 8280 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_455
timestamp 1
transform 1 0 13432 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_456
timestamp 1
transform 1 0 18584 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_457
timestamp 1
transform 1 0 23736 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_458
timestamp 1
transform 1 0 28888 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_459
timestamp 1
transform 1 0 5704 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_460
timestamp 1
transform 1 0 10856 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_461
timestamp 1
transform 1 0 16008 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_462
timestamp 1
transform 1 0 21160 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_463
timestamp 1
transform 1 0 26312 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_464
timestamp 1
transform 1 0 3128 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_465
timestamp 1
transform 1 0 8280 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_466
timestamp 1
transform 1 0 13432 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_467
timestamp 1
transform 1 0 18584 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_468
timestamp 1
transform 1 0 23736 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_469
timestamp 1
transform 1 0 28888 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_470
timestamp 1
transform 1 0 5704 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_471
timestamp 1
transform 1 0 10856 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_472
timestamp 1
transform 1 0 16008 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_473
timestamp 1
transform 1 0 21160 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_474
timestamp 1
transform 1 0 26312 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_475
timestamp 1
transform 1 0 3128 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_476
timestamp 1
transform 1 0 8280 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_477
timestamp 1
transform 1 0 13432 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_478
timestamp 1
transform 1 0 18584 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_479
timestamp 1
transform 1 0 23736 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_480
timestamp 1
transform 1 0 28888 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_481
timestamp 1
transform 1 0 5704 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_482
timestamp 1
transform 1 0 10856 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_483
timestamp 1
transform 1 0 16008 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_484
timestamp 1
transform 1 0 21160 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_485
timestamp 1
transform 1 0 26312 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_486
timestamp 1
transform 1 0 3128 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_487
timestamp 1
transform 1 0 8280 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_488
timestamp 1
transform 1 0 13432 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_489
timestamp 1
transform 1 0 18584 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_490
timestamp 1
transform 1 0 23736 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_491
timestamp 1
transform 1 0 28888 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_492
timestamp 1
transform 1 0 5704 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_493
timestamp 1
transform 1 0 10856 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_494
timestamp 1
transform 1 0 16008 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_495
timestamp 1
transform 1 0 21160 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_496
timestamp 1
transform 1 0 26312 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_497
timestamp 1
transform 1 0 3128 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_498
timestamp 1
transform 1 0 8280 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_499
timestamp 1
transform 1 0 13432 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_500
timestamp 1
transform 1 0 18584 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_501
timestamp 1
transform 1 0 23736 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_502
timestamp 1
transform 1 0 28888 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_503
timestamp 1
transform 1 0 5704 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_504
timestamp 1
transform 1 0 10856 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_505
timestamp 1
transform 1 0 16008 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_506
timestamp 1
transform 1 0 21160 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_507
timestamp 1
transform 1 0 26312 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_508
timestamp 1
transform 1 0 3128 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_509
timestamp 1
transform 1 0 8280 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_510
timestamp 1
transform 1 0 13432 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_511
timestamp 1
transform 1 0 18584 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_512
timestamp 1
transform 1 0 23736 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_513
timestamp 1
transform 1 0 28888 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_514
timestamp 1
transform 1 0 5704 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_515
timestamp 1
transform 1 0 10856 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_516
timestamp 1
transform 1 0 16008 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_517
timestamp 1
transform 1 0 21160 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_518
timestamp 1
transform 1 0 26312 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_519
timestamp 1
transform 1 0 3128 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_520
timestamp 1
transform 1 0 8280 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_521
timestamp 1
transform 1 0 13432 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_522
timestamp 1
transform 1 0 18584 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_523
timestamp 1
transform 1 0 23736 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_524
timestamp 1
transform 1 0 28888 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_525
timestamp 1
transform 1 0 5704 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_526
timestamp 1
transform 1 0 10856 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_527
timestamp 1
transform 1 0 16008 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_528
timestamp 1
transform 1 0 21160 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_529
timestamp 1
transform 1 0 26312 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_530
timestamp 1
transform 1 0 3128 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_531
timestamp 1
transform 1 0 8280 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_532
timestamp 1
transform 1 0 13432 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_533
timestamp 1
transform 1 0 18584 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_534
timestamp 1
transform 1 0 23736 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_535
timestamp 1
transform 1 0 28888 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_536
timestamp 1
transform 1 0 5704 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_537
timestamp 1
transform 1 0 10856 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_538
timestamp 1
transform 1 0 16008 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_539
timestamp 1
transform 1 0 21160 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_540
timestamp 1
transform 1 0 26312 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_541
timestamp 1
transform 1 0 3128 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_542
timestamp 1
transform 1 0 8280 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_543
timestamp 1
transform 1 0 13432 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_544
timestamp 1
transform 1 0 18584 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_545
timestamp 1
transform 1 0 23736 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_546
timestamp 1
transform 1 0 28888 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_547
timestamp 1
transform 1 0 5704 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_548
timestamp 1
transform 1 0 10856 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_549
timestamp 1
transform 1 0 16008 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_550
timestamp 1
transform 1 0 21160 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_551
timestamp 1
transform 1 0 26312 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_552
timestamp 1
transform 1 0 3128 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_553
timestamp 1
transform 1 0 8280 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_554
timestamp 1
transform 1 0 13432 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_555
timestamp 1
transform 1 0 18584 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_556
timestamp 1
transform 1 0 23736 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_557
timestamp 1
transform 1 0 28888 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_558
timestamp 1
transform 1 0 5704 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_559
timestamp 1
transform 1 0 10856 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_560
timestamp 1
transform 1 0 16008 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_561
timestamp 1
transform 1 0 21160 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_562
timestamp 1
transform 1 0 26312 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_563
timestamp 1
transform 1 0 3128 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_564
timestamp 1
transform 1 0 8280 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_565
timestamp 1
transform 1 0 13432 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_566
timestamp 1
transform 1 0 18584 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_567
timestamp 1
transform 1 0 23736 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_568
timestamp 1
transform 1 0 28888 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_569
timestamp 1
transform 1 0 5704 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_570
timestamp 1
transform 1 0 10856 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_571
timestamp 1
transform 1 0 16008 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_572
timestamp 1
transform 1 0 21160 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_573
timestamp 1
transform 1 0 26312 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_574
timestamp 1
transform 1 0 3128 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_575
timestamp 1
transform 1 0 8280 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_576
timestamp 1
transform 1 0 13432 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_577
timestamp 1
transform 1 0 18584 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_578
timestamp 1
transform 1 0 23736 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_579
timestamp 1
transform 1 0 28888 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_580
timestamp 1
transform 1 0 5704 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_581
timestamp 1
transform 1 0 10856 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_582
timestamp 1
transform 1 0 16008 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_583
timestamp 1
transform 1 0 21160 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_584
timestamp 1
transform 1 0 26312 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_585
timestamp 1
transform 1 0 3128 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_586
timestamp 1
transform 1 0 8280 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_587
timestamp 1
transform 1 0 13432 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_588
timestamp 1
transform 1 0 18584 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_589
timestamp 1
transform 1 0 23736 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_590
timestamp 1
transform 1 0 28888 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_591
timestamp 1
transform 1 0 5704 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_592
timestamp 1
transform 1 0 10856 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_593
timestamp 1
transform 1 0 16008 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_594
timestamp 1
transform 1 0 21160 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_595
timestamp 1
transform 1 0 26312 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_596
timestamp 1
transform 1 0 3128 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_597
timestamp 1
transform 1 0 8280 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_598
timestamp 1
transform 1 0 13432 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_599
timestamp 1
transform 1 0 18584 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_600
timestamp 1
transform 1 0 23736 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_601
timestamp 1
transform 1 0 28888 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_602
timestamp 1
transform 1 0 5704 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_603
timestamp 1
transform 1 0 10856 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_604
timestamp 1
transform 1 0 16008 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_605
timestamp 1
transform 1 0 21160 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_606
timestamp 1
transform 1 0 26312 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_607
timestamp 1
transform 1 0 3128 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_608
timestamp 1
transform 1 0 5704 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_609
timestamp 1
transform 1 0 8280 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_610
timestamp 1
transform 1 0 10856 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_611
timestamp 1
transform 1 0 13432 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_612
timestamp 1
transform 1 0 16008 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_613
timestamp 1
transform 1 0 18584 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_614
timestamp 1
transform 1 0 21160 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_615
timestamp 1
transform 1 0 23736 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_616
timestamp 1
transform 1 0 26312 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_617
timestamp 1
transform 1 0 28888 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_63
timestamp 1
transform 1 0 7728 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_64
timestamp 1
transform 1 0 7452 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_65
timestamp 1
transform -1 0 7452 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_66
timestamp 1
transform -1 0 13064 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_67
timestamp 1
transform -1 0 13340 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_68
timestamp 1
transform -1 0 11960 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire17
timestamp 1
transform -1 0 26220 0 -1 33184
box -38 -48 314 592
<< labels >>
flabel metal4 s 4316 496 4636 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12090 496 12410 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19864 496 20184 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27638 496 27958 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11430 496 11750 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19204 496 19524 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26978 496 27298 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
