VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 71.750 BY 20.300 ;
  OBS
      LAYER met1 ;
        RECT 0.000 19.950 8.050 20.300 ;
      LAYER met1 ;
        RECT 8.050 19.950 11.550 20.300 ;
      LAYER met1 ;
        RECT 11.550 19.950 22.050 20.300 ;
      LAYER met1 ;
        RECT 22.050 19.950 24.500 20.300 ;
      LAYER met1 ;
        RECT 24.500 19.950 31.500 20.300 ;
      LAYER met1 ;
        RECT 31.500 19.950 33.950 20.300 ;
      LAYER met1 ;
        RECT 33.950 19.950 52.500 20.300 ;
      LAYER met1 ;
        RECT 52.500 19.950 54.950 20.300 ;
      LAYER met1 ;
        RECT 54.950 19.950 67.200 20.300 ;
      LAYER met1 ;
        RECT 67.200 19.950 69.650 20.300 ;
      LAYER met1 ;
        RECT 69.650 19.950 71.750 20.300 ;
        RECT 0.000 19.600 6.650 19.950 ;
      LAYER met1 ;
        RECT 6.650 19.600 12.950 19.950 ;
      LAYER met1 ;
        RECT 12.950 19.600 21.700 19.950 ;
      LAYER met1 ;
        RECT 21.700 19.600 24.500 19.950 ;
      LAYER met1 ;
        RECT 24.500 19.600 30.450 19.950 ;
      LAYER met1 ;
        RECT 30.450 19.600 34.650 19.950 ;
      LAYER met1 ;
        RECT 34.650 19.600 40.950 19.950 ;
      LAYER met1 ;
        RECT 40.950 19.600 43.750 19.950 ;
      LAYER met1 ;
        RECT 43.750 19.600 46.900 19.950 ;
      LAYER met1 ;
        RECT 46.900 19.600 49.700 19.950 ;
      LAYER met1 ;
        RECT 49.700 19.600 51.800 19.950 ;
      LAYER met1 ;
        RECT 51.800 19.600 55.650 19.950 ;
      LAYER met1 ;
        RECT 55.650 19.600 57.050 19.950 ;
      LAYER met1 ;
        RECT 57.050 19.600 60.200 19.950 ;
      LAYER met1 ;
        RECT 60.200 19.600 66.500 19.950 ;
      LAYER met1 ;
        RECT 66.500 19.600 70.350 19.950 ;
      LAYER met1 ;
        RECT 70.350 19.600 71.750 19.950 ;
        RECT 0.000 19.250 5.600 19.600 ;
      LAYER met1 ;
        RECT 5.600 19.250 13.650 19.600 ;
      LAYER met1 ;
        RECT 13.650 19.250 21.000 19.600 ;
      LAYER met1 ;
        RECT 21.000 19.250 24.500 19.600 ;
      LAYER met1 ;
        RECT 24.500 19.250 30.100 19.600 ;
      LAYER met1 ;
        RECT 30.100 19.250 32.200 19.600 ;
      LAYER met1 ;
        RECT 32.200 19.250 33.250 19.600 ;
      LAYER met1 ;
        RECT 33.250 19.250 35.350 19.600 ;
      LAYER met1 ;
        RECT 35.350 19.250 41.650 19.600 ;
      LAYER met1 ;
        RECT 41.650 19.250 43.050 19.600 ;
      LAYER met1 ;
        RECT 0.000 18.900 4.900 19.250 ;
      LAYER met1 ;
        RECT 4.900 18.900 14.350 19.250 ;
      LAYER met1 ;
        RECT 14.350 18.900 20.300 19.250 ;
      LAYER met1 ;
        RECT 20.300 18.900 24.500 19.250 ;
      LAYER met1 ;
        RECT 24.500 18.900 29.750 19.250 ;
      LAYER met1 ;
        RECT 29.750 18.900 31.850 19.250 ;
      LAYER met1 ;
        RECT 31.850 18.900 33.600 19.250 ;
      LAYER met1 ;
        RECT 33.600 18.900 35.700 19.250 ;
      LAYER met1 ;
        RECT 35.700 18.900 42.000 19.250 ;
      LAYER met1 ;
        RECT 42.000 18.900 43.050 19.250 ;
      LAYER met1 ;
        RECT 43.050 18.900 47.600 19.600 ;
      LAYER met1 ;
        RECT 47.600 18.900 48.650 19.600 ;
      LAYER met1 ;
        RECT 48.650 19.250 51.450 19.600 ;
      LAYER met1 ;
        RECT 51.450 19.250 52.500 19.600 ;
      LAYER met1 ;
        RECT 52.500 19.250 53.900 19.600 ;
      LAYER met1 ;
        RECT 53.900 19.250 55.650 19.600 ;
      LAYER met1 ;
        RECT 55.650 19.250 57.750 19.600 ;
      LAYER met1 ;
        RECT 57.750 19.250 59.500 19.600 ;
      LAYER met1 ;
        RECT 59.500 19.250 65.800 19.600 ;
      LAYER met1 ;
        RECT 65.800 19.250 67.200 19.600 ;
      LAYER met1 ;
        RECT 67.200 19.250 68.250 19.600 ;
      LAYER met1 ;
        RECT 68.250 19.250 70.700 19.600 ;
      LAYER met1 ;
        RECT 70.700 19.250 71.750 19.600 ;
        RECT 48.650 18.900 51.100 19.250 ;
      LAYER met1 ;
        RECT 51.100 18.900 52.150 19.250 ;
      LAYER met1 ;
        RECT 52.150 18.900 54.600 19.250 ;
      LAYER met1 ;
        RECT 54.600 18.900 55.650 19.250 ;
      LAYER met1 ;
        RECT 55.650 18.900 58.100 19.250 ;
        RECT 0.000 18.550 4.550 18.900 ;
      LAYER met1 ;
        RECT 4.550 18.550 8.750 18.900 ;
      LAYER met1 ;
        RECT 8.750 18.550 10.850 18.900 ;
      LAYER met1 ;
        RECT 10.850 18.550 15.050 18.900 ;
      LAYER met1 ;
        RECT 15.050 18.550 19.950 18.900 ;
      LAYER met1 ;
        RECT 19.950 18.550 21.700 18.900 ;
      LAYER met1 ;
        RECT 21.700 18.550 22.050 18.900 ;
        RECT 0.000 18.200 3.850 18.550 ;
      LAYER met1 ;
        RECT 3.850 18.200 7.000 18.550 ;
      LAYER met1 ;
        RECT 7.000 18.200 12.250 18.550 ;
      LAYER met1 ;
        RECT 12.250 18.200 15.400 18.550 ;
      LAYER met1 ;
        RECT 15.400 18.200 19.950 18.550 ;
      LAYER met1 ;
        RECT 19.950 18.200 21.000 18.550 ;
      LAYER met1 ;
        RECT 21.000 18.200 22.050 18.550 ;
        RECT 0.000 17.850 3.500 18.200 ;
      LAYER met1 ;
        RECT 3.500 17.850 6.300 18.200 ;
      LAYER met1 ;
        RECT 6.300 17.850 13.300 18.200 ;
      LAYER met1 ;
        RECT 13.300 17.850 16.100 18.200 ;
      LAYER met1 ;
        RECT 16.100 17.850 19.950 18.200 ;
      LAYER met1 ;
        RECT 19.950 17.850 20.300 18.200 ;
      LAYER met1 ;
        RECT 20.300 17.850 22.050 18.200 ;
        RECT 0.000 17.500 3.150 17.850 ;
      LAYER met1 ;
        RECT 3.150 17.500 5.600 17.850 ;
      LAYER met1 ;
        RECT 5.600 17.500 14.000 17.850 ;
      LAYER met1 ;
        RECT 14.000 17.500 16.450 17.850 ;
      LAYER met1 ;
        RECT 16.450 17.500 22.050 17.850 ;
        RECT 0.000 17.150 2.800 17.500 ;
      LAYER met1 ;
        RECT 2.800 17.150 4.900 17.500 ;
      LAYER met1 ;
        RECT 4.900 17.150 14.350 17.500 ;
      LAYER met1 ;
        RECT 14.350 17.150 16.800 17.500 ;
      LAYER met1 ;
        RECT 16.800 17.150 22.050 17.500 ;
        RECT 0.000 16.800 2.450 17.150 ;
      LAYER met1 ;
        RECT 2.450 16.800 4.550 17.150 ;
      LAYER met1 ;
        RECT 4.550 16.800 15.050 17.150 ;
      LAYER met1 ;
        RECT 15.050 16.800 17.150 17.150 ;
      LAYER met1 ;
        RECT 17.150 16.800 22.050 17.150 ;
        RECT 0.000 16.450 2.100 16.800 ;
      LAYER met1 ;
        RECT 2.100 16.450 4.200 16.800 ;
      LAYER met1 ;
        RECT 4.200 16.450 15.400 16.800 ;
      LAYER met1 ;
        RECT 15.400 16.450 17.500 16.800 ;
      LAYER met1 ;
        RECT 0.000 15.750 1.750 16.450 ;
      LAYER met1 ;
        RECT 1.750 16.100 3.850 16.450 ;
      LAYER met1 ;
        RECT 3.850 16.100 15.750 16.450 ;
      LAYER met1 ;
        RECT 15.750 16.100 17.500 16.450 ;
      LAYER met1 ;
        RECT 17.500 16.100 22.050 16.800 ;
      LAYER met1 ;
        RECT 1.750 15.750 11.550 16.100 ;
      LAYER met1 ;
        RECT 0.000 15.050 1.400 15.750 ;
      LAYER met1 ;
        RECT 1.400 15.050 11.550 15.750 ;
      LAYER met1 ;
        RECT 11.550 15.400 16.100 16.100 ;
      LAYER met1 ;
        RECT 16.100 15.750 17.850 16.100 ;
      LAYER met1 ;
        RECT 17.850 15.750 22.050 16.100 ;
      LAYER met1 ;
        RECT 16.100 15.400 18.200 15.750 ;
      LAYER met1 ;
        RECT 11.550 15.050 16.450 15.400 ;
      LAYER met1 ;
        RECT 16.450 15.050 18.200 15.400 ;
      LAYER met1 ;
        RECT 18.200 15.050 22.050 15.750 ;
        RECT 0.000 14.350 1.050 15.050 ;
      LAYER met1 ;
        RECT 1.050 14.350 11.550 15.050 ;
      LAYER met1 ;
        RECT 11.550 14.350 16.800 15.050 ;
      LAYER met1 ;
        RECT 16.800 14.350 18.550 15.050 ;
      LAYER met1 ;
        RECT 18.550 14.350 22.050 15.050 ;
        RECT 0.000 13.650 0.700 14.350 ;
      LAYER met1 ;
        RECT 0.700 13.650 11.550 14.350 ;
      LAYER met1 ;
        RECT 11.550 13.650 17.150 14.350 ;
      LAYER met1 ;
        RECT 17.150 13.650 18.900 14.350 ;
      LAYER met1 ;
        RECT 0.000 13.300 5.600 13.650 ;
      LAYER met1 ;
        RECT 5.600 13.300 8.750 13.650 ;
      LAYER met1 ;
        RECT 0.000 12.600 5.950 13.300 ;
        RECT 0.000 12.250 0.350 12.600 ;
      LAYER met1 ;
        RECT 0.350 12.250 1.750 12.600 ;
        RECT 0.000 11.550 1.750 12.250 ;
      LAYER met1 ;
        RECT 1.750 11.550 5.950 12.600 ;
      LAYER met1 ;
        RECT 0.000 9.450 1.400 11.550 ;
      LAYER met1 ;
        RECT 1.400 9.450 5.950 11.550 ;
      LAYER met1 ;
        RECT 5.950 11.200 8.750 13.300 ;
      LAYER met1 ;
        RECT 8.750 12.950 17.500 13.650 ;
      LAYER met1 ;
        RECT 17.500 13.300 18.900 13.650 ;
      LAYER met1 ;
        RECT 18.900 13.300 22.050 14.350 ;
      LAYER met1 ;
        RECT 17.500 12.950 19.250 13.300 ;
      LAYER met1 ;
        RECT 8.750 11.200 17.850 12.950 ;
      LAYER met1 ;
        RECT 17.850 11.550 19.250 12.950 ;
      LAYER met1 ;
        RECT 19.250 11.550 22.050 13.300 ;
      LAYER met1 ;
        RECT 0.000 8.750 1.750 9.450 ;
      LAYER met1 ;
        RECT 0.000 7.350 0.350 8.750 ;
      LAYER met1 ;
        RECT 0.350 7.700 1.750 8.750 ;
      LAYER met1 ;
        RECT 1.750 7.700 5.950 9.450 ;
      LAYER met1 ;
        RECT 5.950 8.750 16.100 11.200 ;
      LAYER met1 ;
        RECT 16.100 8.750 17.850 11.200 ;
      LAYER met1 ;
        RECT 17.850 9.450 19.600 11.550 ;
      LAYER met1 ;
        RECT 19.600 10.850 22.050 11.550 ;
      LAYER met1 ;
        RECT 22.050 10.850 24.500 18.900 ;
      LAYER met1 ;
        RECT 24.500 18.200 29.400 18.900 ;
      LAYER met1 ;
        RECT 29.400 18.200 31.500 18.900 ;
      LAYER met1 ;
        RECT 24.500 17.500 29.050 18.200 ;
      LAYER met1 ;
        RECT 29.050 17.500 31.500 18.200 ;
      LAYER met1 ;
        RECT 24.500 15.400 28.700 17.500 ;
      LAYER met1 ;
        RECT 28.700 17.150 31.500 17.500 ;
      LAYER met1 ;
        RECT 31.500 17.150 33.950 18.900 ;
      LAYER met1 ;
        RECT 33.950 18.200 36.050 18.900 ;
      LAYER met1 ;
        RECT 36.050 18.200 42.000 18.900 ;
      LAYER met1 ;
        RECT 42.000 18.200 43.400 18.900 ;
      LAYER met1 ;
        RECT 43.400 18.550 47.600 18.900 ;
      LAYER met1 ;
        RECT 47.600 18.550 48.300 18.900 ;
      LAYER met1 ;
        RECT 43.400 18.200 47.250 18.550 ;
      LAYER met1 ;
        RECT 33.950 17.150 36.400 18.200 ;
      LAYER met1 ;
        RECT 36.400 17.150 42.350 18.200 ;
      LAYER met1 ;
        RECT 42.350 17.150 43.750 18.200 ;
      LAYER met1 ;
        RECT 43.750 17.500 47.250 18.200 ;
      LAYER met1 ;
        RECT 47.250 17.850 48.300 18.550 ;
      LAYER met1 ;
        RECT 48.300 17.850 50.750 18.900 ;
      LAYER met1 ;
        RECT 50.750 17.850 51.800 18.900 ;
      LAYER met1 ;
        RECT 51.800 18.550 54.950 18.900 ;
      LAYER met1 ;
        RECT 54.950 18.550 55.300 18.900 ;
      LAYER met1 ;
        RECT 55.300 18.550 58.100 18.900 ;
        RECT 51.800 17.850 58.100 18.550 ;
      LAYER met1 ;
        RECT 47.250 17.500 47.950 17.850 ;
      LAYER met1 ;
        RECT 43.750 17.150 46.900 17.500 ;
      LAYER met1 ;
        RECT 46.900 17.150 47.950 17.500 ;
      LAYER met1 ;
        RECT 47.950 17.150 50.750 17.850 ;
      LAYER met1 ;
        RECT 50.750 17.500 52.150 17.850 ;
      LAYER met1 ;
        RECT 52.150 17.500 58.100 17.850 ;
      LAYER met1 ;
        RECT 50.750 17.150 52.500 17.500 ;
      LAYER met1 ;
        RECT 52.500 17.150 58.100 17.500 ;
      LAYER met1 ;
        RECT 28.700 15.400 31.150 17.150 ;
      LAYER met1 ;
        RECT 24.500 14.700 28.350 15.400 ;
      LAYER met1 ;
        RECT 28.350 14.700 31.150 15.400 ;
      LAYER met1 ;
        RECT 24.500 12.600 28.700 14.700 ;
      LAYER met1 ;
        RECT 28.700 12.950 31.150 14.700 ;
      LAYER met1 ;
        RECT 31.150 12.950 33.950 17.150 ;
      LAYER met1 ;
        RECT 28.700 12.600 31.500 12.950 ;
      LAYER met1 ;
        RECT 24.500 11.550 29.050 12.600 ;
      LAYER met1 ;
        RECT 29.050 11.550 31.500 12.600 ;
      LAYER met1 ;
        RECT 24.500 11.200 29.400 11.550 ;
      LAYER met1 ;
        RECT 29.400 11.200 31.500 11.550 ;
      LAYER met1 ;
        RECT 31.500 11.200 33.950 12.950 ;
      LAYER met1 ;
        RECT 33.950 12.600 36.750 17.150 ;
      LAYER met1 ;
        RECT 36.750 16.450 42.700 17.150 ;
      LAYER met1 ;
        RECT 42.700 16.450 44.100 17.150 ;
      LAYER met1 ;
        RECT 44.100 16.450 46.900 17.150 ;
      LAYER met1 ;
        RECT 46.900 16.450 47.600 17.150 ;
      LAYER met1 ;
        RECT 47.600 16.800 51.100 17.150 ;
      LAYER met1 ;
        RECT 51.100 16.800 53.200 17.150 ;
      LAYER met1 ;
        RECT 53.200 16.800 58.100 17.150 ;
        RECT 47.600 16.450 51.450 16.800 ;
      LAYER met1 ;
        RECT 51.450 16.450 53.900 16.800 ;
      LAYER met1 ;
        RECT 53.900 16.450 58.100 16.800 ;
        RECT 36.750 15.400 43.050 16.450 ;
      LAYER met1 ;
        RECT 43.050 16.100 44.100 16.450 ;
      LAYER met1 ;
        RECT 44.100 16.100 46.550 16.450 ;
      LAYER met1 ;
        RECT 46.550 16.100 47.600 16.450 ;
      LAYER met1 ;
        RECT 47.600 16.100 51.800 16.450 ;
      LAYER met1 ;
        RECT 51.800 16.100 54.600 16.450 ;
      LAYER met1 ;
        RECT 54.600 16.100 58.100 16.450 ;
      LAYER met1 ;
        RECT 43.050 15.400 44.450 16.100 ;
      LAYER met1 ;
        RECT 44.450 15.400 46.550 16.100 ;
      LAYER met1 ;
        RECT 46.550 15.400 47.250 16.100 ;
      LAYER met1 ;
        RECT 47.250 15.750 52.500 16.100 ;
      LAYER met1 ;
        RECT 52.500 15.750 54.950 16.100 ;
      LAYER met1 ;
        RECT 54.950 15.750 58.100 16.100 ;
        RECT 47.250 15.400 53.200 15.750 ;
      LAYER met1 ;
        RECT 53.200 15.400 55.650 15.750 ;
      LAYER met1 ;
        RECT 36.750 14.350 43.400 15.400 ;
      LAYER met1 ;
        RECT 43.400 14.350 44.800 15.400 ;
      LAYER met1 ;
        RECT 44.800 14.700 46.200 15.400 ;
      LAYER met1 ;
        RECT 46.200 15.050 47.250 15.400 ;
      LAYER met1 ;
        RECT 47.250 15.050 53.900 15.400 ;
      LAYER met1 ;
        RECT 53.900 15.050 55.650 15.400 ;
      LAYER met1 ;
        RECT 55.650 15.050 58.100 15.750 ;
      LAYER met1 ;
        RECT 46.200 14.700 46.900 15.050 ;
      LAYER met1 ;
        RECT 46.900 14.700 54.250 15.050 ;
      LAYER met1 ;
        RECT 54.250 14.700 56.000 15.050 ;
      LAYER met1 ;
        RECT 44.800 14.350 45.850 14.700 ;
        RECT 36.750 13.650 43.750 14.350 ;
      LAYER met1 ;
        RECT 43.750 13.650 45.150 14.350 ;
      LAYER met1 ;
        RECT 45.150 13.650 45.850 14.350 ;
      LAYER met1 ;
        RECT 45.850 14.000 46.900 14.700 ;
      LAYER met1 ;
        RECT 46.900 14.350 54.600 14.700 ;
      LAYER met1 ;
        RECT 54.600 14.350 56.000 14.700 ;
      LAYER met1 ;
        RECT 46.900 14.000 54.950 14.350 ;
      LAYER met1 ;
        RECT 45.850 13.650 46.550 14.000 ;
      LAYER met1 ;
        RECT 46.550 13.650 54.950 14.000 ;
        RECT 36.750 12.600 44.100 13.650 ;
      LAYER met1 ;
        RECT 44.100 13.300 45.150 13.650 ;
      LAYER met1 ;
        RECT 45.150 13.300 45.500 13.650 ;
      LAYER met1 ;
        RECT 45.500 13.300 46.550 13.650 ;
        RECT 44.100 12.950 46.550 13.300 ;
      LAYER met1 ;
        RECT 46.550 12.950 50.750 13.650 ;
      LAYER met1 ;
        RECT 50.750 13.300 51.100 13.650 ;
      LAYER met1 ;
        RECT 51.100 13.300 54.950 13.650 ;
      LAYER met1 ;
        RECT 50.750 12.950 51.450 13.300 ;
      LAYER met1 ;
        RECT 51.450 12.950 54.950 13.300 ;
      LAYER met1 ;
        RECT 54.950 12.950 56.000 14.350 ;
        RECT 44.100 12.600 46.200 12.950 ;
        RECT 33.950 11.900 36.400 12.600 ;
      LAYER met1 ;
        RECT 36.400 11.900 44.450 12.600 ;
      LAYER met1 ;
        RECT 44.450 11.900 46.200 12.600 ;
      LAYER met1 ;
        RECT 46.200 11.900 50.750 12.950 ;
      LAYER met1 ;
        RECT 50.750 12.600 51.800 12.950 ;
      LAYER met1 ;
        RECT 51.800 12.600 54.600 12.950 ;
      LAYER met1 ;
        RECT 54.600 12.600 56.000 12.950 ;
      LAYER met1 ;
        RECT 56.000 12.600 58.100 15.050 ;
      LAYER met1 ;
        RECT 50.750 12.250 52.150 12.600 ;
      LAYER met1 ;
        RECT 52.150 12.250 54.250 12.600 ;
      LAYER met1 ;
        RECT 54.250 12.250 55.650 12.600 ;
      LAYER met1 ;
        RECT 55.650 12.250 58.100 12.600 ;
      LAYER met1 ;
        RECT 58.100 12.250 59.500 19.250 ;
      LAYER met1 ;
        RECT 59.500 18.900 65.450 19.250 ;
      LAYER met1 ;
        RECT 65.450 18.900 66.500 19.250 ;
      LAYER met1 ;
        RECT 66.500 18.900 68.950 19.250 ;
      LAYER met1 ;
        RECT 68.950 18.900 70.350 19.250 ;
      LAYER met1 ;
        RECT 70.350 18.900 71.750 19.250 ;
        RECT 59.500 18.550 65.100 18.900 ;
      LAYER met1 ;
        RECT 65.100 18.550 66.150 18.900 ;
      LAYER met1 ;
        RECT 66.150 18.550 69.650 18.900 ;
      LAYER met1 ;
        RECT 69.650 18.550 70.000 18.900 ;
      LAYER met1 ;
        RECT 70.000 18.550 71.750 18.900 ;
        RECT 59.500 17.850 64.750 18.550 ;
      LAYER met1 ;
        RECT 64.750 18.200 66.150 18.550 ;
      LAYER met1 ;
        RECT 66.150 18.200 71.750 18.550 ;
      LAYER met1 ;
        RECT 64.750 17.850 65.800 18.200 ;
      LAYER met1 ;
        RECT 59.500 16.800 64.400 17.850 ;
      LAYER met1 ;
        RECT 64.400 17.500 65.800 17.850 ;
      LAYER met1 ;
        RECT 65.800 17.500 71.750 18.200 ;
      LAYER met1 ;
        RECT 64.400 16.800 65.450 17.500 ;
      LAYER met1 ;
        RECT 59.500 14.000 64.050 16.800 ;
      LAYER met1 ;
        RECT 64.050 14.000 65.450 16.800 ;
      LAYER met1 ;
        RECT 65.450 14.000 71.750 17.500 ;
        RECT 59.500 13.300 64.400 14.000 ;
      LAYER met1 ;
        RECT 64.400 13.300 65.800 14.000 ;
      LAYER met1 ;
        RECT 65.800 13.300 71.750 14.000 ;
        RECT 59.500 12.950 63.000 13.300 ;
      LAYER met1 ;
        RECT 63.000 12.950 63.350 13.300 ;
      LAYER met1 ;
        RECT 59.500 12.250 62.650 12.950 ;
      LAYER met1 ;
        RECT 62.650 12.250 63.350 12.950 ;
      LAYER met1 ;
        RECT 63.350 12.600 64.750 13.300 ;
      LAYER met1 ;
        RECT 64.750 12.950 66.150 13.300 ;
      LAYER met1 ;
        RECT 66.150 12.950 71.750 13.300 ;
      LAYER met1 ;
        RECT 64.750 12.600 66.500 12.950 ;
      LAYER met1 ;
        RECT 66.500 12.600 70.000 12.950 ;
      LAYER met1 ;
        RECT 70.000 12.600 70.700 12.950 ;
      LAYER met1 ;
        RECT 70.700 12.600 71.750 12.950 ;
        RECT 63.350 12.250 65.100 12.600 ;
      LAYER met1 ;
        RECT 65.100 12.250 66.850 12.600 ;
      LAYER met1 ;
        RECT 66.850 12.250 69.300 12.600 ;
      LAYER met1 ;
        RECT 69.300 12.250 70.350 12.600 ;
      LAYER met1 ;
        RECT 70.350 12.250 71.750 12.600 ;
      LAYER met1 ;
        RECT 50.750 11.900 53.200 12.250 ;
      LAYER met1 ;
        RECT 53.200 11.900 53.550 12.250 ;
      LAYER met1 ;
        RECT 53.550 11.900 55.300 12.250 ;
      LAYER met1 ;
        RECT 55.300 11.900 58.100 12.250 ;
      LAYER met1 ;
        RECT 58.100 11.900 60.550 12.250 ;
      LAYER met1 ;
        RECT 60.550 11.900 61.600 12.250 ;
      LAYER met1 ;
        RECT 61.600 11.900 63.350 12.250 ;
      LAYER met1 ;
        RECT 63.350 11.900 65.450 12.250 ;
      LAYER met1 ;
        RECT 65.450 11.900 70.000 12.250 ;
      LAYER met1 ;
        RECT 70.000 11.900 71.750 12.250 ;
      LAYER met1 ;
        RECT 33.950 11.200 36.050 11.900 ;
      LAYER met1 ;
        RECT 36.050 11.550 44.450 11.900 ;
      LAYER met1 ;
        RECT 44.450 11.550 45.850 11.900 ;
      LAYER met1 ;
        RECT 45.850 11.550 51.100 11.900 ;
      LAYER met1 ;
        RECT 51.100 11.550 54.950 11.900 ;
      LAYER met1 ;
        RECT 54.950 11.550 57.050 11.900 ;
      LAYER met1 ;
        RECT 57.050 11.550 63.350 11.900 ;
      LAYER met1 ;
        RECT 63.350 11.550 65.800 11.900 ;
      LAYER met1 ;
        RECT 65.800 11.550 69.300 11.900 ;
      LAYER met1 ;
        RECT 69.300 11.550 71.750 11.900 ;
        RECT 36.050 11.200 44.800 11.550 ;
      LAYER met1 ;
        RECT 44.800 11.200 45.500 11.550 ;
      LAYER met1 ;
        RECT 45.500 11.200 51.800 11.550 ;
      LAYER met1 ;
        RECT 51.800 11.200 54.250 11.550 ;
      LAYER met1 ;
        RECT 54.250 11.200 57.400 11.550 ;
      LAYER met1 ;
        RECT 57.400 11.200 63.000 11.550 ;
      LAYER met1 ;
        RECT 63.000 11.200 66.500 11.550 ;
      LAYER met1 ;
        RECT 66.500 11.200 68.600 11.550 ;
      LAYER met1 ;
        RECT 68.600 11.200 71.750 11.550 ;
        RECT 24.500 10.850 29.750 11.200 ;
      LAYER met1 ;
        RECT 29.750 10.850 31.850 11.200 ;
      LAYER met1 ;
        RECT 31.850 10.850 33.600 11.200 ;
      LAYER met1 ;
        RECT 33.600 10.850 35.700 11.200 ;
      LAYER met1 ;
        RECT 35.700 10.850 71.750 11.200 ;
        RECT 19.600 10.500 20.300 10.850 ;
      LAYER met1 ;
        RECT 20.300 10.500 26.250 10.850 ;
      LAYER met1 ;
        RECT 26.250 10.500 30.100 10.850 ;
      LAYER met1 ;
        RECT 30.100 10.500 32.200 10.850 ;
      LAYER met1 ;
        RECT 32.200 10.500 33.250 10.850 ;
      LAYER met1 ;
        RECT 33.250 10.500 35.350 10.850 ;
      LAYER met1 ;
        RECT 35.350 10.500 71.750 10.850 ;
        RECT 19.600 10.150 19.950 10.500 ;
      LAYER met1 ;
        RECT 19.950 10.150 26.600 10.500 ;
      LAYER met1 ;
        RECT 26.600 10.150 30.450 10.500 ;
      LAYER met1 ;
        RECT 30.450 10.150 35.000 10.500 ;
      LAYER met1 ;
        RECT 35.000 10.150 71.750 10.500 ;
        RECT 19.600 9.800 20.300 10.150 ;
      LAYER met1 ;
        RECT 20.300 9.800 26.250 10.150 ;
      LAYER met1 ;
        RECT 26.250 9.800 31.150 10.150 ;
      LAYER met1 ;
        RECT 31.150 9.800 34.300 10.150 ;
      LAYER met1 ;
        RECT 34.300 9.800 71.750 10.150 ;
        RECT 19.600 9.450 45.850 9.800 ;
      LAYER met1 ;
        RECT 0.350 7.350 2.100 7.700 ;
      LAYER met1 ;
        RECT 0.000 6.300 0.700 7.350 ;
      LAYER met1 ;
        RECT 0.700 7.000 2.100 7.350 ;
      LAYER met1 ;
        RECT 2.100 7.000 5.950 7.700 ;
      LAYER met1 ;
        RECT 5.950 7.000 8.750 8.750 ;
      LAYER met1 ;
        RECT 8.750 7.000 10.500 8.750 ;
      LAYER met1 ;
        RECT 0.700 6.300 2.450 7.000 ;
      LAYER met1 ;
        RECT 2.450 6.300 10.500 7.000 ;
        RECT 0.000 5.600 1.050 6.300 ;
      LAYER met1 ;
        RECT 1.050 5.600 2.800 6.300 ;
      LAYER met1 ;
        RECT 2.800 5.600 10.500 6.300 ;
        RECT 0.000 5.250 1.400 5.600 ;
      LAYER met1 ;
        RECT 1.400 5.250 3.150 5.600 ;
      LAYER met1 ;
        RECT 3.150 5.250 10.500 5.600 ;
        RECT 0.000 4.550 1.750 5.250 ;
      LAYER met1 ;
        RECT 1.750 4.900 3.500 5.250 ;
      LAYER met1 ;
        RECT 3.500 4.900 10.500 5.250 ;
      LAYER met1 ;
        RECT 1.750 4.550 3.850 4.900 ;
      LAYER met1 ;
        RECT 3.850 4.550 10.500 4.900 ;
        RECT 0.000 4.200 2.100 4.550 ;
      LAYER met1 ;
        RECT 2.100 4.200 4.200 4.550 ;
      LAYER met1 ;
        RECT 4.200 4.200 10.500 4.550 ;
        RECT 0.000 3.850 2.450 4.200 ;
      LAYER met1 ;
        RECT 2.450 3.850 4.550 4.200 ;
      LAYER met1 ;
        RECT 4.550 3.850 10.500 4.200 ;
        RECT 0.000 3.500 2.800 3.850 ;
      LAYER met1 ;
        RECT 2.800 3.500 4.900 3.850 ;
      LAYER met1 ;
        RECT 4.900 3.500 10.500 3.850 ;
        RECT 0.000 3.150 3.150 3.500 ;
      LAYER met1 ;
        RECT 3.150 3.150 5.600 3.500 ;
      LAYER met1 ;
        RECT 5.600 3.150 10.500 3.500 ;
        RECT 0.000 2.800 3.500 3.150 ;
      LAYER met1 ;
        RECT 3.500 2.800 6.300 3.150 ;
      LAYER met1 ;
        RECT 6.300 2.800 10.500 3.150 ;
        RECT 0.000 2.450 3.850 2.800 ;
      LAYER met1 ;
        RECT 3.850 2.450 7.000 2.800 ;
      LAYER met1 ;
        RECT 7.000 2.450 10.500 2.800 ;
        RECT 0.000 2.100 4.550 2.450 ;
      LAYER met1 ;
        RECT 4.550 2.100 8.400 2.450 ;
      LAYER met1 ;
        RECT 8.400 2.100 10.500 2.450 ;
      LAYER met1 ;
        RECT 10.500 2.100 13.300 8.750 ;
      LAYER met1 ;
        RECT 13.300 8.050 17.850 8.750 ;
      LAYER met1 ;
        RECT 17.850 8.050 19.250 9.450 ;
      LAYER met1 ;
        RECT 19.250 8.400 45.850 9.450 ;
      LAYER met1 ;
        RECT 45.850 8.400 51.800 9.800 ;
      LAYER met1 ;
        RECT 19.250 8.050 49.700 8.400 ;
      LAYER met1 ;
        RECT 49.700 8.050 51.800 8.400 ;
      LAYER met1 ;
        RECT 51.800 8.050 52.850 9.800 ;
      LAYER met1 ;
        RECT 52.850 8.400 58.800 9.800 ;
      LAYER met1 ;
        RECT 58.800 8.400 59.500 9.800 ;
      LAYER met1 ;
        RECT 52.850 8.050 54.600 8.400 ;
      LAYER met1 ;
        RECT 54.600 8.050 59.500 8.400 ;
        RECT 13.300 7.350 17.500 8.050 ;
      LAYER met1 ;
        RECT 17.500 7.700 19.250 8.050 ;
      LAYER met1 ;
        RECT 19.250 7.700 50.050 8.050 ;
      LAYER met1 ;
        RECT 17.500 7.350 18.900 7.700 ;
      LAYER met1 ;
        RECT 18.900 7.350 50.050 7.700 ;
        RECT 13.300 6.300 17.150 7.350 ;
      LAYER met1 ;
        RECT 17.150 6.650 18.900 7.350 ;
      LAYER met1 ;
        RECT 18.900 7.000 21.000 7.350 ;
      LAYER met1 ;
        RECT 21.000 7.000 22.750 7.350 ;
      LAYER met1 ;
        RECT 22.750 7.000 25.550 7.350 ;
      LAYER met1 ;
        RECT 25.550 7.000 26.950 7.350 ;
      LAYER met1 ;
        RECT 26.950 7.000 29.400 7.350 ;
      LAYER met1 ;
        RECT 29.400 7.000 31.150 7.350 ;
      LAYER met1 ;
        RECT 31.150 7.000 33.250 7.350 ;
        RECT 18.900 6.650 20.300 7.000 ;
      LAYER met1 ;
        RECT 20.300 6.650 23.100 7.000 ;
      LAYER met1 ;
        RECT 23.100 6.650 25.200 7.000 ;
      LAYER met1 ;
        RECT 25.200 6.650 27.300 7.000 ;
      LAYER met1 ;
        RECT 27.300 6.650 29.050 7.000 ;
      LAYER met1 ;
        RECT 29.050 6.650 31.850 7.000 ;
        RECT 17.150 6.300 18.550 6.650 ;
      LAYER met1 ;
        RECT 18.550 6.300 20.300 6.650 ;
      LAYER met1 ;
        RECT 20.300 6.300 21.350 6.650 ;
      LAYER met1 ;
        RECT 21.350 6.300 22.050 6.650 ;
      LAYER met1 ;
        RECT 22.050 6.300 23.450 6.650 ;
      LAYER met1 ;
        RECT 13.300 5.950 16.800 6.300 ;
      LAYER met1 ;
        RECT 16.800 5.950 18.550 6.300 ;
      LAYER met1 ;
        RECT 18.550 5.950 22.400 6.300 ;
        RECT 13.300 5.250 16.450 5.950 ;
      LAYER met1 ;
        RECT 16.450 5.250 18.200 5.950 ;
      LAYER met1 ;
        RECT 18.200 5.250 22.400 5.950 ;
        RECT 13.300 4.900 16.100 5.250 ;
      LAYER met1 ;
        RECT 16.100 4.900 17.850 5.250 ;
      LAYER met1 ;
        RECT 17.850 4.900 22.400 5.250 ;
      LAYER met1 ;
        RECT 22.400 4.900 23.450 6.300 ;
      LAYER met1 ;
        RECT 23.450 5.600 24.850 6.650 ;
      LAYER met1 ;
        RECT 24.850 6.300 27.650 6.650 ;
      LAYER met1 ;
        RECT 27.650 6.300 29.050 6.650 ;
      LAYER met1 ;
        RECT 29.050 6.300 29.750 6.650 ;
      LAYER met1 ;
        RECT 29.750 6.300 30.450 6.650 ;
      LAYER met1 ;
        RECT 30.450 6.300 31.850 6.650 ;
      LAYER met1 ;
        RECT 31.850 6.300 33.250 7.000 ;
      LAYER met1 ;
        RECT 33.250 6.300 36.050 7.350 ;
      LAYER met1 ;
        RECT 36.050 6.300 50.050 7.350 ;
      LAYER met1 ;
        RECT 24.850 5.600 25.900 6.300 ;
      LAYER met1 ;
        RECT 25.900 5.950 26.600 6.300 ;
      LAYER met1 ;
        RECT 26.600 5.950 27.650 6.300 ;
      LAYER met1 ;
        RECT 27.650 5.950 30.800 6.300 ;
      LAYER met1 ;
        RECT 30.800 5.950 32.200 6.300 ;
      LAYER met1 ;
        RECT 25.900 5.600 26.950 5.950 ;
        RECT 23.450 4.900 24.500 5.600 ;
        RECT 13.300 4.550 15.750 4.900 ;
      LAYER met1 ;
        RECT 15.750 4.550 17.500 4.900 ;
      LAYER met1 ;
        RECT 17.500 4.550 22.050 4.900 ;
      LAYER met1 ;
        RECT 22.050 4.550 23.100 4.900 ;
      LAYER met1 ;
        RECT 23.100 4.550 24.500 4.900 ;
        RECT 13.300 4.200 15.400 4.550 ;
      LAYER met1 ;
        RECT 15.400 4.200 17.500 4.550 ;
      LAYER met1 ;
        RECT 17.500 4.200 21.700 4.550 ;
      LAYER met1 ;
        RECT 21.700 4.200 22.750 4.550 ;
      LAYER met1 ;
        RECT 22.750 4.200 24.500 4.550 ;
        RECT 13.300 3.850 15.050 4.200 ;
      LAYER met1 ;
        RECT 15.050 3.850 17.150 4.200 ;
      LAYER met1 ;
        RECT 17.150 3.850 21.350 4.200 ;
      LAYER met1 ;
        RECT 21.350 3.850 22.400 4.200 ;
      LAYER met1 ;
        RECT 22.400 3.850 24.500 4.200 ;
      LAYER met1 ;
        RECT 24.500 3.850 25.550 5.600 ;
      LAYER met1 ;
        RECT 25.550 4.900 26.950 5.600 ;
        RECT 25.550 4.200 25.900 4.900 ;
      LAYER met1 ;
        RECT 25.900 4.200 26.600 4.900 ;
      LAYER met1 ;
        RECT 26.600 4.200 26.950 4.900 ;
        RECT 13.300 3.500 14.350 3.850 ;
      LAYER met1 ;
        RECT 14.350 3.500 16.800 3.850 ;
      LAYER met1 ;
        RECT 16.800 3.500 21.000 3.850 ;
      LAYER met1 ;
        RECT 21.000 3.500 22.050 3.850 ;
      LAYER met1 ;
        RECT 22.050 3.500 24.850 3.850 ;
      LAYER met1 ;
        RECT 24.850 3.500 25.550 3.850 ;
      LAYER met1 ;
        RECT 25.550 3.500 26.950 4.200 ;
        RECT 0.000 1.750 4.900 2.100 ;
      LAYER met1 ;
        RECT 4.900 1.750 13.300 2.100 ;
      LAYER met1 ;
        RECT 13.300 1.750 14.000 3.500 ;
      LAYER met1 ;
        RECT 14.000 3.150 16.450 3.500 ;
      LAYER met1 ;
        RECT 16.450 3.150 20.650 3.500 ;
      LAYER met1 ;
        RECT 20.650 3.150 21.700 3.500 ;
      LAYER met1 ;
        RECT 21.700 3.150 24.850 3.500 ;
      LAYER met1 ;
        RECT 14.000 2.800 16.100 3.150 ;
      LAYER met1 ;
        RECT 16.100 2.800 20.300 3.150 ;
      LAYER met1 ;
        RECT 14.000 2.450 15.750 2.800 ;
      LAYER met1 ;
        RECT 15.750 2.450 20.300 2.800 ;
      LAYER met1 ;
        RECT 14.000 2.100 15.050 2.450 ;
      LAYER met1 ;
        RECT 15.050 2.100 20.300 2.450 ;
      LAYER met1 ;
        RECT 20.300 2.100 23.450 3.150 ;
      LAYER met1 ;
        RECT 23.450 2.800 24.850 3.150 ;
      LAYER met1 ;
        RECT 24.850 2.800 25.900 3.500 ;
      LAYER met1 ;
        RECT 25.900 3.150 26.950 3.500 ;
      LAYER met1 ;
        RECT 26.950 3.150 28.000 5.950 ;
      LAYER met1 ;
        RECT 28.000 5.600 31.150 5.950 ;
      LAYER met1 ;
        RECT 31.150 5.600 32.200 5.950 ;
      LAYER met1 ;
        RECT 32.200 5.600 33.250 6.300 ;
      LAYER met1 ;
        RECT 33.250 5.600 34.300 6.300 ;
      LAYER met1 ;
        RECT 34.300 5.600 50.050 6.300 ;
        RECT 28.000 4.900 30.800 5.600 ;
      LAYER met1 ;
        RECT 30.800 4.900 31.850 5.600 ;
      LAYER met1 ;
        RECT 31.850 4.900 33.250 5.600 ;
      LAYER met1 ;
        RECT 33.250 5.250 35.000 5.600 ;
      LAYER met1 ;
        RECT 35.000 5.250 50.050 5.600 ;
      LAYER met1 ;
        RECT 33.250 4.900 35.700 5.250 ;
      LAYER met1 ;
        RECT 35.700 4.900 50.050 5.250 ;
        RECT 28.000 4.550 30.450 4.900 ;
      LAYER met1 ;
        RECT 30.450 4.550 31.500 4.900 ;
      LAYER met1 ;
        RECT 31.500 4.550 33.250 4.900 ;
      LAYER met1 ;
        RECT 33.250 4.550 36.050 4.900 ;
      LAYER met1 ;
        RECT 36.050 4.550 50.050 4.900 ;
        RECT 28.000 4.200 30.100 4.550 ;
      LAYER met1 ;
        RECT 30.100 4.200 31.150 4.550 ;
      LAYER met1 ;
        RECT 31.150 4.200 35.000 4.550 ;
      LAYER met1 ;
        RECT 35.000 4.200 36.400 4.550 ;
      LAYER met1 ;
        RECT 28.000 3.850 29.750 4.200 ;
      LAYER met1 ;
        RECT 29.750 3.850 30.800 4.200 ;
      LAYER met1 ;
        RECT 30.800 3.850 35.350 4.200 ;
        RECT 28.000 3.500 29.400 3.850 ;
      LAYER met1 ;
        RECT 29.400 3.500 30.450 3.850 ;
      LAYER met1 ;
        RECT 30.450 3.500 35.350 3.850 ;
        RECT 28.000 3.150 29.050 3.500 ;
      LAYER met1 ;
        RECT 29.050 3.150 30.100 3.500 ;
      LAYER met1 ;
        RECT 30.100 3.150 35.350 3.500 ;
      LAYER met1 ;
        RECT 35.350 3.150 36.400 4.200 ;
      LAYER met1 ;
        RECT 36.400 3.850 50.050 4.550 ;
        RECT 25.900 2.800 26.600 3.150 ;
      LAYER met1 ;
        RECT 26.600 2.800 27.650 3.150 ;
      LAYER met1 ;
        RECT 23.450 2.450 25.200 2.800 ;
      LAYER met1 ;
        RECT 25.200 2.450 27.650 2.800 ;
      LAYER met1 ;
        RECT 27.650 2.450 28.700 3.150 ;
      LAYER met1 ;
        RECT 28.700 2.800 31.850 3.150 ;
      LAYER met1 ;
        RECT 31.850 2.800 33.250 3.150 ;
      LAYER met1 ;
        RECT 33.250 2.800 33.600 3.150 ;
      LAYER met1 ;
        RECT 33.600 2.800 35.000 3.150 ;
      LAYER met1 ;
        RECT 35.000 2.800 36.400 3.150 ;
      LAYER met1 ;
        RECT 36.400 2.800 45.850 3.850 ;
      LAYER met1 ;
        RECT 45.850 3.500 47.250 3.850 ;
      LAYER met1 ;
        RECT 47.250 3.500 50.050 3.850 ;
        RECT 23.450 2.100 25.550 2.450 ;
      LAYER met1 ;
        RECT 25.550 2.100 27.300 2.450 ;
      LAYER met1 ;
        RECT 27.300 2.100 28.700 2.450 ;
      LAYER met1 ;
        RECT 28.700 2.100 32.200 2.800 ;
      LAYER met1 ;
        RECT 32.200 2.100 33.250 2.800 ;
      LAYER met1 ;
        RECT 33.250 2.450 36.050 2.800 ;
      LAYER met1 ;
        RECT 36.050 2.450 45.850 2.800 ;
      LAYER met1 ;
        RECT 33.250 2.100 35.700 2.450 ;
      LAYER met1 ;
        RECT 35.700 2.100 45.850 2.450 ;
      LAYER met1 ;
        RECT 14.000 1.750 14.350 2.100 ;
      LAYER met1 ;
        RECT 14.350 1.750 45.850 2.100 ;
      LAYER met1 ;
        RECT 45.850 1.750 47.600 3.500 ;
      LAYER met1 ;
        RECT 47.600 1.750 50.050 3.500 ;
      LAYER met1 ;
        RECT 50.050 1.750 51.450 8.050 ;
      LAYER met1 ;
        RECT 51.450 3.850 52.850 8.050 ;
      LAYER met1 ;
        RECT 52.850 5.600 54.250 8.050 ;
      LAYER met1 ;
        RECT 54.250 5.600 59.500 8.050 ;
      LAYER met1 ;
        RECT 59.500 6.650 61.250 9.800 ;
      LAYER met1 ;
        RECT 61.250 9.450 64.400 9.800 ;
      LAYER met1 ;
        RECT 64.400 9.450 65.100 9.800 ;
      LAYER met1 ;
        RECT 65.100 9.450 71.750 9.800 ;
        RECT 61.250 9.100 64.050 9.450 ;
      LAYER met1 ;
        RECT 64.050 9.100 65.450 9.450 ;
      LAYER met1 ;
        RECT 65.450 9.100 71.750 9.450 ;
        RECT 61.250 8.750 63.700 9.100 ;
      LAYER met1 ;
        RECT 63.700 8.750 65.800 9.100 ;
      LAYER met1 ;
        RECT 65.800 8.750 71.750 9.100 ;
        RECT 61.250 8.400 63.350 8.750 ;
      LAYER met1 ;
        RECT 63.350 8.400 65.450 8.750 ;
      LAYER met1 ;
        RECT 65.450 8.400 71.750 8.750 ;
        RECT 61.250 8.050 63.000 8.400 ;
      LAYER met1 ;
        RECT 63.000 8.050 65.100 8.400 ;
      LAYER met1 ;
        RECT 65.100 8.050 71.750 8.400 ;
        RECT 61.250 7.700 62.650 8.050 ;
      LAYER met1 ;
        RECT 62.650 7.700 64.750 8.050 ;
      LAYER met1 ;
        RECT 64.750 7.700 71.750 8.050 ;
        RECT 61.250 7.350 62.300 7.700 ;
      LAYER met1 ;
        RECT 62.300 7.350 64.400 7.700 ;
      LAYER met1 ;
        RECT 61.250 7.000 61.950 7.350 ;
      LAYER met1 ;
        RECT 61.950 7.000 64.400 7.350 ;
      LAYER met1 ;
        RECT 64.400 7.000 71.750 7.700 ;
        RECT 61.250 6.650 61.600 7.000 ;
      LAYER met1 ;
        RECT 61.600 6.650 64.050 7.000 ;
      LAYER met1 ;
        RECT 64.050 6.650 71.750 7.000 ;
      LAYER met1 ;
        RECT 59.500 6.300 63.700 6.650 ;
      LAYER met1 ;
        RECT 63.700 6.300 71.750 6.650 ;
      LAYER met1 ;
        RECT 59.500 5.950 63.350 6.300 ;
      LAYER met1 ;
        RECT 63.350 5.950 71.750 6.300 ;
      LAYER met1 ;
        RECT 59.500 5.600 63.000 5.950 ;
      LAYER met1 ;
        RECT 63.000 5.600 71.750 5.950 ;
      LAYER met1 ;
        RECT 52.850 5.250 54.600 5.600 ;
      LAYER met1 ;
        RECT 54.600 5.250 59.500 5.600 ;
      LAYER met1 ;
        RECT 59.500 5.250 62.650 5.600 ;
      LAYER met1 ;
        RECT 62.650 5.250 71.750 5.600 ;
      LAYER met1 ;
        RECT 52.850 3.850 58.800 5.250 ;
      LAYER met1 ;
        RECT 51.450 1.750 57.050 3.850 ;
      LAYER met1 ;
        RECT 57.050 1.750 58.800 3.850 ;
      LAYER met1 ;
        RECT 0.000 1.400 5.600 1.750 ;
      LAYER met1 ;
        RECT 5.600 1.400 13.300 1.750 ;
      LAYER met1 ;
        RECT 13.300 1.400 45.850 1.750 ;
        RECT 0.000 1.050 6.650 1.400 ;
      LAYER met1 ;
        RECT 6.650 1.050 12.950 1.400 ;
      LAYER met1 ;
        RECT 12.950 1.050 45.850 1.400 ;
        RECT 0.000 0.700 7.700 1.050 ;
      LAYER met1 ;
        RECT 7.700 0.700 11.900 1.050 ;
      LAYER met1 ;
        RECT 11.900 0.700 45.850 1.050 ;
        RECT 0.000 0.000 45.850 0.700 ;
      LAYER met1 ;
        RECT 45.850 0.000 51.450 1.750 ;
      LAYER met1 ;
        RECT 51.450 0.000 52.850 1.750 ;
      LAYER met1 ;
        RECT 52.850 0.000 58.800 1.750 ;
      LAYER met1 ;
        RECT 58.800 0.350 59.500 5.250 ;
      LAYER met1 ;
        RECT 59.500 4.900 62.300 5.250 ;
      LAYER met1 ;
        RECT 62.300 4.900 71.750 5.250 ;
      LAYER met1 ;
        RECT 59.500 4.200 62.650 4.900 ;
      LAYER met1 ;
        RECT 62.650 4.200 71.750 4.900 ;
      LAYER met1 ;
        RECT 59.500 3.850 63.000 4.200 ;
      LAYER met1 ;
        RECT 63.000 3.850 71.750 4.200 ;
      LAYER met1 ;
        RECT 59.500 3.500 63.350 3.850 ;
      LAYER met1 ;
        RECT 63.350 3.500 71.750 3.850 ;
      LAYER met1 ;
        RECT 59.500 0.350 61.250 3.500 ;
      LAYER met1 ;
        RECT 61.250 3.150 61.600 3.500 ;
      LAYER met1 ;
        RECT 61.600 3.150 63.700 3.500 ;
      LAYER met1 ;
        RECT 63.700 3.150 71.750 3.500 ;
        RECT 61.250 2.800 61.950 3.150 ;
      LAYER met1 ;
        RECT 61.950 2.800 64.050 3.150 ;
      LAYER met1 ;
        RECT 64.050 2.800 71.750 3.150 ;
        RECT 61.250 2.450 62.300 2.800 ;
      LAYER met1 ;
        RECT 62.300 2.450 64.400 2.800 ;
      LAYER met1 ;
        RECT 64.400 2.450 71.750 2.800 ;
        RECT 61.250 1.750 62.650 2.450 ;
      LAYER met1 ;
        RECT 62.650 2.100 64.750 2.450 ;
      LAYER met1 ;
        RECT 64.750 2.100 71.750 2.450 ;
      LAYER met1 ;
        RECT 62.650 1.750 65.100 2.100 ;
      LAYER met1 ;
        RECT 65.100 1.750 71.750 2.100 ;
        RECT 61.250 1.400 63.000 1.750 ;
      LAYER met1 ;
        RECT 63.000 1.400 65.450 1.750 ;
      LAYER met1 ;
        RECT 65.450 1.400 71.750 1.750 ;
        RECT 61.250 1.050 63.350 1.400 ;
      LAYER met1 ;
        RECT 63.350 1.050 65.800 1.400 ;
      LAYER met1 ;
        RECT 65.800 1.050 71.750 1.400 ;
        RECT 61.250 0.700 63.700 1.050 ;
      LAYER met1 ;
        RECT 63.700 0.700 65.450 1.050 ;
      LAYER met1 ;
        RECT 61.250 0.350 64.050 0.700 ;
      LAYER met1 ;
        RECT 64.050 0.350 65.450 0.700 ;
      LAYER met1 ;
        RECT 65.450 0.350 71.750 1.050 ;
        RECT 58.800 0.000 59.850 0.350 ;
      LAYER met1 ;
        RECT 59.850 0.000 61.250 0.350 ;
      LAYER met1 ;
        RECT 61.250 0.000 64.400 0.350 ;
      LAYER met1 ;
        RECT 64.400 0.000 64.750 0.350 ;
      LAYER met1 ;
        RECT 64.750 0.000 71.750 0.350 ;
  END
END my_logo
END LIBRARY

