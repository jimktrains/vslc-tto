VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO jsk
  CLASS BLOCK ;
  FOREIGN jsk ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 15.120 ;
  OBS
      LAYER met1 ;
        RECT 0.000 14.840 11.760 15.120 ;
        RECT 0.000 14.560 2.520 14.840 ;
      LAYER met1 ;
        RECT 2.520 14.560 3.640 14.840 ;
      LAYER met1 ;
        RECT 3.640 14.560 5.040 14.840 ;
      LAYER met1 ;
        RECT 5.040 14.560 5.600 14.840 ;
      LAYER met1 ;
        RECT 5.600 14.560 7.000 14.840 ;
      LAYER met1 ;
        RECT 7.000 14.560 8.120 14.840 ;
      LAYER met1 ;
        RECT 8.120 14.560 8.960 14.840 ;
      LAYER met1 ;
        RECT 8.960 14.560 10.640 14.840 ;
      LAYER met1 ;
        RECT 0.000 14.000 2.240 14.560 ;
      LAYER met1 ;
        RECT 2.240 14.280 2.800 14.560 ;
      LAYER met1 ;
        RECT 2.800 14.280 3.360 14.560 ;
      LAYER met1 ;
        RECT 2.240 14.000 2.520 14.280 ;
      LAYER met1 ;
        RECT 2.520 14.000 3.360 14.280 ;
        RECT 0.000 13.440 3.360 14.000 ;
      LAYER met1 ;
        RECT 3.360 13.720 3.920 14.560 ;
      LAYER met1 ;
        RECT 3.920 14.000 4.760 14.560 ;
      LAYER met1 ;
        RECT 4.760 14.280 5.880 14.560 ;
        RECT 4.760 14.000 5.040 14.280 ;
      LAYER met1 ;
        RECT 5.040 14.000 5.600 14.280 ;
      LAYER met1 ;
        RECT 5.600 14.000 5.880 14.280 ;
      LAYER met1 ;
        RECT 5.880 14.000 6.720 14.560 ;
      LAYER met1 ;
        RECT 6.720 14.280 7.280 14.560 ;
      LAYER met1 ;
        RECT 7.280 14.280 7.840 14.560 ;
      LAYER met1 ;
        RECT 6.720 14.000 7.000 14.280 ;
      LAYER met1 ;
        RECT 7.000 14.000 7.840 14.280 ;
        RECT 3.920 13.720 4.480 14.000 ;
      LAYER met1 ;
        RECT 4.480 13.720 5.320 14.000 ;
      LAYER met1 ;
        RECT 5.320 13.720 5.600 14.000 ;
      LAYER met1 ;
        RECT 5.600 13.720 6.160 14.000 ;
        RECT 3.360 13.440 3.640 13.720 ;
      LAYER met1 ;
        RECT 0.000 13.160 3.080 13.440 ;
      LAYER met1 ;
        RECT 3.080 13.160 3.640 13.440 ;
      LAYER met1 ;
        RECT 3.640 13.160 4.480 13.720 ;
        RECT 0.000 12.600 2.800 13.160 ;
      LAYER met1 ;
        RECT 2.800 12.600 3.360 13.160 ;
      LAYER met1 ;
        RECT 3.360 12.600 4.480 13.160 ;
      LAYER met1 ;
        RECT 4.480 12.880 4.760 13.720 ;
      LAYER met1 ;
        RECT 4.760 13.160 5.040 13.720 ;
      LAYER met1 ;
        RECT 5.040 13.440 5.320 13.720 ;
      LAYER met1 ;
        RECT 5.320 13.440 5.880 13.720 ;
      LAYER met1 ;
        RECT 5.040 13.160 5.600 13.440 ;
      LAYER met1 ;
        RECT 4.760 12.880 5.320 13.160 ;
      LAYER met1 ;
        RECT 5.320 12.880 5.600 13.160 ;
      LAYER met1 ;
        RECT 5.600 12.880 5.880 13.440 ;
      LAYER met1 ;
        RECT 5.880 12.880 6.160 13.720 ;
      LAYER met1 ;
        RECT 6.160 13.440 7.840 14.000 ;
      LAYER met1 ;
        RECT 7.840 13.720 8.400 14.560 ;
      LAYER met1 ;
        RECT 8.400 13.720 8.960 14.560 ;
      LAYER met1 ;
        RECT 8.960 13.720 9.520 14.560 ;
      LAYER met1 ;
        RECT 9.520 14.280 10.080 14.560 ;
      LAYER met1 ;
        RECT 10.080 14.280 10.640 14.560 ;
      LAYER met1 ;
        RECT 10.640 14.280 11.760 14.840 ;
        RECT 9.520 13.720 11.760 14.280 ;
      LAYER met1 ;
        RECT 7.840 13.440 8.120 13.720 ;
      LAYER met1 ;
        RECT 8.120 13.440 8.960 13.720 ;
      LAYER met1 ;
        RECT 8.960 13.440 10.360 13.720 ;
      LAYER met1 ;
        RECT 10.360 13.440 11.760 13.720 ;
        RECT 6.160 13.160 7.560 13.440 ;
      LAYER met1 ;
        RECT 7.560 13.160 8.120 13.440 ;
      LAYER met1 ;
        RECT 8.120 13.160 10.080 13.440 ;
      LAYER met1 ;
        RECT 4.480 12.600 5.040 12.880 ;
      LAYER met1 ;
        RECT 5.040 12.600 5.320 12.880 ;
      LAYER met1 ;
        RECT 5.320 12.600 6.160 12.880 ;
      LAYER met1 ;
        RECT 6.160 12.600 7.280 13.160 ;
      LAYER met1 ;
        RECT 7.280 12.600 7.840 13.160 ;
      LAYER met1 ;
        RECT 7.840 12.600 10.080 13.160 ;
        RECT 0.000 12.040 2.520 12.600 ;
      LAYER met1 ;
        RECT 2.520 12.320 3.080 12.600 ;
      LAYER met1 ;
        RECT 3.080 12.320 4.760 12.600 ;
      LAYER met1 ;
        RECT 4.760 12.320 5.040 12.600 ;
      LAYER met1 ;
        RECT 5.040 12.320 5.600 12.600 ;
      LAYER met1 ;
        RECT 5.600 12.320 5.880 12.600 ;
        RECT 2.520 12.040 3.640 12.320 ;
      LAYER met1 ;
        RECT 3.640 12.040 4.760 12.320 ;
      LAYER met1 ;
        RECT 4.760 12.040 5.880 12.320 ;
      LAYER met1 ;
        RECT 5.880 12.040 7.000 12.600 ;
      LAYER met1 ;
        RECT 7.000 12.320 7.560 12.600 ;
      LAYER met1 ;
        RECT 7.560 12.320 8.960 12.600 ;
      LAYER met1 ;
        RECT 8.960 12.320 9.520 12.600 ;
      LAYER met1 ;
        RECT 9.520 12.320 10.080 12.600 ;
      LAYER met1 ;
        RECT 10.080 12.320 10.640 13.440 ;
      LAYER met1 ;
        RECT 10.640 12.320 11.760 13.440 ;
      LAYER met1 ;
        RECT 7.000 12.040 8.120 12.320 ;
      LAYER met1 ;
        RECT 8.120 12.040 8.960 12.320 ;
      LAYER met1 ;
        RECT 8.960 12.040 10.360 12.320 ;
      LAYER met1 ;
        RECT 0.000 11.760 2.240 12.040 ;
      LAYER met1 ;
        RECT 2.240 11.760 3.920 12.040 ;
      LAYER met1 ;
        RECT 3.920 11.760 5.040 12.040 ;
      LAYER met1 ;
        RECT 5.040 11.760 5.600 12.040 ;
      LAYER met1 ;
        RECT 5.600 11.760 6.720 12.040 ;
      LAYER met1 ;
        RECT 6.720 11.760 8.400 12.040 ;
      LAYER met1 ;
        RECT 8.400 11.760 9.240 12.040 ;
      LAYER met1 ;
        RECT 9.240 11.760 10.360 12.040 ;
      LAYER met1 ;
        RECT 10.360 11.760 11.760 12.320 ;
        RECT 0.000 11.200 11.760 11.760 ;
        RECT 0.000 10.080 1.120 11.200 ;
      LAYER met1 ;
        RECT 1.120 10.080 3.640 11.200 ;
      LAYER met1 ;
        RECT 3.640 10.080 11.760 11.200 ;
        RECT 0.000 7.280 1.680 10.080 ;
        RECT 0.000 7.000 0.280 7.280 ;
      LAYER met1 ;
        RECT 0.280 7.000 1.120 7.280 ;
      LAYER met1 ;
        RECT 1.120 7.000 1.680 7.280 ;
      LAYER met1 ;
        RECT 0.000 6.160 1.400 7.000 ;
      LAYER met1 ;
        RECT 1.400 6.160 1.680 7.000 ;
      LAYER met1 ;
        RECT 1.680 6.160 3.080 10.080 ;
      LAYER met1 ;
        RECT 3.080 9.240 4.200 10.080 ;
      LAYER met1 ;
        RECT 4.200 9.240 7.280 10.080 ;
      LAYER met1 ;
        RECT 7.280 9.240 11.760 10.080 ;
        RECT 3.080 7.560 3.640 9.240 ;
      LAYER met1 ;
        RECT 3.640 8.960 7.560 9.240 ;
        RECT 3.640 7.560 5.040 8.960 ;
      LAYER met1 ;
        RECT 5.040 8.400 6.160 8.960 ;
      LAYER met1 ;
        RECT 6.160 8.400 7.560 8.960 ;
      LAYER met1 ;
        RECT 5.040 8.120 6.440 8.400 ;
      LAYER met1 ;
        RECT 6.440 8.120 7.560 8.400 ;
      LAYER met1 ;
        RECT 7.560 8.120 8.120 9.240 ;
        RECT 5.040 7.560 8.120 8.120 ;
        RECT 3.080 7.280 3.920 7.560 ;
      LAYER met1 ;
        RECT 3.920 7.280 7.280 7.560 ;
      LAYER met1 ;
        RECT 3.080 6.440 4.200 7.280 ;
      LAYER met1 ;
        RECT 4.200 6.720 7.280 7.280 ;
      LAYER met1 ;
        RECT 7.280 6.720 8.120 7.560 ;
      LAYER met1 ;
        RECT 8.120 6.720 9.520 9.240 ;
      LAYER met1 ;
        RECT 9.520 8.400 10.640 9.240 ;
      LAYER met1 ;
        RECT 10.640 8.400 11.760 9.240 ;
      LAYER met1 ;
        RECT 9.520 7.560 10.360 8.400 ;
      LAYER met1 ;
        RECT 10.360 7.560 11.760 8.400 ;
      LAYER met1 ;
        RECT 9.520 6.720 9.800 7.560 ;
      LAYER met1 ;
        RECT 9.800 7.280 11.760 7.560 ;
        RECT 9.800 6.720 11.200 7.280 ;
        RECT 4.200 6.440 7.560 6.720 ;
      LAYER met1 ;
        RECT 3.080 6.160 6.160 6.440 ;
        RECT 0.000 5.880 0.280 6.160 ;
      LAYER met1 ;
        RECT 0.280 5.880 3.080 6.160 ;
      LAYER met1 ;
        RECT 3.080 5.880 3.920 6.160 ;
      LAYER met1 ;
        RECT 3.920 5.880 4.760 6.160 ;
      LAYER met1 ;
        RECT 4.760 5.880 6.160 6.160 ;
        RECT 0.000 5.040 0.560 5.880 ;
      LAYER met1 ;
        RECT 0.560 5.320 2.800 5.880 ;
      LAYER met1 ;
        RECT 2.800 5.320 3.640 5.880 ;
      LAYER met1 ;
        RECT 0.560 5.040 2.520 5.320 ;
      LAYER met1 ;
        RECT 2.520 5.040 3.640 5.320 ;
      LAYER met1 ;
        RECT 3.640 5.040 5.040 5.880 ;
      LAYER met1 ;
        RECT 5.040 5.040 6.160 5.880 ;
      LAYER met1 ;
        RECT 6.160 5.040 7.560 6.440 ;
      LAYER met1 ;
        RECT 0.000 4.760 3.920 5.040 ;
      LAYER met1 ;
        RECT 3.920 4.760 7.560 5.040 ;
      LAYER met1 ;
        RECT 7.560 4.760 8.120 6.720 ;
      LAYER met1 ;
        RECT 8.120 6.440 11.200 6.720 ;
      LAYER met1 ;
        RECT 11.200 6.440 11.760 7.280 ;
      LAYER met1 ;
        RECT 8.120 5.880 10.640 6.440 ;
      LAYER met1 ;
        RECT 10.640 5.880 11.760 6.440 ;
      LAYER met1 ;
        RECT 8.120 5.600 11.200 5.880 ;
      LAYER met1 ;
        RECT 0.000 3.920 4.200 4.760 ;
      LAYER met1 ;
        RECT 4.200 4.200 7.280 4.760 ;
      LAYER met1 ;
        RECT 7.280 4.200 8.120 4.760 ;
      LAYER met1 ;
        RECT 4.200 3.920 7.000 4.200 ;
      LAYER met1 ;
        RECT 7.000 3.920 8.120 4.200 ;
        RECT 0.000 3.360 8.120 3.920 ;
      LAYER met1 ;
        RECT 8.120 3.360 9.520 5.600 ;
      LAYER met1 ;
        RECT 9.520 4.760 9.800 5.600 ;
      LAYER met1 ;
        RECT 9.800 5.040 11.200 5.600 ;
      LAYER met1 ;
        RECT 11.200 5.040 11.760 5.880 ;
      LAYER met1 ;
        RECT 9.800 4.760 11.760 5.040 ;
      LAYER met1 ;
        RECT 9.520 3.920 10.360 4.760 ;
      LAYER met1 ;
        RECT 10.360 3.920 11.760 4.760 ;
      LAYER met1 ;
        RECT 9.520 3.360 10.640 3.920 ;
      LAYER met1 ;
        RECT 10.640 3.360 11.760 3.920 ;
      LAYER met1 ;
        RECT 0.000 3.080 8.400 3.360 ;
      LAYER met1 ;
        RECT 8.400 3.080 9.520 3.360 ;
      LAYER met1 ;
        RECT 9.520 3.080 10.920 3.360 ;
      LAYER met1 ;
        RECT 10.920 3.080 11.760 3.360 ;
      LAYER met1 ;
        RECT 0.000 2.800 11.760 3.080 ;
        RECT 0.000 2.240 2.240 2.800 ;
      LAYER met1 ;
        RECT 2.240 2.240 5.880 2.800 ;
      LAYER met1 ;
        RECT 5.880 2.520 6.720 2.800 ;
      LAYER met1 ;
        RECT 6.720 2.520 7.280 2.800 ;
      LAYER met1 ;
        RECT 7.280 2.520 8.680 2.800 ;
      LAYER met1 ;
        RECT 8.680 2.520 9.240 2.800 ;
      LAYER met1 ;
        RECT 9.240 2.520 11.760 2.800 ;
        RECT 5.880 2.240 6.440 2.520 ;
        RECT 0.000 0.000 2.800 2.240 ;
      LAYER met1 ;
        RECT 2.800 0.000 3.360 2.240 ;
      LAYER met1 ;
        RECT 3.360 0.000 4.760 2.240 ;
      LAYER met1 ;
        RECT 4.760 0.000 5.320 2.240 ;
      LAYER met1 ;
        RECT 5.320 1.960 6.440 2.240 ;
      LAYER met1 ;
        RECT 6.440 1.960 7.280 2.520 ;
      LAYER met1 ;
        RECT 7.280 1.960 8.400 2.520 ;
      LAYER met1 ;
        RECT 8.400 2.240 9.520 2.520 ;
        RECT 8.400 1.960 8.680 2.240 ;
      LAYER met1 ;
        RECT 8.680 1.960 9.240 2.240 ;
      LAYER met1 ;
        RECT 9.240 1.960 9.520 2.240 ;
      LAYER met1 ;
        RECT 9.520 1.960 11.760 2.520 ;
        RECT 5.320 0.280 6.720 1.960 ;
      LAYER met1 ;
        RECT 6.720 0.280 7.280 1.960 ;
      LAYER met1 ;
        RECT 7.280 0.560 8.120 1.960 ;
      LAYER met1 ;
        RECT 8.120 1.680 8.960 1.960 ;
      LAYER met1 ;
        RECT 8.960 1.680 9.240 1.960 ;
      LAYER met1 ;
        RECT 9.240 1.680 9.800 1.960 ;
        RECT 8.120 0.840 8.400 1.680 ;
      LAYER met1 ;
        RECT 8.400 1.120 8.680 1.680 ;
      LAYER met1 ;
        RECT 8.680 1.400 8.960 1.680 ;
      LAYER met1 ;
        RECT 8.960 1.400 9.520 1.680 ;
      LAYER met1 ;
        RECT 8.680 1.120 9.240 1.400 ;
      LAYER met1 ;
        RECT 8.400 0.840 8.960 1.120 ;
      LAYER met1 ;
        RECT 8.960 0.840 9.240 1.120 ;
      LAYER met1 ;
        RECT 9.240 0.840 9.520 1.400 ;
      LAYER met1 ;
        RECT 9.520 0.840 9.800 1.680 ;
        RECT 8.120 0.560 8.680 0.840 ;
      LAYER met1 ;
        RECT 8.680 0.560 8.960 0.840 ;
      LAYER met1 ;
        RECT 8.960 0.560 9.800 0.840 ;
      LAYER met1 ;
        RECT 9.800 0.560 11.760 1.960 ;
        RECT 7.280 0.280 8.400 0.560 ;
      LAYER met1 ;
        RECT 8.400 0.280 8.680 0.560 ;
      LAYER met1 ;
        RECT 8.680 0.280 9.240 0.560 ;
      LAYER met1 ;
        RECT 9.240 0.280 9.520 0.560 ;
      LAYER met1 ;
        RECT 5.320 0.000 6.160 0.280 ;
      LAYER met1 ;
        RECT 6.160 0.000 7.840 0.280 ;
      LAYER met1 ;
        RECT 7.840 0.000 8.400 0.280 ;
      LAYER met1 ;
        RECT 8.400 0.000 9.520 0.280 ;
      LAYER met1 ;
        RECT 9.520 0.000 11.760 0.560 ;
      LAYER met2 ;
        RECT 0.000 14.840 11.760 15.120 ;
        RECT 0.000 14.560 2.520 14.840 ;
      LAYER met2 ;
        RECT 2.520 14.560 3.640 14.840 ;
      LAYER met2 ;
        RECT 3.640 14.560 5.040 14.840 ;
      LAYER met2 ;
        RECT 5.040 14.560 5.600 14.840 ;
      LAYER met2 ;
        RECT 5.600 14.560 7.000 14.840 ;
      LAYER met2 ;
        RECT 7.000 14.560 8.120 14.840 ;
      LAYER met2 ;
        RECT 8.120 14.560 8.960 14.840 ;
      LAYER met2 ;
        RECT 8.960 14.560 10.640 14.840 ;
      LAYER met2 ;
        RECT 0.000 14.000 2.240 14.560 ;
      LAYER met2 ;
        RECT 2.240 14.280 2.800 14.560 ;
      LAYER met2 ;
        RECT 2.800 14.280 3.360 14.560 ;
      LAYER met2 ;
        RECT 2.240 14.000 2.520 14.280 ;
      LAYER met2 ;
        RECT 2.520 14.000 3.360 14.280 ;
        RECT 0.000 13.440 3.360 14.000 ;
      LAYER met2 ;
        RECT 3.360 13.720 3.920 14.560 ;
      LAYER met2 ;
        RECT 3.920 14.000 4.760 14.560 ;
      LAYER met2 ;
        RECT 4.760 14.280 5.880 14.560 ;
        RECT 4.760 14.000 5.040 14.280 ;
      LAYER met2 ;
        RECT 5.040 14.000 5.600 14.280 ;
      LAYER met2 ;
        RECT 5.600 14.000 5.880 14.280 ;
      LAYER met2 ;
        RECT 5.880 14.000 6.720 14.560 ;
      LAYER met2 ;
        RECT 6.720 14.280 7.280 14.560 ;
      LAYER met2 ;
        RECT 7.280 14.280 7.840 14.560 ;
      LAYER met2 ;
        RECT 6.720 14.000 7.000 14.280 ;
      LAYER met2 ;
        RECT 7.000 14.000 7.840 14.280 ;
        RECT 3.920 13.720 4.480 14.000 ;
      LAYER met2 ;
        RECT 4.480 13.720 5.320 14.000 ;
      LAYER met2 ;
        RECT 5.320 13.720 5.600 14.000 ;
      LAYER met2 ;
        RECT 5.600 13.720 6.160 14.000 ;
        RECT 3.360 13.440 3.640 13.720 ;
      LAYER met2 ;
        RECT 0.000 13.160 3.080 13.440 ;
      LAYER met2 ;
        RECT 3.080 13.160 3.640 13.440 ;
      LAYER met2 ;
        RECT 3.640 13.160 4.480 13.720 ;
        RECT 0.000 12.600 2.800 13.160 ;
      LAYER met2 ;
        RECT 2.800 12.600 3.360 13.160 ;
      LAYER met2 ;
        RECT 3.360 12.600 4.480 13.160 ;
      LAYER met2 ;
        RECT 4.480 12.880 4.760 13.720 ;
      LAYER met2 ;
        RECT 4.760 13.160 5.040 13.720 ;
      LAYER met2 ;
        RECT 5.040 13.440 5.320 13.720 ;
      LAYER met2 ;
        RECT 5.320 13.440 5.880 13.720 ;
      LAYER met2 ;
        RECT 5.040 13.160 5.600 13.440 ;
      LAYER met2 ;
        RECT 4.760 12.880 5.320 13.160 ;
      LAYER met2 ;
        RECT 5.320 12.880 5.600 13.160 ;
      LAYER met2 ;
        RECT 5.600 12.880 5.880 13.440 ;
      LAYER met2 ;
        RECT 5.880 12.880 6.160 13.720 ;
      LAYER met2 ;
        RECT 6.160 13.440 7.840 14.000 ;
      LAYER met2 ;
        RECT 7.840 13.720 8.400 14.560 ;
      LAYER met2 ;
        RECT 8.400 13.720 8.960 14.560 ;
      LAYER met2 ;
        RECT 8.960 13.720 9.520 14.560 ;
      LAYER met2 ;
        RECT 9.520 14.280 10.080 14.560 ;
      LAYER met2 ;
        RECT 10.080 14.280 10.640 14.560 ;
      LAYER met2 ;
        RECT 10.640 14.280 11.760 14.840 ;
        RECT 9.520 13.720 11.760 14.280 ;
      LAYER met2 ;
        RECT 7.840 13.440 8.120 13.720 ;
      LAYER met2 ;
        RECT 8.120 13.440 8.960 13.720 ;
      LAYER met2 ;
        RECT 8.960 13.440 10.360 13.720 ;
      LAYER met2 ;
        RECT 10.360 13.440 11.760 13.720 ;
        RECT 6.160 13.160 7.560 13.440 ;
      LAYER met2 ;
        RECT 7.560 13.160 8.120 13.440 ;
      LAYER met2 ;
        RECT 8.120 13.160 10.080 13.440 ;
      LAYER met2 ;
        RECT 4.480 12.600 5.040 12.880 ;
      LAYER met2 ;
        RECT 5.040 12.600 5.320 12.880 ;
      LAYER met2 ;
        RECT 5.320 12.600 6.160 12.880 ;
      LAYER met2 ;
        RECT 6.160 12.600 7.280 13.160 ;
      LAYER met2 ;
        RECT 7.280 12.600 7.840 13.160 ;
      LAYER met2 ;
        RECT 7.840 12.600 10.080 13.160 ;
        RECT 0.000 12.040 2.520 12.600 ;
      LAYER met2 ;
        RECT 2.520 12.320 3.080 12.600 ;
      LAYER met2 ;
        RECT 3.080 12.320 4.760 12.600 ;
      LAYER met2 ;
        RECT 4.760 12.320 5.040 12.600 ;
      LAYER met2 ;
        RECT 5.040 12.320 5.600 12.600 ;
      LAYER met2 ;
        RECT 5.600 12.320 5.880 12.600 ;
        RECT 2.520 12.040 3.640 12.320 ;
      LAYER met2 ;
        RECT 3.640 12.040 4.760 12.320 ;
      LAYER met2 ;
        RECT 4.760 12.040 5.880 12.320 ;
      LAYER met2 ;
        RECT 5.880 12.040 7.000 12.600 ;
      LAYER met2 ;
        RECT 7.000 12.320 7.560 12.600 ;
      LAYER met2 ;
        RECT 7.560 12.320 8.960 12.600 ;
      LAYER met2 ;
        RECT 8.960 12.320 9.520 12.600 ;
      LAYER met2 ;
        RECT 9.520 12.320 10.080 12.600 ;
      LAYER met2 ;
        RECT 10.080 12.320 10.640 13.440 ;
      LAYER met2 ;
        RECT 10.640 12.320 11.760 13.440 ;
      LAYER met2 ;
        RECT 7.000 12.040 8.120 12.320 ;
      LAYER met2 ;
        RECT 8.120 12.040 8.960 12.320 ;
      LAYER met2 ;
        RECT 8.960 12.040 10.360 12.320 ;
      LAYER met2 ;
        RECT 0.000 11.760 2.240 12.040 ;
      LAYER met2 ;
        RECT 2.240 11.760 3.920 12.040 ;
      LAYER met2 ;
        RECT 3.920 11.760 5.040 12.040 ;
      LAYER met2 ;
        RECT 5.040 11.760 5.600 12.040 ;
      LAYER met2 ;
        RECT 5.600 11.760 6.720 12.040 ;
      LAYER met2 ;
        RECT 6.720 11.760 8.400 12.040 ;
      LAYER met2 ;
        RECT 8.400 11.760 9.240 12.040 ;
      LAYER met2 ;
        RECT 9.240 11.760 10.360 12.040 ;
      LAYER met2 ;
        RECT 10.360 11.760 11.760 12.320 ;
        RECT 0.000 11.200 11.760 11.760 ;
        RECT 0.000 10.080 1.120 11.200 ;
      LAYER met2 ;
        RECT 1.120 10.080 3.640 11.200 ;
      LAYER met2 ;
        RECT 3.640 10.080 11.760 11.200 ;
        RECT 0.000 7.280 1.680 10.080 ;
        RECT 0.000 7.000 0.280 7.280 ;
      LAYER met2 ;
        RECT 0.280 7.000 1.120 7.280 ;
      LAYER met2 ;
        RECT 1.120 7.000 1.680 7.280 ;
      LAYER met2 ;
        RECT 0.000 6.160 1.400 7.000 ;
      LAYER met2 ;
        RECT 1.400 6.160 1.680 7.000 ;
      LAYER met2 ;
        RECT 1.680 6.160 3.080 10.080 ;
      LAYER met2 ;
        RECT 3.080 9.240 4.200 10.080 ;
      LAYER met2 ;
        RECT 4.200 9.240 7.280 10.080 ;
      LAYER met2 ;
        RECT 7.280 9.240 11.760 10.080 ;
        RECT 3.080 7.560 3.640 9.240 ;
      LAYER met2 ;
        RECT 3.640 8.960 7.560 9.240 ;
        RECT 3.640 7.560 5.040 8.960 ;
      LAYER met2 ;
        RECT 5.040 8.400 6.160 8.960 ;
      LAYER met2 ;
        RECT 6.160 8.400 7.560 8.960 ;
      LAYER met2 ;
        RECT 5.040 8.120 6.440 8.400 ;
      LAYER met2 ;
        RECT 6.440 8.120 7.560 8.400 ;
      LAYER met2 ;
        RECT 7.560 8.120 8.120 9.240 ;
        RECT 5.040 7.560 8.120 8.120 ;
        RECT 3.080 7.280 3.920 7.560 ;
      LAYER met2 ;
        RECT 3.920 7.280 7.280 7.560 ;
      LAYER met2 ;
        RECT 3.080 6.440 4.200 7.280 ;
      LAYER met2 ;
        RECT 4.200 6.720 7.280 7.280 ;
      LAYER met2 ;
        RECT 7.280 6.720 8.120 7.560 ;
      LAYER met2 ;
        RECT 8.120 6.720 9.520 9.240 ;
      LAYER met2 ;
        RECT 9.520 8.400 10.640 9.240 ;
      LAYER met2 ;
        RECT 10.640 8.400 11.760 9.240 ;
      LAYER met2 ;
        RECT 9.520 7.560 10.360 8.400 ;
      LAYER met2 ;
        RECT 10.360 7.560 11.760 8.400 ;
      LAYER met2 ;
        RECT 9.520 6.720 9.800 7.560 ;
      LAYER met2 ;
        RECT 9.800 7.280 11.760 7.560 ;
        RECT 9.800 6.720 11.200 7.280 ;
        RECT 4.200 6.440 7.560 6.720 ;
      LAYER met2 ;
        RECT 3.080 6.160 6.160 6.440 ;
        RECT 0.000 5.880 0.280 6.160 ;
      LAYER met2 ;
        RECT 0.280 5.880 3.080 6.160 ;
      LAYER met2 ;
        RECT 3.080 5.880 3.920 6.160 ;
      LAYER met2 ;
        RECT 3.920 5.880 4.760 6.160 ;
      LAYER met2 ;
        RECT 4.760 5.880 6.160 6.160 ;
        RECT 0.000 5.040 0.560 5.880 ;
      LAYER met2 ;
        RECT 0.560 5.320 2.800 5.880 ;
      LAYER met2 ;
        RECT 2.800 5.320 3.640 5.880 ;
      LAYER met2 ;
        RECT 0.560 5.040 2.520 5.320 ;
      LAYER met2 ;
        RECT 2.520 5.040 3.640 5.320 ;
      LAYER met2 ;
        RECT 3.640 5.040 5.040 5.880 ;
      LAYER met2 ;
        RECT 5.040 5.040 6.160 5.880 ;
      LAYER met2 ;
        RECT 6.160 5.040 7.560 6.440 ;
      LAYER met2 ;
        RECT 0.000 4.760 3.920 5.040 ;
      LAYER met2 ;
        RECT 3.920 4.760 7.560 5.040 ;
      LAYER met2 ;
        RECT 7.560 4.760 8.120 6.720 ;
      LAYER met2 ;
        RECT 8.120 6.440 11.200 6.720 ;
      LAYER met2 ;
        RECT 11.200 6.440 11.760 7.280 ;
      LAYER met2 ;
        RECT 8.120 5.880 10.640 6.440 ;
      LAYER met2 ;
        RECT 10.640 5.880 11.760 6.440 ;
      LAYER met2 ;
        RECT 8.120 5.600 11.200 5.880 ;
      LAYER met2 ;
        RECT 0.000 3.920 4.200 4.760 ;
      LAYER met2 ;
        RECT 4.200 4.200 7.280 4.760 ;
      LAYER met2 ;
        RECT 7.280 4.200 8.120 4.760 ;
      LAYER met2 ;
        RECT 4.200 3.920 7.000 4.200 ;
      LAYER met2 ;
        RECT 7.000 3.920 8.120 4.200 ;
        RECT 0.000 3.360 8.120 3.920 ;
      LAYER met2 ;
        RECT 8.120 3.360 9.520 5.600 ;
      LAYER met2 ;
        RECT 9.520 4.760 9.800 5.600 ;
      LAYER met2 ;
        RECT 9.800 5.040 11.200 5.600 ;
      LAYER met2 ;
        RECT 11.200 5.040 11.760 5.880 ;
      LAYER met2 ;
        RECT 9.800 4.760 11.760 5.040 ;
      LAYER met2 ;
        RECT 9.520 3.920 10.360 4.760 ;
      LAYER met2 ;
        RECT 10.360 3.920 11.760 4.760 ;
      LAYER met2 ;
        RECT 9.520 3.360 10.640 3.920 ;
      LAYER met2 ;
        RECT 10.640 3.360 11.760 3.920 ;
      LAYER met2 ;
        RECT 0.000 3.080 8.400 3.360 ;
      LAYER met2 ;
        RECT 8.400 3.080 9.520 3.360 ;
      LAYER met2 ;
        RECT 9.520 3.080 10.920 3.360 ;
      LAYER met2 ;
        RECT 10.920 3.080 11.760 3.360 ;
      LAYER met2 ;
        RECT 0.000 2.800 11.760 3.080 ;
        RECT 0.000 2.240 2.240 2.800 ;
      LAYER met2 ;
        RECT 2.240 2.240 5.880 2.800 ;
      LAYER met2 ;
        RECT 5.880 2.520 6.720 2.800 ;
      LAYER met2 ;
        RECT 6.720 2.520 7.280 2.800 ;
      LAYER met2 ;
        RECT 7.280 2.520 8.680 2.800 ;
      LAYER met2 ;
        RECT 8.680 2.520 9.240 2.800 ;
      LAYER met2 ;
        RECT 9.240 2.520 11.760 2.800 ;
        RECT 5.880 2.240 6.440 2.520 ;
        RECT 0.000 0.000 2.800 2.240 ;
      LAYER met2 ;
        RECT 2.800 0.000 3.360 2.240 ;
      LAYER met2 ;
        RECT 3.360 0.000 4.760 2.240 ;
      LAYER met2 ;
        RECT 4.760 0.000 5.320 2.240 ;
      LAYER met2 ;
        RECT 5.320 1.960 6.440 2.240 ;
      LAYER met2 ;
        RECT 6.440 1.960 7.280 2.520 ;
      LAYER met2 ;
        RECT 7.280 1.960 8.400 2.520 ;
      LAYER met2 ;
        RECT 8.400 2.240 9.520 2.520 ;
        RECT 8.400 1.960 8.680 2.240 ;
      LAYER met2 ;
        RECT 8.680 1.960 9.240 2.240 ;
      LAYER met2 ;
        RECT 9.240 1.960 9.520 2.240 ;
      LAYER met2 ;
        RECT 9.520 1.960 11.760 2.520 ;
        RECT 5.320 0.280 6.720 1.960 ;
      LAYER met2 ;
        RECT 6.720 0.280 7.280 1.960 ;
      LAYER met2 ;
        RECT 7.280 0.560 8.120 1.960 ;
      LAYER met2 ;
        RECT 8.120 1.680 8.960 1.960 ;
      LAYER met2 ;
        RECT 8.960 1.680 9.240 1.960 ;
      LAYER met2 ;
        RECT 9.240 1.680 9.800 1.960 ;
        RECT 8.120 0.840 8.400 1.680 ;
      LAYER met2 ;
        RECT 8.400 1.120 8.680 1.680 ;
      LAYER met2 ;
        RECT 8.680 1.400 8.960 1.680 ;
      LAYER met2 ;
        RECT 8.960 1.400 9.520 1.680 ;
      LAYER met2 ;
        RECT 8.680 1.120 9.240 1.400 ;
      LAYER met2 ;
        RECT 8.400 0.840 8.960 1.120 ;
      LAYER met2 ;
        RECT 8.960 0.840 9.240 1.120 ;
      LAYER met2 ;
        RECT 9.240 0.840 9.520 1.400 ;
      LAYER met2 ;
        RECT 9.520 0.840 9.800 1.680 ;
        RECT 8.120 0.560 8.680 0.840 ;
      LAYER met2 ;
        RECT 8.680 0.560 8.960 0.840 ;
      LAYER met2 ;
        RECT 8.960 0.560 9.800 0.840 ;
      LAYER met2 ;
        RECT 9.800 0.560 11.760 1.960 ;
        RECT 7.280 0.280 8.400 0.560 ;
      LAYER met2 ;
        RECT 8.400 0.280 8.680 0.560 ;
      LAYER met2 ;
        RECT 8.680 0.280 9.240 0.560 ;
      LAYER met2 ;
        RECT 9.240 0.280 9.520 0.560 ;
      LAYER met2 ;
        RECT 5.320 0.000 6.160 0.280 ;
      LAYER met2 ;
        RECT 6.160 0.000 7.840 0.280 ;
      LAYER met2 ;
        RECT 7.840 0.000 8.400 0.280 ;
      LAYER met2 ;
        RECT 8.400 0.000 9.520 0.280 ;
      LAYER met2 ;
        RECT 9.520 0.000 11.760 0.560 ;
      LAYER met3 ;
        RECT 0.000 0.000 11.760 15.120 ;
      LAYER met4 ;
        RECT 0.000 0.000 11.760 15.120 ;
      LAYER met5 ;
        RECT 0.000 0.000 11.760 15.120 ;
  END
END jsk
END LIBRARY

