magic
tech sky130A
magscale 1 2
timestamp 1738298459
<< viali >>
rect 6469 21641 6503 21675
rect 7297 21641 7331 21675
rect 8401 21641 8435 21675
rect 8677 21641 8711 21675
rect 9413 21641 9447 21675
rect 10333 21641 10367 21675
rect 11805 21641 11839 21675
rect 12265 21641 12299 21675
rect 12817 21641 12851 21675
rect 25697 21573 25731 21607
rect 3525 21505 3559 21539
rect 11161 21505 11195 21539
rect 29009 21505 29043 21539
rect 2789 21437 2823 21471
rect 3065 21437 3099 21471
rect 3249 21437 3283 21471
rect 3341 21437 3375 21471
rect 3985 21437 4019 21471
rect 4077 21437 4111 21471
rect 4261 21437 4295 21471
rect 6101 21437 6135 21471
rect 6653 21437 6687 21471
rect 8217 21437 8251 21471
rect 9229 21437 9263 21471
rect 9597 21437 9631 21471
rect 9689 21437 9723 21471
rect 9873 21437 9907 21471
rect 9965 21437 9999 21471
rect 10517 21437 10551 21471
rect 11253 21437 11287 21471
rect 11345 21437 11379 21471
rect 11529 21437 11563 21471
rect 15669 21437 15703 21471
rect 16405 21437 16439 21471
rect 16681 21437 16715 21471
rect 16957 21437 16991 21471
rect 19165 21437 19199 21471
rect 19533 21437 19567 21471
rect 19809 21437 19843 21471
rect 21649 21437 21683 21471
rect 23857 21437 23891 21471
rect 24409 21437 24443 21471
rect 24961 21437 24995 21471
rect 25513 21437 25547 21471
rect 25789 21437 25823 21471
rect 26065 21437 26099 21471
rect 27905 21437 27939 21471
rect 27997 21437 28031 21471
rect 28273 21437 28307 21471
rect 29285 21437 29319 21471
rect 2973 21369 3007 21403
rect 3893 21369 3927 21403
rect 6929 21369 6963 21403
rect 7113 21369 7147 21403
rect 7573 21369 7607 21403
rect 16865 21369 16899 21403
rect 19257 21369 19291 21403
rect 19349 21369 19383 21403
rect 27638 21369 27672 21403
rect 2697 21301 2731 21335
rect 3525 21301 3559 21335
rect 4077 21301 4111 21335
rect 6193 21301 6227 21335
rect 6745 21301 6779 21335
rect 10149 21301 10183 21335
rect 11621 21301 11655 21335
rect 15577 21301 15611 21335
rect 16497 21301 16531 21335
rect 17049 21301 17083 21335
rect 18981 21301 19015 21335
rect 19717 21301 19751 21335
rect 21833 21301 21867 21335
rect 24041 21301 24075 21335
rect 24593 21301 24627 21335
rect 25145 21301 25179 21335
rect 25973 21301 26007 21335
rect 26249 21301 26283 21335
rect 26525 21301 26559 21335
rect 28181 21301 28215 21335
rect 28457 21301 28491 21335
rect 1041 21097 1075 21131
rect 4261 21097 4295 21131
rect 6285 21097 6319 21131
rect 7941 21097 7975 21131
rect 8493 21097 8527 21131
rect 10149 21097 10183 21131
rect 12633 21097 12667 21131
rect 16405 21097 16439 21131
rect 20085 21097 20119 21131
rect 11713 21029 11747 21063
rect 18153 21029 18187 21063
rect 23888 21029 23922 21063
rect 27546 21029 27580 21063
rect 29018 21029 29052 21063
rect 2165 20961 2199 20995
rect 2421 20961 2455 20995
rect 2513 20961 2547 20995
rect 2789 20961 2823 20995
rect 4169 20961 4203 20995
rect 4445 20961 4479 20995
rect 4629 20961 4663 20995
rect 5549 20961 5583 20995
rect 6101 20961 6135 20995
rect 6469 20961 6503 20995
rect 6561 20961 6595 20995
rect 6828 20961 6862 20995
rect 8309 20961 8343 20995
rect 8861 20961 8895 20995
rect 9137 20961 9171 20995
rect 9321 20961 9355 20995
rect 9413 20961 9447 20995
rect 10057 20961 10091 20995
rect 11253 20961 11287 20995
rect 12081 20961 12115 20995
rect 12357 20961 12391 20995
rect 12817 20961 12851 20995
rect 13829 20961 13863 20995
rect 15209 20961 15243 20995
rect 15301 20961 15335 20995
rect 15485 20961 15519 20995
rect 15761 20961 15795 20995
rect 15945 20961 15979 20995
rect 17785 20961 17819 20995
rect 18015 20961 18049 20995
rect 18245 20961 18279 20995
rect 18373 20961 18407 20995
rect 18521 20961 18555 20995
rect 18705 20961 18739 20995
rect 22394 20961 22428 20995
rect 22661 20961 22695 20995
rect 24133 20961 24167 20995
rect 25338 20961 25372 20995
rect 30490 20961 30524 20995
rect 30757 20961 30791 20995
rect 10701 20893 10735 20927
rect 17509 20893 17543 20927
rect 18981 20893 19015 20927
rect 25605 20893 25639 20927
rect 27813 20893 27847 20927
rect 29285 20893 29319 20927
rect 11529 20825 11563 20859
rect 13001 20825 13035 20859
rect 5457 20757 5491 20791
rect 5917 20757 5951 20791
rect 8677 20757 8711 20791
rect 13737 20757 13771 20791
rect 15669 20757 15703 20791
rect 15853 20757 15887 20791
rect 17877 20757 17911 20791
rect 21281 20757 21315 20791
rect 22753 20757 22787 20791
rect 24225 20757 24259 20791
rect 26433 20757 26467 20791
rect 27905 20757 27939 20791
rect 29377 20757 29411 20791
rect 2605 20553 2639 20587
rect 4353 20553 4387 20587
rect 8585 20553 8619 20587
rect 10333 20553 10367 20587
rect 11989 20553 12023 20587
rect 16957 20553 16991 20587
rect 17141 20553 17175 20587
rect 20269 20553 20303 20587
rect 17877 20485 17911 20519
rect 5273 20417 5307 20451
rect 6653 20417 6687 20451
rect 13553 20417 13587 20451
rect 15393 20417 15427 20451
rect 18705 20417 18739 20451
rect 20453 20417 20487 20451
rect 29101 20417 29135 20451
rect 29561 20417 29595 20451
rect 2237 20349 2271 20383
rect 2789 20349 2823 20383
rect 3065 20349 3099 20383
rect 4077 20349 4111 20383
rect 4537 20349 4571 20383
rect 4629 20349 4663 20383
rect 4721 20349 4755 20383
rect 4997 20349 5031 20383
rect 5181 20349 5215 20383
rect 5549 20349 5583 20383
rect 8033 20349 8067 20383
rect 8401 20349 8435 20383
rect 8953 20349 8987 20383
rect 9220 20349 9254 20383
rect 10609 20349 10643 20383
rect 12173 20349 12207 20383
rect 12265 20349 12299 20383
rect 13185 20349 13219 20383
rect 13829 20349 13863 20383
rect 15669 20349 15703 20383
rect 17417 20349 17451 20383
rect 17509 20349 17543 20383
rect 17601 20349 17635 20383
rect 17785 20349 17819 20383
rect 18153 20349 18187 20383
rect 18245 20349 18279 20383
rect 18337 20349 18371 20383
rect 18521 20349 18555 20383
rect 18981 20349 19015 20383
rect 20637 20349 20671 20383
rect 20913 20349 20947 20383
rect 21925 20349 21959 20383
rect 22293 20349 22327 20383
rect 22569 20349 22603 20383
rect 22661 20349 22695 20383
rect 22845 20349 22879 20383
rect 22937 20349 22971 20383
rect 25522 20349 25556 20383
rect 25789 20349 25823 20383
rect 27261 20349 27295 20383
rect 29009 20349 29043 20383
rect 29285 20349 29319 20383
rect 2973 20281 3007 20315
rect 4353 20281 4387 20315
rect 10876 20281 10910 20315
rect 20821 20281 20855 20315
rect 22109 20281 22143 20315
rect 22201 20281 22235 20315
rect 26994 20281 27028 20315
rect 29806 20281 29840 20315
rect 2145 20213 2179 20247
rect 3433 20213 3467 20247
rect 4813 20213 4847 20247
rect 8125 20213 8159 20247
rect 13277 20213 13311 20247
rect 15117 20213 15151 20247
rect 22477 20213 22511 20247
rect 23121 20213 23155 20247
rect 24409 20213 24443 20247
rect 25881 20213 25915 20247
rect 29377 20213 29411 20247
rect 30941 20213 30975 20247
rect 5273 20009 5307 20043
rect 7573 20009 7607 20043
rect 8493 20009 8527 20043
rect 10149 20009 10183 20043
rect 11069 20009 11103 20043
rect 14933 20009 14967 20043
rect 17233 20009 17267 20043
rect 18245 20009 18279 20043
rect 18705 20009 18739 20043
rect 19809 20009 19843 20043
rect 29469 20009 29503 20043
rect 2228 19941 2262 19975
rect 5825 19941 5859 19975
rect 9036 19941 9070 19975
rect 15577 19941 15611 19975
rect 16497 19941 16531 19975
rect 17601 19941 17635 19975
rect 23857 19941 23891 19975
rect 27905 19941 27939 19975
rect 1961 19873 1995 19907
rect 3433 19873 3467 19907
rect 3689 19873 3723 19907
rect 5273 19873 5307 19907
rect 5457 19873 5491 19907
rect 6009 19873 6043 19907
rect 6193 19873 6227 19907
rect 6285 19873 6319 19907
rect 7389 19873 7423 19907
rect 8401 19873 8435 19907
rect 8769 19873 8803 19907
rect 11345 19873 11379 19907
rect 11437 19873 11471 19907
rect 11529 19873 11563 19907
rect 11713 19873 11747 19907
rect 13369 19873 13403 19907
rect 15393 19873 15427 19907
rect 15485 19873 15519 19907
rect 15761 19873 15795 19907
rect 16129 19873 16163 19907
rect 16277 19873 16311 19907
rect 16405 19873 16439 19907
rect 16635 19873 16669 19907
rect 17049 19873 17083 19907
rect 17325 19873 17359 19907
rect 18153 19873 18187 19907
rect 18429 19873 18463 19907
rect 18613 19873 18647 19907
rect 18981 19873 19015 19907
rect 19073 19873 19107 19907
rect 19165 19873 19199 19907
rect 19349 19873 19383 19907
rect 19625 19873 19659 19907
rect 19901 19873 19935 19907
rect 21557 19873 21591 19907
rect 22293 19873 22327 19907
rect 22385 19873 22419 19907
rect 22496 19873 22530 19907
rect 22661 19879 22695 19913
rect 23121 19873 23155 19907
rect 23213 19873 23247 19907
rect 23397 19873 23431 19907
rect 23489 19873 23523 19907
rect 23765 19873 23799 19907
rect 23949 19873 23983 19907
rect 24133 19873 24167 19907
rect 27721 19873 27755 19907
rect 28825 19873 28859 19907
rect 29009 19873 29043 19907
rect 29101 19873 29135 19907
rect 29193 19873 29227 19907
rect 29561 19873 29595 19907
rect 29828 19873 29862 19907
rect 6377 19805 6411 19839
rect 7113 19805 7147 19839
rect 7205 19805 7239 19839
rect 7297 19805 7331 19839
rect 13645 19805 13679 19839
rect 17417 19805 17451 19839
rect 19441 19805 19475 19839
rect 22937 19805 22971 19839
rect 25697 19805 25731 19839
rect 15945 19737 15979 19771
rect 16773 19737 16807 19771
rect 18521 19737 18555 19771
rect 3341 19669 3375 19703
rect 4813 19669 4847 19703
rect 15209 19669 15243 19703
rect 16865 19669 16899 19703
rect 21465 19669 21499 19703
rect 22845 19669 22879 19703
rect 23581 19669 23615 19703
rect 25145 19669 25179 19703
rect 27629 19669 27663 19703
rect 27997 19669 28031 19703
rect 30941 19669 30975 19703
rect 2421 19465 2455 19499
rect 6469 19465 6503 19499
rect 9045 19465 9079 19499
rect 16129 19465 16163 19499
rect 16313 19465 16347 19499
rect 16589 19465 16623 19499
rect 16773 19465 16807 19499
rect 17601 19465 17635 19499
rect 17693 19465 17727 19499
rect 19073 19465 19107 19499
rect 29745 19465 29779 19499
rect 22017 19397 22051 19431
rect 3985 19329 4019 19363
rect 15025 19329 15059 19363
rect 17693 19329 17727 19363
rect 22293 19329 22327 19363
rect 25881 19329 25915 19363
rect 1961 19261 1995 19295
rect 2053 19261 2087 19295
rect 2145 19261 2179 19295
rect 2329 19261 2363 19295
rect 2697 19261 2731 19295
rect 2789 19261 2823 19295
rect 2881 19261 2915 19295
rect 3065 19261 3099 19295
rect 3433 19261 3467 19295
rect 4169 19261 4203 19295
rect 5825 19261 5859 19295
rect 5973 19261 6007 19295
rect 6331 19261 6365 19295
rect 6561 19261 6595 19295
rect 6753 19271 6787 19305
rect 9045 19261 9079 19295
rect 9229 19261 9263 19295
rect 11161 19261 11195 19295
rect 14565 19261 14599 19295
rect 14749 19261 14783 19295
rect 14933 19261 14967 19295
rect 15117 19261 15151 19295
rect 15301 19261 15335 19295
rect 15669 19261 15703 19295
rect 15761 19261 15795 19295
rect 15853 19261 15887 19295
rect 16037 19261 16071 19295
rect 16865 19261 16899 19295
rect 17141 19261 17175 19295
rect 17233 19261 17267 19295
rect 17427 19261 17461 19295
rect 17555 19261 17589 19295
rect 17877 19261 17911 19295
rect 18981 19261 19015 19295
rect 19165 19261 19199 19295
rect 21833 19261 21867 19295
rect 22477 19261 22511 19295
rect 22569 19261 22603 19295
rect 22753 19261 22787 19295
rect 22845 19261 22879 19295
rect 24409 19261 24443 19295
rect 25329 19261 25363 19295
rect 25488 19261 25522 19295
rect 25605 19261 25639 19295
rect 26341 19261 26375 19295
rect 26525 19261 26559 19295
rect 26709 19261 26743 19295
rect 26893 19261 26927 19295
rect 26985 19261 27019 19295
rect 27077 19261 27111 19295
rect 27445 19261 27479 19295
rect 29101 19261 29135 19295
rect 29285 19261 29319 19295
rect 29377 19261 29411 19295
rect 29469 19261 29503 19295
rect 30021 19261 30055 19295
rect 30113 19261 30147 19295
rect 30297 19261 30331 19295
rect 30389 19261 30423 19295
rect 30481 19261 30515 19295
rect 3249 19193 3283 19227
rect 3617 19193 3651 19227
rect 6101 19193 6135 19227
rect 6193 19193 6227 19227
rect 6653 19193 6687 19227
rect 15393 19193 15427 19227
rect 16297 19193 16331 19227
rect 16497 19193 16531 19227
rect 21097 19193 21131 19227
rect 21649 19193 21683 19227
rect 23121 19193 23155 19227
rect 27353 19193 27387 19227
rect 27690 19193 27724 19227
rect 1685 19125 1719 19159
rect 4077 19125 4111 19159
rect 4537 19125 4571 19159
rect 11253 19125 11287 19159
rect 17233 19125 17267 19159
rect 21005 19125 21039 19159
rect 21373 19125 21407 19159
rect 23029 19125 23063 19159
rect 24501 19125 24535 19159
rect 24685 19125 24719 19159
rect 28825 19125 28859 19159
rect 29837 19125 29871 19159
rect 30665 19125 30699 19159
rect 2329 18921 2363 18955
rect 5089 18921 5123 18955
rect 6469 18921 6503 18955
rect 7205 18921 7239 18955
rect 11253 18921 11287 18955
rect 14473 18921 14507 18955
rect 16497 18921 16531 18955
rect 17509 18921 17543 18955
rect 22661 18921 22695 18955
rect 25973 18921 26007 18955
rect 26709 18921 26743 18955
rect 27261 18921 27295 18955
rect 29377 18921 29411 18955
rect 29469 18921 29503 18955
rect 29837 18921 29871 18955
rect 29929 18921 29963 18955
rect 6377 18853 6411 18887
rect 11437 18853 11471 18887
rect 21548 18853 21582 18887
rect 24501 18853 24535 18887
rect 24838 18853 24872 18887
rect 29009 18853 29043 18887
rect 1961 18785 1995 18819
rect 2145 18785 2179 18819
rect 2421 18785 2455 18819
rect 2605 18785 2639 18819
rect 2697 18785 2731 18819
rect 2789 18785 2823 18819
rect 4261 18785 4295 18819
rect 4997 18785 5031 18819
rect 5181 18785 5215 18819
rect 6193 18785 6227 18819
rect 6469 18785 6503 18819
rect 7389 18785 7423 18819
rect 7573 18785 7607 18819
rect 11621 18785 11655 18819
rect 11897 18785 11931 18819
rect 14749 18785 14783 18819
rect 14841 18785 14875 18819
rect 14933 18785 14967 18819
rect 15117 18785 15151 18819
rect 15393 18785 15427 18819
rect 15485 18785 15519 18819
rect 15669 18785 15703 18819
rect 15761 18785 15795 18819
rect 16129 18785 16163 18819
rect 16313 18785 16347 18819
rect 16589 18785 16623 18819
rect 16681 18785 16715 18819
rect 16865 18785 16899 18819
rect 16957 18785 16991 18819
rect 17141 18785 17175 18819
rect 17233 18785 17267 18819
rect 17325 18785 17359 18819
rect 20085 18785 20119 18819
rect 20269 18785 20303 18819
rect 20453 18785 20487 18819
rect 20637 18785 20671 18819
rect 20729 18785 20763 18819
rect 20821 18785 20855 18819
rect 21281 18785 21315 18819
rect 22937 18785 22971 18819
rect 23857 18785 23891 18819
rect 24041 18785 24075 18819
rect 24133 18785 24167 18819
rect 24225 18785 24259 18819
rect 24593 18785 24627 18819
rect 26801 18785 26835 18819
rect 27445 18785 27479 18819
rect 27537 18785 27571 18819
rect 27721 18785 27755 18819
rect 27813 18785 27847 18819
rect 28365 18785 28399 18819
rect 28549 18785 28583 18819
rect 28641 18785 28675 18819
rect 28733 18785 28767 18819
rect 30113 18785 30147 18819
rect 30205 18785 30239 18819
rect 30389 18785 30423 18819
rect 30481 18785 30515 18819
rect 3801 18717 3835 18751
rect 3985 18717 4019 18751
rect 4169 18717 4203 18751
rect 15209 18717 15243 18751
rect 26525 18717 26559 18751
rect 29193 18717 29227 18751
rect 3157 18649 3191 18683
rect 4629 18649 4663 18683
rect 11713 18649 11747 18683
rect 27169 18649 27203 18683
rect 3065 18581 3099 18615
rect 16773 18581 16807 18615
rect 20177 18581 20211 18615
rect 21097 18581 21131 18615
rect 22845 18581 22879 18615
rect 1501 18377 1535 18411
rect 10977 18377 11011 18411
rect 15301 18377 15335 18411
rect 20545 18377 20579 18411
rect 24133 18377 24167 18411
rect 26985 18377 27019 18411
rect 28089 18377 28123 18411
rect 28825 18377 28859 18411
rect 30205 18377 30239 18411
rect 6929 18309 6963 18343
rect 16589 18309 16623 18343
rect 17785 18309 17819 18343
rect 10149 18241 10183 18275
rect 16313 18241 16347 18275
rect 16681 18241 16715 18275
rect 17049 18241 17083 18275
rect 17417 18241 17451 18275
rect 17509 18241 17543 18275
rect 21005 18241 21039 18275
rect 21097 18241 21131 18275
rect 21189 18241 21223 18275
rect 25329 18241 25363 18275
rect 29377 18241 29411 18275
rect 29561 18241 29595 18275
rect 29745 18241 29779 18275
rect 1409 18173 1443 18207
rect 2973 18173 3007 18207
rect 4629 18173 4663 18207
rect 7205 18173 7239 18207
rect 7757 18173 7791 18207
rect 7849 18173 7883 18207
rect 7941 18173 7975 18207
rect 8125 18173 8159 18207
rect 9413 18173 9447 18207
rect 10057 18173 10091 18207
rect 10517 18173 10551 18207
rect 10701 18173 10735 18207
rect 12357 18173 12391 18207
rect 12541 18173 12575 18207
rect 12633 18173 12667 18207
rect 13645 18173 13679 18207
rect 13737 18173 13771 18207
rect 13921 18173 13955 18207
rect 14197 18173 14231 18207
rect 15853 18173 15887 18207
rect 15945 18173 15979 18207
rect 16129 18173 16163 18207
rect 16221 18173 16255 18207
rect 16497 18173 16531 18207
rect 16773 18173 16807 18207
rect 16957 18173 16991 18207
rect 17233 18173 17267 18207
rect 17325 18173 17359 18207
rect 17693 18173 17727 18207
rect 17877 18183 17911 18217
rect 19901 18173 19935 18207
rect 20085 18173 20119 18207
rect 20453 18173 20487 18207
rect 20637 18173 20671 18207
rect 20913 18173 20947 18207
rect 23489 18173 23523 18207
rect 24317 18173 24351 18207
rect 24409 18173 24443 18207
rect 24593 18173 24627 18207
rect 24685 18173 24719 18207
rect 25881 18173 25915 18207
rect 26065 18173 26099 18207
rect 26249 18173 26283 18207
rect 26341 18173 26375 18207
rect 26525 18173 26559 18207
rect 26617 18173 26651 18207
rect 26709 18173 26743 18207
rect 28181 18173 28215 18207
rect 28365 18173 28399 18207
rect 28457 18173 28491 18207
rect 28549 18173 28583 18207
rect 29837 18173 29871 18207
rect 1685 18105 1719 18139
rect 1869 18105 1903 18139
rect 1961 18105 1995 18139
rect 2145 18105 2179 18139
rect 2329 18105 2363 18139
rect 4362 18105 4396 18139
rect 6561 18105 6595 18139
rect 12090 18105 12124 18139
rect 15669 18105 15703 18139
rect 19349 18105 19383 18139
rect 19533 18105 19567 18139
rect 23305 18105 23339 18139
rect 27721 18105 27755 18139
rect 27905 18105 27939 18139
rect 29009 18105 29043 18139
rect 29193 18105 29227 18139
rect 1317 18037 1351 18071
rect 2421 18037 2455 18071
rect 3249 18037 3283 18071
rect 7021 18037 7055 18071
rect 7297 18037 7331 18071
rect 7481 18037 7515 18071
rect 19441 18037 19475 18071
rect 21373 18037 21407 18071
rect 23673 18037 23707 18071
rect 24777 18037 24811 18071
rect 25145 18037 25179 18071
rect 25237 18037 25271 18071
rect 3341 17833 3375 17867
rect 4261 17833 4295 17867
rect 9505 17833 9539 17867
rect 10149 17833 10183 17867
rect 10701 17833 10735 17867
rect 11621 17833 11655 17867
rect 13277 17833 13311 17867
rect 14657 17833 14691 17867
rect 16129 17833 16163 17867
rect 25237 17833 25271 17867
rect 29377 17833 29411 17867
rect 5825 17765 5859 17799
rect 1961 17697 1995 17731
rect 2228 17697 2262 17731
rect 3617 17697 3651 17731
rect 3801 17697 3835 17731
rect 3893 17697 3927 17731
rect 4169 17697 4203 17731
rect 6009 17697 6043 17731
rect 6101 17697 6135 17731
rect 6469 17697 6503 17731
rect 6653 17697 6687 17731
rect 6745 17697 6779 17731
rect 6837 17697 6871 17731
rect 7297 17697 7331 17731
rect 7564 17697 7598 17731
rect 9873 17697 9907 17731
rect 10241 17697 10275 17731
rect 10333 17697 10367 17731
rect 10517 17697 10551 17731
rect 10977 17697 11011 17731
rect 11161 17697 11195 17731
rect 11253 17697 11287 17731
rect 11345 17697 11379 17731
rect 12081 17697 12115 17731
rect 12357 17697 12391 17731
rect 12541 17697 12575 17731
rect 13553 17697 13587 17731
rect 13829 17697 13863 17731
rect 14933 17697 14967 17731
rect 15025 17697 15059 17731
rect 15117 17697 15151 17731
rect 15301 17697 15335 17731
rect 15761 17697 15795 17731
rect 16405 17697 16439 17731
rect 16497 17697 16531 17731
rect 16589 17697 16623 17731
rect 16773 17697 16807 17731
rect 17233 17697 17267 17731
rect 20545 17697 20579 17731
rect 20637 17697 20671 17731
rect 20729 17697 20763 17731
rect 20913 17697 20947 17731
rect 21925 17697 21959 17731
rect 22201 17697 22235 17731
rect 23213 17697 23247 17731
rect 23397 17697 23431 17731
rect 24409 17697 24443 17731
rect 24501 17697 24535 17731
rect 24593 17697 24627 17731
rect 24777 17697 24811 17731
rect 24869 17697 24903 17731
rect 24961 17697 24995 17731
rect 27537 17719 27571 17753
rect 27629 17697 27663 17731
rect 27813 17697 27847 17731
rect 27905 17697 27939 17731
rect 29285 17697 29319 17731
rect 30297 17697 30331 17731
rect 30481 17697 30515 17731
rect 11713 17629 11747 17663
rect 11897 17629 11931 17663
rect 11989 17629 12023 17663
rect 12173 17629 12207 17663
rect 12817 17629 12851 17663
rect 22084 17629 22118 17663
rect 22937 17629 22971 17663
rect 23121 17629 23155 17663
rect 28825 17629 28859 17663
rect 29469 17629 29503 17663
rect 9965 17561 9999 17595
rect 13185 17561 13219 17595
rect 13829 17561 13863 17595
rect 17049 17561 17083 17595
rect 21281 17561 21315 17595
rect 22477 17561 22511 17595
rect 28089 17561 28123 17595
rect 28917 17561 28951 17595
rect 3893 17493 3927 17527
rect 4077 17493 4111 17527
rect 6101 17493 6135 17527
rect 7021 17493 7055 17527
rect 8677 17493 8711 17527
rect 9781 17493 9815 17527
rect 10333 17493 10367 17527
rect 12449 17493 12483 17527
rect 15669 17493 15703 17527
rect 20269 17493 20303 17527
rect 23581 17493 23615 17527
rect 28181 17493 28215 17527
rect 29745 17493 29779 17527
rect 30573 17493 30607 17527
rect 2421 17289 2455 17323
rect 3249 17289 3283 17323
rect 4353 17289 4387 17323
rect 7481 17289 7515 17323
rect 7665 17289 7699 17323
rect 16865 17289 16899 17323
rect 21005 17289 21039 17323
rect 29285 17289 29319 17323
rect 3709 17221 3743 17255
rect 7941 17221 7975 17255
rect 21281 17221 21315 17255
rect 6561 17153 6595 17187
rect 10609 17153 10643 17187
rect 12725 17153 12759 17187
rect 13645 17153 13679 17187
rect 17785 17153 17819 17187
rect 22661 17153 22695 17187
rect 23581 17153 23615 17187
rect 24409 17153 24443 17187
rect 25421 17153 25455 17187
rect 30665 17153 30699 17187
rect 2697 17085 2731 17119
rect 2789 17085 2823 17119
rect 2881 17085 2915 17119
rect 3065 17085 3099 17119
rect 3433 17085 3467 17119
rect 3525 17085 3559 17119
rect 4169 17085 4203 17119
rect 4353 17085 4387 17119
rect 7941 17085 7975 17119
rect 8125 17085 8159 17119
rect 10057 17085 10091 17119
rect 10149 17085 10183 17119
rect 10333 17085 10367 17119
rect 10425 17085 10459 17119
rect 10701 17085 10735 17119
rect 12449 17085 12483 17119
rect 12541 17085 12575 17119
rect 12633 17085 12667 17119
rect 13001 17085 13035 17119
rect 15025 17085 15059 17119
rect 15117 17085 15151 17119
rect 15209 17085 15243 17119
rect 15393 17085 15427 17119
rect 15485 17085 15519 17119
rect 15761 17085 15795 17119
rect 17693 17085 17727 17119
rect 20177 17085 20211 17119
rect 20361 17085 20395 17119
rect 20453 17085 20487 17119
rect 20545 17085 20579 17119
rect 20729 17085 20763 17119
rect 21189 17085 21223 17119
rect 22753 17085 22787 17119
rect 22937 17085 22971 17119
rect 23029 17085 23063 17119
rect 23121 17085 23155 17119
rect 23673 17085 23707 17119
rect 24961 17085 24995 17119
rect 25145 17085 25179 17119
rect 26065 17085 26099 17119
rect 26249 17085 26283 17119
rect 26341 17085 26375 17119
rect 26433 17085 26467 17119
rect 27905 17085 27939 17119
rect 28181 17085 28215 17119
rect 28365 17085 28399 17119
rect 28457 17085 28491 17119
rect 28549 17085 28583 17119
rect 29193 17085 29227 17119
rect 3249 17017 3283 17051
rect 7389 17017 7423 17051
rect 7849 17017 7883 17051
rect 14473 17017 14507 17051
rect 22416 17017 22450 17051
rect 23397 17017 23431 17051
rect 24317 17017 24351 17051
rect 24777 17017 24811 17051
rect 25513 17017 25547 17051
rect 25605 17017 25639 17051
rect 26709 17017 26743 17051
rect 27721 17017 27755 17051
rect 28825 17017 28859 17051
rect 30398 17017 30432 17051
rect 7649 16949 7683 16983
rect 9873 16949 9907 16983
rect 12909 16949 12943 16983
rect 14749 16949 14783 16983
rect 17233 16949 17267 16983
rect 17601 16949 17635 16983
rect 19993 16949 20027 16983
rect 23857 16949 23891 16983
rect 24225 16949 24259 16983
rect 25973 16949 26007 16983
rect 28089 16949 28123 16983
rect 29101 16949 29135 16983
rect 2237 16745 2271 16779
rect 4905 16745 4939 16779
rect 8585 16745 8619 16779
rect 15577 16745 15611 16779
rect 16129 16745 16163 16779
rect 16497 16745 16531 16779
rect 16589 16745 16623 16779
rect 17417 16745 17451 16779
rect 18521 16745 18555 16779
rect 25605 16745 25639 16779
rect 30389 16745 30423 16779
rect 1869 16677 1903 16711
rect 2053 16677 2087 16711
rect 2329 16677 2363 16711
rect 6285 16677 6319 16711
rect 8401 16677 8435 16711
rect 13645 16677 13679 16711
rect 19165 16677 19199 16711
rect 22109 16677 22143 16711
rect 26433 16677 26467 16711
rect 29929 16677 29963 16711
rect 1593 16609 1627 16643
rect 3065 16609 3099 16643
rect 3249 16609 3283 16643
rect 4261 16609 4295 16643
rect 7113 16609 7147 16643
rect 7297 16609 7331 16643
rect 8217 16609 8251 16643
rect 8493 16609 8527 16643
rect 8677 16609 8711 16643
rect 9505 16609 9539 16643
rect 9689 16609 9723 16643
rect 10517 16609 10551 16643
rect 12817 16609 12851 16643
rect 12909 16609 12943 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 17141 16609 17175 16643
rect 17233 16609 17267 16643
rect 17417 16609 17451 16643
rect 18797 16609 18831 16643
rect 19257 16609 19291 16643
rect 19441 16609 19475 16643
rect 21281 16609 21315 16643
rect 22753 16609 22787 16643
rect 23305 16609 23339 16643
rect 23397 16609 23431 16643
rect 23489 16609 23523 16643
rect 23685 16609 23719 16643
rect 24225 16609 24259 16643
rect 24492 16609 24526 16643
rect 25697 16609 25731 16643
rect 25789 16609 25823 16643
rect 25973 16609 26007 16643
rect 26065 16609 26099 16643
rect 26709 16609 26743 16643
rect 26801 16609 26835 16643
rect 26893 16609 26927 16643
rect 27077 16609 27111 16643
rect 27445 16609 27479 16643
rect 27629 16609 27663 16643
rect 27721 16609 27755 16643
rect 27813 16609 27847 16643
rect 28181 16609 28215 16643
rect 28437 16609 28471 16643
rect 30021 16609 30055 16643
rect 30481 16609 30515 16643
rect 30573 16609 30607 16643
rect 30757 16609 30791 16643
rect 30849 16609 30883 16643
rect 2973 16541 3007 16575
rect 3985 16541 4019 16575
rect 4102 16541 4136 16575
rect 8033 16541 8067 16575
rect 8125 16541 8159 16575
rect 9873 16541 9907 16575
rect 10241 16541 10275 16575
rect 16773 16541 16807 16575
rect 18685 16541 18719 16575
rect 19073 16541 19107 16575
rect 20177 16541 20211 16575
rect 20315 16541 20349 16575
rect 20453 16541 20487 16575
rect 26249 16541 26283 16575
rect 28089 16541 28123 16575
rect 29745 16541 29779 16575
rect 31033 16541 31067 16575
rect 3709 16473 3743 16507
rect 10425 16473 10459 16507
rect 19901 16473 19935 16507
rect 1685 16405 1719 16439
rect 9781 16405 9815 16439
rect 9965 16405 9999 16439
rect 17049 16405 17083 16439
rect 21097 16405 21131 16439
rect 23029 16405 23063 16439
rect 29561 16405 29595 16439
rect 3065 16201 3099 16235
rect 8125 16201 8159 16235
rect 9505 16201 9539 16235
rect 9873 16201 9907 16235
rect 10057 16201 10091 16235
rect 10425 16201 10459 16235
rect 11253 16201 11287 16235
rect 16221 16201 16255 16235
rect 22661 16201 22695 16235
rect 24501 16201 24535 16235
rect 26157 16201 26191 16235
rect 28825 16201 28859 16235
rect 29653 16201 29687 16235
rect 6745 16133 6779 16167
rect 9321 16133 9355 16167
rect 10333 16133 10367 16167
rect 11069 16133 11103 16167
rect 15761 16133 15795 16167
rect 22017 16133 22051 16167
rect 16589 16065 16623 16099
rect 16681 16065 16715 16099
rect 21373 16065 21407 16099
rect 21557 16065 21591 16099
rect 1409 15997 1443 16031
rect 1501 15997 1535 16031
rect 1685 15997 1719 16031
rect 3341 15997 3375 16031
rect 4261 15997 4295 16031
rect 4353 15997 4387 16031
rect 4445 15997 4479 16031
rect 4629 15997 4663 16031
rect 7481 15997 7515 16031
rect 7665 15997 7699 16031
rect 7757 15997 7791 16031
rect 7849 15997 7883 16031
rect 7941 15997 7975 16031
rect 9597 15997 9631 16031
rect 9965 15997 9999 16031
rect 10609 15997 10643 16031
rect 10701 15997 10735 16031
rect 10885 15997 10919 16031
rect 10977 15997 11011 16031
rect 12357 15997 12391 16031
rect 12541 15997 12575 16031
rect 12633 15997 12667 16031
rect 12725 15997 12759 16031
rect 13185 15997 13219 16031
rect 13277 15997 13311 16031
rect 13553 15997 13587 16031
rect 15577 15997 15611 16031
rect 15761 15997 15795 16031
rect 16465 15997 16499 16031
rect 18705 15997 18739 16031
rect 18797 15997 18831 16031
rect 18981 15997 19015 16031
rect 19248 15997 19282 16031
rect 20545 15997 20579 16031
rect 20729 15997 20763 16031
rect 20821 15997 20855 16031
rect 20913 15997 20947 16031
rect 22109 15997 22143 16031
rect 22201 15997 22235 16031
rect 22385 15997 22419 16031
rect 22477 15997 22511 16031
rect 22753 15997 22787 16031
rect 23121 15997 23155 16031
rect 23213 15997 23247 16031
rect 23397 15997 23431 16031
rect 23489 15997 23523 16031
rect 23857 15997 23891 16031
rect 24041 15997 24075 16031
rect 24133 15997 24167 16031
rect 24225 15997 24259 16031
rect 24777 15997 24811 16031
rect 25044 15997 25078 16031
rect 27629 15997 27663 16031
rect 28181 15997 28215 16031
rect 28365 15997 28399 16031
rect 28457 15997 28491 16031
rect 28549 15997 28583 16031
rect 29009 15997 29043 16031
rect 29193 15997 29227 16031
rect 29285 15997 29319 16031
rect 29377 15997 29411 16031
rect 29929 15997 29963 16031
rect 1952 15929 1986 15963
rect 6745 15929 6779 15963
rect 9045 15929 9079 15963
rect 11437 15929 11471 15963
rect 13001 15929 13035 15963
rect 13798 15929 13832 15963
rect 16129 15929 16163 15963
rect 17049 15929 17083 15963
rect 17509 15929 17543 15963
rect 17877 15929 17911 15963
rect 21189 15929 21223 15963
rect 23673 15929 23707 15963
rect 26617 15929 26651 15963
rect 27353 15929 27387 15963
rect 29745 15929 29779 15963
rect 30113 15929 30147 15963
rect 3893 15861 3927 15895
rect 3985 15861 4019 15895
rect 7205 15861 7239 15895
rect 7297 15861 7331 15895
rect 9689 15861 9723 15895
rect 11237 15861 11271 15895
rect 14933 15861 14967 15895
rect 17141 15861 17175 15895
rect 20361 15861 20395 15895
rect 21649 15861 21683 15895
rect 22937 15861 22971 15895
rect 3433 15657 3467 15691
rect 4537 15657 4571 15691
rect 14197 15657 14231 15691
rect 16129 15657 16163 15691
rect 18245 15657 18279 15691
rect 19073 15657 19107 15691
rect 19165 15657 19199 15691
rect 20545 15657 20579 15691
rect 20913 15657 20947 15691
rect 22293 15657 22327 15691
rect 22661 15657 22695 15691
rect 24961 15657 24995 15691
rect 2228 15589 2262 15623
rect 4169 15589 4203 15623
rect 4353 15589 4387 15623
rect 7113 15589 7147 15623
rect 9597 15589 9631 15623
rect 10701 15589 10735 15623
rect 20269 15589 20303 15623
rect 26433 15589 26467 15623
rect 27629 15589 27663 15623
rect 28825 15589 28859 15623
rect 1961 15521 1995 15555
rect 3709 15521 3743 15555
rect 3801 15521 3835 15555
rect 3893 15521 3927 15555
rect 4077 15521 4111 15555
rect 7665 15521 7699 15555
rect 7849 15521 7883 15555
rect 10425 15521 10459 15555
rect 10609 15521 10643 15555
rect 11529 15521 11563 15555
rect 14381 15521 14415 15555
rect 14657 15521 14691 15555
rect 16313 15521 16347 15555
rect 16589 15521 16623 15555
rect 16865 15521 16899 15555
rect 17121 15521 17155 15555
rect 18521 15521 18555 15555
rect 18889 15521 18923 15555
rect 19349 15521 19383 15555
rect 19533 15521 19567 15555
rect 19809 15521 19843 15555
rect 20729 15521 20763 15555
rect 21005 15521 21039 15555
rect 21465 15521 21499 15555
rect 21649 15521 21683 15555
rect 21833 15521 21867 15555
rect 22109 15521 22143 15555
rect 22845 15521 22879 15555
rect 24041 15521 24075 15555
rect 24225 15521 24259 15555
rect 24869 15521 24903 15555
rect 25237 15521 25271 15555
rect 26157 15521 26191 15555
rect 27169 15521 27203 15555
rect 27813 15521 27847 15555
rect 28181 15521 28215 15555
rect 28273 15521 28307 15555
rect 28457 15521 28491 15555
rect 28549 15521 28583 15555
rect 29101 15521 29135 15555
rect 29193 15521 29227 15555
rect 29290 15521 29324 15555
rect 29469 15521 29503 15555
rect 5549 15453 5583 15487
rect 6193 15453 6227 15487
rect 10057 15453 10091 15487
rect 18429 15453 18463 15487
rect 20453 15453 20487 15487
rect 3341 15385 3375 15419
rect 7389 15385 7423 15419
rect 9965 15385 9999 15419
rect 10241 15385 10275 15419
rect 14565 15385 14599 15419
rect 21281 15385 21315 15419
rect 4997 15317 5031 15351
rect 6837 15317 6871 15351
rect 7573 15317 7607 15351
rect 7757 15317 7791 15351
rect 12081 15317 12115 15351
rect 16497 15317 16531 15351
rect 18797 15317 18831 15351
rect 19717 15317 19751 15351
rect 21925 15317 21959 15351
rect 24409 15317 24443 15351
rect 25513 15317 25547 15351
rect 27997 15317 28031 15351
rect 28733 15317 28767 15351
rect 5457 15113 5491 15147
rect 9965 15113 9999 15147
rect 15393 15113 15427 15147
rect 16405 15113 16439 15147
rect 29101 15113 29135 15147
rect 30297 15113 30331 15147
rect 6285 15045 6319 15079
rect 9781 15045 9815 15079
rect 10057 15045 10091 15079
rect 16037 15045 16071 15079
rect 16681 15045 16715 15079
rect 18429 15045 18463 15079
rect 21189 15045 21223 15079
rect 22385 15045 22419 15079
rect 4813 14977 4847 15011
rect 6101 14977 6135 15011
rect 6745 14977 6779 15011
rect 6837 14977 6871 15011
rect 10517 14977 10551 15011
rect 11529 14977 11563 15011
rect 11621 14977 11655 15011
rect 14013 14977 14047 15011
rect 17785 14977 17819 15011
rect 22293 14977 22327 15011
rect 26617 14977 26651 15011
rect 29653 14977 29687 15011
rect 1961 14909 1995 14943
rect 2513 14909 2547 14943
rect 2605 14909 2639 14943
rect 2697 14909 2731 14943
rect 2881 14909 2915 14943
rect 3249 14909 3283 14943
rect 4353 14909 4387 14943
rect 4629 14909 4663 14943
rect 5365 14909 5399 14943
rect 5917 14909 5951 14943
rect 7849 14909 7883 14943
rect 8033 14909 8067 14943
rect 8217 14909 8251 14943
rect 9505 14909 9539 14943
rect 10241 14909 10275 14943
rect 10425 14909 10459 14943
rect 10609 14909 10643 14943
rect 10793 14909 10827 14943
rect 10977 14909 11011 14943
rect 11345 14909 11379 14943
rect 11805 14909 11839 14943
rect 13645 14909 13679 14943
rect 15761 14909 15795 14943
rect 16037 14909 16071 14943
rect 16405 14909 16439 14943
rect 16589 14909 16623 14943
rect 16957 14909 16991 14943
rect 17049 14909 17083 14943
rect 17141 14909 17175 14943
rect 17325 14909 17359 14943
rect 17601 14909 17635 14943
rect 18245 14909 18279 14943
rect 21005 14909 21039 14943
rect 22017 14909 22051 14943
rect 22661 14909 22695 14943
rect 22845 14909 22879 14943
rect 22937 14909 22971 14943
rect 23213 14909 23247 14943
rect 24225 14909 24259 14943
rect 24317 14909 24351 14943
rect 24409 14909 24443 14943
rect 24593 14909 24627 14943
rect 24961 14909 24995 14943
rect 25053 14909 25087 14943
rect 25237 14909 25271 14943
rect 25329 14909 25363 14943
rect 27169 14909 27203 14943
rect 27261 14909 27295 14943
rect 27445 14909 27479 14943
rect 27537 14909 27571 14943
rect 28641 14909 28675 14943
rect 29561 14909 29595 14943
rect 30113 14909 30147 14943
rect 30481 14909 30515 14943
rect 30665 14909 30699 14943
rect 30757 14909 30791 14943
rect 30849 14909 30883 14943
rect 3893 14841 3927 14875
rect 4169 14841 4203 14875
rect 8125 14841 8159 14875
rect 14280 14841 14314 14875
rect 17417 14841 17451 14875
rect 17969 14841 18003 14875
rect 20821 14841 20855 14875
rect 23029 14841 23063 14875
rect 29929 14841 29963 14875
rect 1869 14773 1903 14807
rect 2237 14773 2271 14807
rect 3985 14773 4019 14807
rect 4537 14773 4571 14807
rect 5825 14773 5859 14807
rect 6653 14773 6687 14807
rect 7297 14773 7331 14807
rect 11345 14773 11379 14807
rect 11989 14773 12023 14807
rect 13829 14773 13863 14807
rect 18061 14773 18095 14807
rect 23397 14773 23431 14807
rect 23949 14773 23983 14807
rect 25513 14773 25547 14807
rect 26065 14773 26099 14807
rect 26985 14773 27019 14807
rect 27997 14773 28031 14807
rect 29469 14773 29503 14807
rect 31125 14773 31159 14807
rect 5549 14569 5583 14603
rect 7113 14569 7147 14603
rect 11437 14569 11471 14603
rect 12265 14569 12299 14603
rect 13277 14569 13311 14603
rect 14381 14569 14415 14603
rect 16773 14569 16807 14603
rect 18521 14569 18555 14603
rect 19073 14569 19107 14603
rect 19165 14569 19199 14603
rect 20729 14569 20763 14603
rect 24501 14569 24535 14603
rect 27905 14569 27939 14603
rect 29377 14569 29411 14603
rect 1952 14501 1986 14535
rect 4436 14501 4470 14535
rect 7021 14501 7055 14535
rect 10793 14501 10827 14535
rect 11897 14501 11931 14535
rect 12097 14501 12131 14535
rect 14841 14501 14875 14535
rect 21465 14501 21499 14535
rect 24869 14501 24903 14535
rect 1685 14433 1719 14467
rect 3433 14433 3467 14467
rect 3525 14433 3559 14467
rect 3617 14433 3651 14467
rect 3801 14433 3835 14467
rect 4169 14433 4203 14467
rect 6009 14433 6043 14467
rect 6561 14433 6595 14467
rect 7849 14433 7883 14467
rect 10425 14433 10459 14467
rect 10609 14433 10643 14467
rect 11253 14433 11287 14467
rect 11345 14433 11379 14467
rect 11713 14433 11747 14467
rect 13093 14433 13127 14467
rect 13737 14433 13771 14467
rect 13921 14433 13955 14467
rect 14013 14433 14047 14467
rect 14105 14433 14139 14467
rect 14657 14433 14691 14467
rect 16221 14433 16255 14467
rect 16589 14433 16623 14467
rect 18153 14433 18187 14467
rect 18307 14433 18341 14467
rect 18981 14433 19015 14467
rect 20545 14433 20579 14467
rect 20821 14433 20855 14467
rect 20913 14433 20947 14467
rect 22661 14433 22695 14467
rect 23029 14433 23063 14467
rect 23581 14433 23615 14467
rect 23673 14433 23707 14467
rect 23765 14433 23799 14467
rect 23949 14433 23983 14467
rect 24409 14433 24443 14467
rect 25881 14433 25915 14467
rect 25973 14433 26007 14467
rect 26065 14433 26099 14467
rect 26249 14433 26283 14467
rect 26709 14433 26743 14467
rect 26801 14433 26835 14467
rect 26893 14433 26927 14467
rect 27077 14433 27111 14467
rect 27169 14433 27203 14467
rect 27353 14433 27387 14467
rect 27445 14433 27479 14467
rect 27537 14433 27571 14467
rect 28181 14433 28215 14467
rect 28273 14433 28307 14467
rect 28365 14433 28399 14467
rect 28549 14433 28583 14467
rect 29285 14433 29319 14467
rect 30481 14433 30515 14467
rect 30665 14433 30699 14467
rect 30757 14433 30791 14467
rect 30849 14433 30883 14467
rect 6101 14365 6135 14399
rect 6377 14365 6411 14399
rect 7205 14365 7239 14399
rect 7941 14365 7975 14399
rect 8033 14365 8067 14399
rect 14473 14365 14507 14399
rect 17601 14365 17635 14399
rect 19349 14365 19383 14399
rect 22201 14365 22235 14399
rect 24685 14365 24719 14399
rect 25421 14365 25455 14399
rect 29561 14365 29595 14399
rect 30297 14365 30331 14399
rect 3065 14297 3099 14331
rect 17969 14297 18003 14331
rect 18061 14297 18095 14331
rect 26433 14297 26467 14331
rect 27813 14297 27847 14331
rect 3157 14229 3191 14263
rect 6653 14229 6687 14263
rect 7481 14229 7515 14263
rect 12081 14229 12115 14263
rect 16405 14229 16439 14263
rect 19073 14229 19107 14263
rect 22477 14229 22511 14263
rect 22937 14229 22971 14263
rect 23305 14229 23339 14263
rect 24041 14229 24075 14263
rect 25605 14229 25639 14263
rect 28917 14229 28951 14263
rect 29745 14229 29779 14263
rect 31125 14229 31159 14263
rect 3065 14025 3099 14059
rect 5641 14025 5675 14059
rect 12081 14025 12115 14059
rect 12265 14025 12299 14059
rect 15945 14025 15979 14059
rect 18061 14025 18095 14059
rect 21005 14025 21039 14059
rect 23489 14025 23523 14059
rect 25237 14025 25271 14059
rect 26709 14025 26743 14059
rect 27169 14025 27203 14059
rect 29377 14025 29411 14059
rect 30941 14025 30975 14059
rect 11345 13957 11379 13991
rect 17877 13957 17911 13991
rect 22661 13957 22695 13991
rect 3801 13889 3835 13923
rect 5825 13889 5859 13923
rect 6285 13889 6319 13923
rect 9781 13889 9815 13923
rect 9965 13889 9999 13923
rect 20913 13889 20947 13923
rect 27629 13889 27663 13923
rect 27721 13889 27755 13923
rect 28825 13889 28859 13923
rect 1409 13821 1443 13855
rect 1501 13821 1535 13855
rect 1685 13821 1719 13855
rect 1952 13821 1986 13855
rect 3985 13821 4019 13855
rect 4077 13821 4111 13855
rect 4261 13821 4295 13855
rect 5733 13821 5767 13855
rect 6193 13821 6227 13855
rect 6552 13821 6586 13855
rect 9873 13821 9907 13855
rect 12633 13821 12667 13855
rect 12817 13821 12851 13855
rect 13093 13821 13127 13855
rect 13277 13821 13311 13855
rect 13829 13821 13863 13855
rect 14013 13821 14047 13855
rect 14105 13821 14139 13855
rect 14197 13821 14231 13855
rect 14565 13821 14599 13855
rect 16221 13821 16255 13855
rect 16497 13821 16531 13855
rect 17969 13821 18003 13855
rect 18153 13821 18187 13855
rect 20637 13821 20671 13855
rect 21281 13821 21315 13855
rect 22753 13821 22787 13855
rect 22845 13821 22879 13855
rect 23029 13821 23063 13855
rect 23673 13821 23707 13855
rect 23857 13821 23891 13855
rect 25329 13821 25363 13855
rect 25596 13821 25630 13855
rect 26893 13821 26927 13855
rect 27537 13821 27571 13855
rect 28181 13821 28215 13855
rect 28365 13821 28399 13855
rect 28457 13821 28491 13855
rect 28549 13821 28583 13855
rect 29193 13821 29227 13855
rect 29561 13821 29595 13855
rect 29828 13821 29862 13855
rect 31033 13821 31067 13855
rect 4528 13753 4562 13787
rect 10232 13753 10266 13787
rect 12449 13753 12483 13787
rect 14473 13753 14507 13787
rect 14810 13753 14844 13787
rect 16037 13753 16071 13787
rect 16764 13753 16798 13787
rect 21548 13753 21582 13787
rect 23213 13753 23247 13787
rect 24102 13753 24136 13787
rect 29009 13753 29043 13787
rect 3249 13685 3283 13719
rect 6101 13685 6135 13719
rect 7665 13685 7699 13719
rect 12249 13685 12283 13719
rect 12633 13685 12667 13719
rect 16405 13685 16439 13719
rect 26985 13685 27019 13719
rect 31125 13685 31159 13719
rect 2881 13481 2915 13515
rect 3893 13481 3927 13515
rect 13093 13481 13127 13515
rect 14841 13481 14875 13515
rect 15485 13481 15519 13515
rect 15761 13481 15795 13515
rect 16865 13481 16899 13515
rect 17049 13481 17083 13515
rect 20637 13481 20671 13515
rect 21741 13481 21775 13515
rect 21909 13481 21943 13515
rect 22293 13481 22327 13515
rect 23765 13481 23799 13515
rect 24501 13481 24535 13515
rect 24869 13481 24903 13515
rect 25145 13481 25179 13515
rect 26065 13481 26099 13515
rect 26801 13481 26835 13515
rect 28549 13481 28583 13515
rect 29009 13481 29043 13515
rect 31309 13481 31343 13515
rect 2697 13413 2731 13447
rect 3709 13413 3743 13447
rect 6276 13413 6310 13447
rect 9505 13413 9539 13447
rect 15025 13413 15059 13447
rect 15209 13413 15243 13447
rect 22109 13413 22143 13447
rect 25513 13413 25547 13447
rect 25605 13413 25639 13447
rect 26617 13413 26651 13447
rect 27436 13413 27470 13447
rect 30306 13413 30340 13447
rect 2513 13345 2547 13379
rect 3525 13345 3559 13379
rect 3801 13345 3835 13379
rect 3985 13345 4019 13379
rect 6009 13345 6043 13379
rect 7849 13345 7883 13379
rect 8033 13345 8067 13379
rect 9137 13345 9171 13379
rect 9413 13345 9447 13379
rect 9873 13345 9907 13379
rect 10057 13345 10091 13379
rect 10333 13345 10367 13379
rect 11069 13345 11103 13379
rect 13369 13345 13403 13379
rect 13829 13345 13863 13379
rect 15301 13345 15335 13379
rect 15853 13345 15887 13379
rect 16221 13345 16255 13379
rect 16405 13345 16439 13379
rect 16497 13345 16531 13379
rect 16589 13345 16623 13379
rect 16957 13345 16991 13379
rect 19165 13345 19199 13379
rect 19625 13345 19659 13379
rect 20085 13345 20119 13379
rect 20361 13345 20395 13379
rect 21649 13345 21683 13379
rect 22385 13345 22419 13379
rect 23949 13345 23983 13379
rect 24041 13345 24075 13379
rect 24225 13345 24259 13379
rect 24317 13345 24351 13379
rect 24685 13345 24719 13379
rect 24777 13345 24811 13379
rect 26157 13345 26191 13379
rect 26433 13345 26467 13379
rect 27169 13345 27203 13379
rect 28917 13345 28951 13379
rect 30573 13345 30607 13379
rect 8585 13277 8619 13311
rect 8953 13277 8987 13311
rect 9045 13277 9079 13311
rect 14105 13277 14139 13311
rect 19809 13277 19843 13311
rect 20177 13277 20211 13311
rect 21097 13277 21131 13311
rect 21557 13277 21591 13311
rect 25697 13277 25731 13311
rect 30757 13277 30791 13311
rect 19441 13209 19475 13243
rect 20729 13209 20763 13243
rect 21281 13209 21315 13243
rect 29193 13209 29227 13243
rect 3433 13141 3467 13175
rect 7389 13141 7423 13175
rect 7941 13141 7975 13175
rect 9965 13141 9999 13175
rect 10517 13141 10551 13175
rect 11161 13141 11195 13175
rect 13737 13141 13771 13175
rect 14749 13141 14783 13175
rect 19073 13141 19107 13175
rect 19809 13141 19843 13175
rect 21465 13141 21499 13175
rect 21925 13141 21959 13175
rect 10241 12937 10275 12971
rect 14933 12937 14967 12971
rect 18889 12937 18923 12971
rect 19625 12937 19659 12971
rect 21649 12937 21683 12971
rect 29009 12937 29043 12971
rect 19165 12869 19199 12903
rect 20177 12869 20211 12903
rect 5549 12801 5583 12835
rect 6009 12801 6043 12835
rect 6101 12801 6135 12835
rect 8861 12801 8895 12835
rect 8953 12801 8987 12835
rect 13553 12801 13587 12835
rect 19073 12801 19107 12835
rect 19441 12801 19475 12835
rect 19809 12801 19843 12835
rect 21373 12801 21407 12835
rect 2237 12733 2271 12767
rect 2605 12733 2639 12767
rect 2789 12733 2823 12767
rect 7205 12733 7239 12767
rect 7665 12733 7699 12767
rect 7849 12733 7883 12767
rect 8585 12733 8619 12767
rect 9597 12733 9631 12767
rect 9873 12733 9907 12767
rect 11621 12733 11655 12767
rect 11805 12733 11839 12767
rect 11897 12733 11931 12767
rect 12725 12733 12759 12767
rect 13184 12733 13218 12767
rect 13277 12733 13311 12767
rect 16037 12733 16071 12767
rect 16313 12733 16347 12767
rect 16497 12733 16531 12767
rect 17049 12733 17083 12767
rect 18797 12733 18831 12767
rect 19717 12733 19751 12767
rect 19993 12733 20027 12767
rect 20085 12733 20119 12767
rect 20269 12733 20303 12767
rect 20821 12733 20855 12767
rect 21465 12733 21499 12767
rect 21649 12733 21683 12767
rect 29193 12733 29227 12767
rect 29285 12733 29319 12767
rect 29469 12733 29503 12767
rect 29561 12733 29595 12767
rect 2421 12665 2455 12699
rect 11354 12665 11388 12699
rect 13820 12665 13854 12699
rect 16865 12665 16899 12699
rect 20637 12665 20671 12699
rect 2145 12597 2179 12631
rect 5733 12597 5767 12631
rect 7665 12597 7699 12631
rect 10057 12597 10091 12631
rect 12633 12597 12667 12631
rect 12909 12597 12943 12631
rect 16313 12597 16347 12631
rect 17141 12597 17175 12631
rect 19073 12597 19107 12631
rect 20729 12597 20763 12631
rect 21189 12597 21223 12631
rect 3433 12393 3467 12427
rect 10609 12393 10643 12427
rect 13921 12393 13955 12427
rect 14381 12393 14415 12427
rect 17969 12393 18003 12427
rect 1869 12325 1903 12359
rect 2206 12325 2240 12359
rect 3801 12325 3835 12359
rect 8795 12325 8829 12359
rect 12716 12325 12750 12359
rect 19156 12325 19190 12359
rect 20545 12325 20579 12359
rect 30297 12325 30331 12359
rect 1685 12257 1719 12291
rect 1961 12257 1995 12291
rect 3617 12257 3651 12291
rect 3709 12257 3743 12291
rect 3939 12257 3973 12291
rect 6929 12257 6963 12291
rect 7113 12257 7147 12291
rect 7481 12257 7515 12291
rect 8033 12257 8067 12291
rect 8217 12257 8251 12291
rect 8309 12257 8343 12291
rect 8493 12257 8527 12291
rect 8585 12257 8619 12291
rect 8677 12257 8711 12291
rect 8953 12257 8987 12291
rect 9229 12257 9263 12291
rect 9597 12257 9631 12291
rect 9965 12257 9999 12291
rect 10149 12257 10183 12291
rect 10241 12257 10275 12291
rect 10333 12257 10367 12291
rect 11253 12257 11287 12291
rect 11529 12257 11563 12291
rect 12449 12257 12483 12291
rect 14289 12257 14323 12291
rect 14749 12257 14783 12291
rect 15025 12257 15059 12291
rect 15485 12257 15519 12291
rect 15669 12257 15703 12291
rect 15761 12257 15795 12291
rect 16405 12257 16439 12291
rect 16589 12257 16623 12291
rect 16856 12257 16890 12291
rect 18705 12257 18739 12291
rect 18889 12257 18923 12291
rect 20361 12257 20395 12291
rect 22385 12257 22419 12291
rect 22845 12257 22879 12291
rect 23029 12257 23063 12291
rect 23121 12257 23155 12291
rect 23213 12257 23247 12291
rect 23765 12257 23799 12291
rect 24133 12257 24167 12291
rect 28273 12257 28307 12291
rect 28549 12257 28583 12291
rect 29469 12257 29503 12291
rect 29561 12257 29595 12291
rect 29745 12257 29779 12291
rect 29837 12257 29871 12291
rect 1501 12189 1535 12223
rect 4077 12189 4111 12223
rect 11713 12189 11747 12223
rect 14565 12189 14599 12223
rect 14841 12189 14875 12223
rect 29101 12189 29135 12223
rect 30941 12189 30975 12223
rect 3341 12121 3375 12155
rect 7021 12121 7055 12155
rect 9045 12121 9079 12155
rect 15209 12121 15243 12155
rect 15853 12121 15887 12155
rect 20729 12121 20763 12155
rect 8125 12053 8159 12087
rect 9413 12053 9447 12087
rect 13829 12053 13863 12087
rect 14749 12053 14783 12087
rect 15577 12053 15611 12087
rect 16313 12053 16347 12087
rect 18613 12053 18647 12087
rect 20269 12053 20303 12087
rect 22293 12053 22327 12087
rect 23489 12053 23523 12087
rect 23673 12053 23707 12087
rect 24041 12053 24075 12087
rect 28181 12053 28215 12087
rect 29377 12053 29411 12087
rect 29745 12053 29779 12087
rect 29929 12053 29963 12087
rect 3985 11849 4019 11883
rect 10057 11849 10091 11883
rect 13829 11849 13863 11883
rect 16221 11849 16255 11883
rect 28825 11849 28859 11883
rect 23305 11781 23339 11815
rect 26433 11781 26467 11815
rect 26617 11781 26651 11815
rect 1501 11713 1535 11747
rect 1685 11713 1719 11747
rect 3893 11713 3927 11747
rect 4629 11713 4663 11747
rect 6837 11713 6871 11747
rect 19349 11713 19383 11747
rect 23857 11713 23891 11747
rect 29193 11713 29227 11747
rect 1593 11645 1627 11679
rect 3433 11645 3467 11679
rect 3755 11645 3789 11679
rect 4170 11623 4204 11657
rect 4491 11645 4525 11679
rect 6101 11645 6135 11679
rect 7021 11645 7055 11679
rect 7481 11645 7515 11679
rect 7665 11645 7699 11679
rect 8033 11645 8067 11679
rect 8125 11645 8159 11679
rect 8401 11645 8435 11679
rect 8657 11645 8691 11679
rect 11437 11645 11471 11679
rect 11621 11645 11655 11679
rect 11713 11645 11747 11679
rect 13001 11645 13035 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 14105 11645 14139 11679
rect 15577 11645 15611 11679
rect 15761 11645 15795 11679
rect 15853 11645 15887 11679
rect 15945 11645 15979 11679
rect 16497 11645 16531 11679
rect 18061 11645 18095 11679
rect 18153 11645 18187 11679
rect 18337 11645 18371 11679
rect 18981 11645 19015 11679
rect 19533 11645 19567 11679
rect 19717 11645 19751 11679
rect 19901 11645 19935 11679
rect 19993 11645 20027 11679
rect 20177 11645 20211 11679
rect 21005 11645 21039 11679
rect 21189 11645 21223 11679
rect 21281 11645 21315 11679
rect 21373 11645 21407 11679
rect 21741 11645 21775 11679
rect 24113 11645 24147 11679
rect 25329 11645 25363 11679
rect 25483 11645 25517 11679
rect 25789 11645 25823 11679
rect 25882 11645 25916 11679
rect 26295 11645 26329 11679
rect 26525 11645 26559 11679
rect 26801 11645 26835 11679
rect 26893 11645 26927 11679
rect 27169 11645 27203 11679
rect 27261 11645 27295 11679
rect 27445 11645 27479 11679
rect 29460 11645 29494 11679
rect 31217 11645 31251 11679
rect 1952 11577 1986 11611
rect 3249 11577 3283 11611
rect 3525 11577 3559 11611
rect 3617 11577 3651 11611
rect 4261 11577 4295 11611
rect 4353 11577 4387 11611
rect 11170 11577 11204 11611
rect 15301 11577 15335 11611
rect 18245 11577 18279 11611
rect 21649 11577 21683 11611
rect 21986 11577 22020 11611
rect 23489 11577 23523 11611
rect 23673 11577 23707 11611
rect 25697 11577 25731 11611
rect 26065 11577 26099 11611
rect 26157 11577 26191 11611
rect 27077 11577 27111 11611
rect 27690 11577 27724 11611
rect 30665 11577 30699 11611
rect 3065 11509 3099 11543
rect 6009 11509 6043 11543
rect 7205 11509 7239 11543
rect 7665 11509 7699 11543
rect 9781 11509 9815 11543
rect 13093 11509 13127 11543
rect 14013 11509 14047 11543
rect 15393 11509 15427 11543
rect 19165 11509 19199 11543
rect 19809 11509 19843 11543
rect 20085 11509 20119 11543
rect 23121 11509 23155 11543
rect 25237 11509 25271 11543
rect 30573 11509 30607 11543
rect 3709 11305 3743 11339
rect 7205 11305 7239 11339
rect 9229 11305 9263 11339
rect 10175 11305 10209 11339
rect 10977 11305 11011 11339
rect 21925 11305 21959 11339
rect 25513 11305 25547 11339
rect 28365 11305 28399 11339
rect 29193 11305 29227 11339
rect 5273 11237 5307 11271
rect 6092 11237 6126 11271
rect 9965 11237 9999 11271
rect 10793 11237 10827 11271
rect 15761 11237 15795 11271
rect 16374 11237 16408 11271
rect 22109 11237 22143 11271
rect 22293 11237 22327 11271
rect 22753 11237 22787 11271
rect 25973 11237 26007 11271
rect 2053 11169 2087 11203
rect 2596 11169 2630 11203
rect 5181 11169 5215 11203
rect 5365 11169 5399 11203
rect 5503 11169 5537 11203
rect 5825 11169 5859 11203
rect 8585 11169 8619 11203
rect 8677 11169 8711 11203
rect 8769 11169 8803 11203
rect 8887 11169 8921 11203
rect 9045 11169 9079 11203
rect 9321 11169 9355 11203
rect 10517 11169 10551 11203
rect 10609 11169 10643 11203
rect 11345 11169 11379 11203
rect 15669 11169 15703 11203
rect 15853 11169 15887 11203
rect 16129 11169 16163 11203
rect 17785 11169 17819 11203
rect 18981 11169 19015 11203
rect 21281 11169 21315 11203
rect 21465 11169 21499 11203
rect 22017 11169 22051 11203
rect 22477 11169 22511 11203
rect 23305 11169 23339 11203
rect 23489 11169 23523 11203
rect 23756 11169 23790 11203
rect 28089 11169 28123 11203
rect 28549 11169 28583 11203
rect 28825 11169 28859 11203
rect 29101 11169 29135 11203
rect 30306 11169 30340 11203
rect 30573 11169 30607 11203
rect 30757 11169 30791 11203
rect 2145 11101 2179 11135
rect 2329 11101 2363 11135
rect 5641 11101 5675 11135
rect 11437 11101 11471 11135
rect 11529 11101 11563 11135
rect 17693 11101 17727 11135
rect 19625 11101 19659 11135
rect 27997 11101 28031 11135
rect 28733 11101 28767 11135
rect 10333 11033 10367 11067
rect 10793 11033 10827 11067
rect 18153 11033 18187 11067
rect 25605 11033 25639 11067
rect 27721 11033 27755 11067
rect 4997 10965 5031 10999
rect 8401 10965 8435 10999
rect 10149 10965 10183 10999
rect 17509 10965 17543 10999
rect 21649 10965 21683 10999
rect 24869 10965 24903 10999
rect 28549 10965 28583 10999
rect 29009 10965 29043 10999
rect 31309 10965 31343 10999
rect 2513 10761 2547 10795
rect 5457 10761 5491 10795
rect 7389 10761 7423 10795
rect 8769 10761 8803 10795
rect 13185 10761 13219 10795
rect 15853 10761 15887 10795
rect 22109 10761 22143 10795
rect 23397 10761 23431 10795
rect 25881 10761 25915 10795
rect 29929 10761 29963 10795
rect 30665 10761 30699 10795
rect 31217 10761 31251 10795
rect 7205 10693 7239 10727
rect 30481 10693 30515 10727
rect 2881 10625 2915 10659
rect 5089 10625 5123 10659
rect 15393 10625 15427 10659
rect 16497 10625 16531 10659
rect 23857 10625 23891 10659
rect 26065 10625 26099 10659
rect 30113 10625 30147 10659
rect 2237 10557 2271 10591
rect 2697 10557 2731 10591
rect 5273 10557 5307 10591
rect 5549 10557 5583 10591
rect 5641 10557 5675 10591
rect 5825 10557 5859 10591
rect 7573 10557 7607 10591
rect 7849 10557 7883 10591
rect 9321 10557 9355 10591
rect 9505 10557 9539 10591
rect 9689 10557 9723 10591
rect 10241 10557 10275 10591
rect 12265 10557 12299 10591
rect 12541 10557 12575 10591
rect 12843 10557 12877 10591
rect 13001 10557 13035 10591
rect 13277 10557 13311 10591
rect 14105 10557 14139 10591
rect 14657 10557 14691 10591
rect 15209 10557 15243 10591
rect 16037 10557 16071 10591
rect 16221 10557 16255 10591
rect 16773 10557 16807 10591
rect 18245 10557 18279 10591
rect 18429 10557 18463 10591
rect 18705 10557 18739 10591
rect 18961 10557 18995 10591
rect 20453 10557 20487 10591
rect 20545 10557 20579 10591
rect 20729 10557 20763 10591
rect 22753 10557 22787 10591
rect 22937 10557 22971 10591
rect 23029 10557 23063 10591
rect 23121 10557 23155 10591
rect 24041 10557 24075 10591
rect 25329 10557 25363 10591
rect 25513 10557 25547 10591
rect 25697 10557 25731 10591
rect 25973 10557 26007 10591
rect 26249 10557 26283 10591
rect 26341 10557 26375 10591
rect 29653 10557 29687 10591
rect 30205 10557 30239 10591
rect 30941 10557 30975 10591
rect 31033 10557 31067 10591
rect 31217 10557 31251 10591
rect 6070 10489 6104 10523
rect 12357 10489 12391 10523
rect 12633 10489 12667 10523
rect 12725 10489 12759 10523
rect 16129 10489 16163 10523
rect 16339 10489 16373 10523
rect 20996 10489 21030 10523
rect 24225 10489 24259 10523
rect 25605 10489 25639 10523
rect 30649 10489 30683 10523
rect 30849 10489 30883 10523
rect 2145 10421 2179 10455
rect 7757 10421 7791 10455
rect 9873 10421 9907 10455
rect 10149 10421 10183 10455
rect 12081 10421 12115 10455
rect 13553 10421 13587 10455
rect 14749 10421 14783 10455
rect 15025 10421 15059 10455
rect 16681 10421 16715 10455
rect 18245 10421 18279 10455
rect 20085 10421 20119 10455
rect 26525 10421 26559 10455
rect 29101 10421 29135 10455
rect 5917 10217 5951 10251
rect 8585 10217 8619 10251
rect 14013 10217 14047 10251
rect 18889 10217 18923 10251
rect 21281 10217 21315 10251
rect 25697 10217 25731 10251
rect 26249 10217 26283 10251
rect 26893 10217 26927 10251
rect 29285 10217 29319 10251
rect 3939 10149 3973 10183
rect 6653 10149 6687 10183
rect 6863 10149 6897 10183
rect 12035 10149 12069 10183
rect 12173 10149 12207 10183
rect 12878 10149 12912 10183
rect 14832 10149 14866 10183
rect 18153 10149 18187 10183
rect 18291 10149 18325 10183
rect 22477 10149 22511 10183
rect 25421 10149 25455 10183
rect 1685 10081 1719 10115
rect 1961 10081 1995 10115
rect 2217 10081 2251 10115
rect 3617 10081 3651 10115
rect 3709 10081 3743 10115
rect 3801 10081 3835 10115
rect 4077 10081 4111 10115
rect 6101 10081 6135 10115
rect 6377 10081 6411 10115
rect 6561 10081 6595 10115
rect 6745 10081 6779 10115
rect 7205 10081 7239 10115
rect 7472 10081 7506 10115
rect 9790 10081 9824 10115
rect 10057 10081 10091 10115
rect 11161 10081 11195 10115
rect 11253 10081 11287 10115
rect 11437 10081 11471 10115
rect 11621 10081 11655 10115
rect 12265 10081 12299 10115
rect 12357 10081 12391 10115
rect 12633 10081 12667 10115
rect 14565 10081 14599 10115
rect 17969 10081 18003 10115
rect 18061 10081 18095 10115
rect 18981 10081 19015 10115
rect 21557 10081 21591 10115
rect 21649 10081 21683 10115
rect 21741 10081 21775 10115
rect 21925 10081 21959 10115
rect 22201 10081 22235 10115
rect 22661 10081 22695 10115
rect 25145 10081 25179 10115
rect 25329 10081 25363 10115
rect 25513 10081 25547 10115
rect 25789 10081 25823 10115
rect 25881 10081 25915 10115
rect 26065 10081 26099 10115
rect 26617 10081 26651 10115
rect 26985 10081 27019 10115
rect 28641 10081 28675 10115
rect 28825 10081 28859 10115
rect 29101 10081 29135 10115
rect 30490 10081 30524 10115
rect 31033 10081 31067 10115
rect 3433 10013 3467 10047
rect 6285 10013 6319 10047
rect 7021 10013 7055 10047
rect 11897 10013 11931 10047
rect 12541 10013 12575 10047
rect 18429 10013 18463 10047
rect 28917 10013 28951 10047
rect 30757 10013 30791 10047
rect 30941 10013 30975 10047
rect 28825 9945 28859 9979
rect 1777 9877 1811 9911
rect 3341 9877 3375 9911
rect 8677 9877 8711 9911
rect 10977 9877 11011 9911
rect 11805 9877 11839 9911
rect 15945 9877 15979 9911
rect 17785 9877 17819 9911
rect 22293 9877 22327 9911
rect 22845 9877 22879 9911
rect 26525 9877 26559 9911
rect 29377 9877 29411 9911
rect 1593 9673 1627 9707
rect 9137 9673 9171 9707
rect 13553 9673 13587 9707
rect 15945 9673 15979 9707
rect 25145 9673 25179 9707
rect 25605 9673 25639 9707
rect 27445 9673 27479 9707
rect 28641 9673 28675 9707
rect 3065 9605 3099 9639
rect 9045 9605 9079 9639
rect 23489 9605 23523 9639
rect 25697 9605 25731 9639
rect 26985 9605 27019 9639
rect 28365 9605 28399 9639
rect 1225 9537 1259 9571
rect 9229 9537 9263 9571
rect 16589 9537 16623 9571
rect 22109 9537 22143 9571
rect 26801 9537 26835 9571
rect 27261 9537 27295 9571
rect 30205 9537 30239 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3249 9469 3283 9503
rect 3709 9469 3743 9503
rect 3893 9469 3927 9503
rect 4169 9469 4203 9503
rect 4353 9469 4387 9503
rect 5273 9469 5307 9503
rect 5365 9469 5399 9503
rect 5549 9469 5583 9503
rect 7205 9469 7239 9503
rect 8401 9469 8435 9503
rect 8769 9469 8803 9503
rect 8861 9469 8895 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 10241 9469 10275 9503
rect 10333 9469 10367 9503
rect 10517 9469 10551 9503
rect 10784 9469 10818 9503
rect 11989 9469 12023 9503
rect 12245 9469 12279 9503
rect 14105 9469 14139 9503
rect 14473 9469 14507 9503
rect 16129 9469 16163 9503
rect 16221 9469 16255 9503
rect 16773 9469 16807 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 18889 9469 18923 9503
rect 19901 9469 19935 9503
rect 20085 9469 20119 9503
rect 20177 9469 20211 9503
rect 20269 9469 20303 9503
rect 20637 9469 20671 9503
rect 24225 9469 24259 9503
rect 24379 9469 24413 9503
rect 25053 9469 25087 9503
rect 25329 9469 25363 9503
rect 25421 9469 25455 9503
rect 26065 9469 26099 9503
rect 26525 9469 26559 9503
rect 26617 9469 26651 9503
rect 26709 9469 26743 9503
rect 27169 9469 27203 9503
rect 28089 9469 28123 9503
rect 28181 9469 28215 9503
rect 28365 9469 28399 9503
rect 29193 9469 29227 9503
rect 29929 9469 29963 9503
rect 30113 9469 30147 9503
rect 30297 9469 30331 9503
rect 1952 9401 1986 9435
rect 3387 9401 3421 9435
rect 3525 9401 3559 9435
rect 3617 9401 3651 9435
rect 5816 9401 5850 9435
rect 8539 9401 8573 9435
rect 8677 9401 8711 9435
rect 14718 9401 14752 9435
rect 16313 9401 16347 9435
rect 16431 9401 16465 9435
rect 17049 9401 17083 9435
rect 17386 9401 17420 9435
rect 20545 9401 20579 9435
rect 20882 9401 20916 9435
rect 22376 9401 22410 9435
rect 25881 9401 25915 9435
rect 26249 9401 26283 9435
rect 27445 9401 27479 9435
rect 28457 9401 28491 9435
rect 29377 9401 29411 9435
rect 3985 9333 4019 9367
rect 6929 9333 6963 9367
rect 7849 9333 7883 9367
rect 9597 9333 9631 9367
rect 11897 9333 11931 9367
rect 13369 9333 13403 9367
rect 15853 9333 15887 9367
rect 18521 9333 18555 9367
rect 18797 9333 18831 9367
rect 22017 9333 22051 9367
rect 24593 9333 24627 9367
rect 25973 9333 26007 9367
rect 26341 9333 26375 9367
rect 28657 9333 28691 9367
rect 28825 9333 28859 9367
rect 29101 9333 29135 9367
rect 1869 9129 1903 9163
rect 3525 9129 3559 9163
rect 7021 9129 7055 9163
rect 9505 9129 9539 9163
rect 10517 9129 10551 9163
rect 12173 9129 12207 9163
rect 13829 9129 13863 9163
rect 15393 9129 15427 9163
rect 17325 9129 17359 9163
rect 20821 9129 20855 9163
rect 21281 9129 21315 9163
rect 22477 9129 22511 9163
rect 25329 9129 25363 9163
rect 28917 9129 28951 9163
rect 3801 9061 3835 9095
rect 4031 9061 4065 9095
rect 4905 9061 4939 9095
rect 7389 9061 7423 9095
rect 7527 9061 7561 9095
rect 11621 9061 11655 9095
rect 11851 9061 11885 9095
rect 14381 9061 14415 9095
rect 14841 9061 14875 9095
rect 15071 9061 15105 9095
rect 21465 9061 21499 9095
rect 21741 9061 21775 9095
rect 23581 9061 23615 9095
rect 24961 9061 24995 9095
rect 26249 9061 26283 9095
rect 26433 9061 26467 9095
rect 26617 9061 26651 9095
rect 1961 8993 1995 9027
rect 2320 8993 2354 9027
rect 3709 8993 3743 9027
rect 3893 8993 3927 9027
rect 4169 8993 4203 9027
rect 5641 8993 5675 9027
rect 6745 8993 6779 9027
rect 7205 8993 7239 9027
rect 7297 8993 7331 9027
rect 7665 8993 7699 9027
rect 9321 8993 9355 9027
rect 9505 8993 9539 9027
rect 9781 8993 9815 9027
rect 10057 8993 10091 9027
rect 10149 8993 10183 9027
rect 10241 8993 10275 9027
rect 11529 8993 11563 9027
rect 11713 8993 11747 9027
rect 11989 8993 12023 9027
rect 12265 8993 12299 9027
rect 13737 8993 13771 9027
rect 14197 8993 14231 9027
rect 14565 8993 14599 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 15209 8993 15243 9027
rect 15393 8993 15427 9027
rect 15577 8993 15611 9027
rect 17417 8993 17451 9027
rect 17969 8993 18003 9027
rect 18236 8993 18270 9027
rect 20913 8993 20947 9027
rect 21649 8993 21683 9027
rect 22753 8993 22787 9027
rect 22845 8993 22879 9027
rect 22937 8993 22971 9027
rect 23121 8993 23155 9027
rect 23213 8993 23247 9027
rect 23306 8993 23340 9027
rect 24685 8993 24719 9027
rect 24778 8993 24812 9027
rect 25053 8993 25087 9027
rect 25191 8993 25225 9027
rect 25513 8993 25547 9027
rect 26985 8993 27019 9027
rect 27905 8993 27939 9027
rect 28457 8993 28491 9027
rect 30030 8993 30064 9027
rect 30297 8993 30331 9027
rect 2053 8925 2087 8959
rect 5917 8925 5951 8959
rect 9965 8925 9999 8959
rect 11345 8925 11379 8959
rect 14013 8925 14047 8959
rect 22385 8925 22419 8959
rect 24409 8925 24443 8959
rect 25973 8857 26007 8891
rect 3433 8789 3467 8823
rect 19349 8789 19383 8823
rect 23765 8789 23799 8823
rect 25605 8789 25639 8823
rect 25789 8789 25823 8823
rect 26893 8789 26927 8823
rect 2329 8585 2363 8619
rect 4721 8585 4755 8619
rect 6377 8585 6411 8619
rect 14013 8585 14047 8619
rect 18153 8585 18187 8619
rect 24501 8585 24535 8619
rect 27169 8585 27203 8619
rect 28825 8585 28859 8619
rect 29929 8585 29963 8619
rect 4905 8517 4939 8551
rect 7113 8517 7147 8551
rect 14197 8517 14231 8551
rect 23857 8517 23891 8551
rect 24593 8517 24627 8551
rect 6101 8449 6135 8483
rect 18705 8449 18739 8483
rect 19349 8449 19383 8483
rect 23673 8449 23707 8483
rect 25421 8449 25455 8483
rect 25789 8449 25823 8483
rect 29009 8449 29043 8483
rect 2513 8381 2547 8415
rect 2697 8381 2731 8415
rect 4537 8381 4571 8415
rect 4721 8381 4755 8415
rect 5273 8381 5307 8415
rect 6285 8381 6319 8415
rect 6377 8381 6411 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 7665 8381 7699 8415
rect 9321 8381 9355 8415
rect 11989 8381 12023 8415
rect 15945 8381 15979 8415
rect 18337 8381 18371 8415
rect 18429 8381 18463 8415
rect 18889 8381 18923 8415
rect 19073 8381 19107 8415
rect 19191 8381 19225 8415
rect 19441 8381 19475 8415
rect 19625 8381 19659 8415
rect 21005 8381 21039 8415
rect 22201 8381 22235 8415
rect 22293 8381 22327 8415
rect 22477 8381 22511 8415
rect 22569 8381 22603 8415
rect 22661 8381 22695 8415
rect 23029 8381 23063 8415
rect 23213 8381 23247 8415
rect 23305 8381 23339 8415
rect 23397 8381 23431 8415
rect 25697 8381 25731 8415
rect 27445 8381 27479 8415
rect 29745 8381 29779 8415
rect 29929 8381 29963 8415
rect 7757 8313 7791 8347
rect 13829 8313 13863 8347
rect 18981 8313 19015 8347
rect 24041 8313 24075 8347
rect 24225 8313 24259 8347
rect 24961 8313 24995 8347
rect 25053 8313 25087 8347
rect 25237 8313 25271 8347
rect 26034 8313 26068 8347
rect 27690 8313 27724 8347
rect 29653 8313 29687 8347
rect 9229 8245 9263 8279
rect 14013 8245 14047 8279
rect 15853 8245 15887 8279
rect 19809 8245 19843 8279
rect 20913 8245 20947 8279
rect 22109 8245 22143 8279
rect 22937 8245 22971 8279
rect 25605 8245 25639 8279
rect 5089 8041 5123 8075
rect 6929 8041 6963 8075
rect 10149 8041 10183 8075
rect 19349 8041 19383 8075
rect 24133 8041 24167 8075
rect 27169 8041 27203 8075
rect 27629 8041 27663 8075
rect 5273 7973 5307 8007
rect 6469 7973 6503 8007
rect 7389 7973 7423 8007
rect 11621 7973 11655 8007
rect 12817 7973 12851 8007
rect 19073 7973 19107 8007
rect 20554 7973 20588 8007
rect 2329 7905 2363 7939
rect 2881 7905 2915 7939
rect 4721 7905 4755 7939
rect 5181 7905 5215 7939
rect 6285 7905 6319 7939
rect 6561 7905 6595 7939
rect 6653 7905 6687 7939
rect 7113 7905 7147 7939
rect 7205 7905 7239 7939
rect 7665 7905 7699 7939
rect 7757 7905 7791 7939
rect 7849 7905 7883 7939
rect 8493 7905 8527 7939
rect 9780 7905 9814 7939
rect 9873 7905 9907 7939
rect 9965 7929 9999 7963
rect 11161 7905 11195 7939
rect 12357 7905 12391 7939
rect 12725 7905 12759 7939
rect 13001 7905 13035 7939
rect 13093 7905 13127 7939
rect 13186 7905 13220 7939
rect 13369 7905 13403 7939
rect 13461 7905 13495 7939
rect 13558 7905 13592 7939
rect 15025 7905 15059 7939
rect 15117 7905 15151 7939
rect 15301 7905 15335 7939
rect 15577 7905 15611 7939
rect 18705 7905 18739 7939
rect 18843 7905 18877 7939
rect 18981 7905 19015 7939
rect 19165 7905 19199 7939
rect 20821 7905 20855 7939
rect 22753 7905 22787 7939
rect 23020 7905 23054 7939
rect 24225 7905 24259 7939
rect 24481 7905 24515 7939
rect 26801 7905 26835 7939
rect 27721 7905 27755 7939
rect 2513 7837 2547 7871
rect 4629 7837 4663 7871
rect 8033 7837 8067 7871
rect 8585 7837 8619 7871
rect 11253 7837 11287 7871
rect 11529 7837 11563 7871
rect 14381 7837 14415 7871
rect 14749 7837 14783 7871
rect 15669 7837 15703 7871
rect 16773 7837 16807 7871
rect 26709 7837 26743 7871
rect 7481 7769 7515 7803
rect 8861 7769 8895 7803
rect 9045 7769 9079 7803
rect 9505 7769 9539 7803
rect 14933 7769 14967 7803
rect 16497 7769 16531 7803
rect 19441 7769 19475 7803
rect 25605 7769 25639 7803
rect 2145 7701 2179 7735
rect 2789 7701 2823 7735
rect 6837 7701 6871 7735
rect 7389 7701 7423 7735
rect 8401 7701 8435 7735
rect 13001 7701 13035 7735
rect 13737 7701 13771 7735
rect 13829 7701 13863 7735
rect 14841 7701 14875 7735
rect 15301 7701 15335 7735
rect 15853 7701 15887 7735
rect 16313 7701 16347 7735
rect 3249 7497 3283 7531
rect 6653 7497 6687 7531
rect 8033 7497 8067 7531
rect 8953 7497 8987 7531
rect 13921 7497 13955 7531
rect 14013 7497 14047 7531
rect 14289 7497 14323 7531
rect 14749 7497 14783 7531
rect 21649 7497 21683 7531
rect 3065 7429 3099 7463
rect 9597 7429 9631 7463
rect 13277 7429 13311 7463
rect 13829 7429 13863 7463
rect 4537 7361 4571 7395
rect 6193 7361 6227 7395
rect 6285 7361 6319 7395
rect 7573 7361 7607 7395
rect 8861 7361 8895 7395
rect 9413 7361 9447 7395
rect 9873 7361 9907 7395
rect 14841 7361 14875 7395
rect 16681 7361 16715 7395
rect 17049 7361 17083 7395
rect 18429 7361 18463 7395
rect 19165 7361 19199 7395
rect 21373 7361 21407 7395
rect 22293 7361 22327 7395
rect 1317 7293 1351 7327
rect 1409 7293 1443 7327
rect 1501 7293 1535 7327
rect 1685 7293 1719 7327
rect 1952 7293 1986 7327
rect 3433 7293 3467 7327
rect 3525 7293 3559 7327
rect 3893 7293 3927 7327
rect 4445 7293 4479 7327
rect 5917 7293 5951 7327
rect 6101 7293 6135 7327
rect 6469 7293 6503 7327
rect 7021 7293 7055 7327
rect 7297 7293 7331 7327
rect 7481 7293 7515 7327
rect 7665 7293 7699 7327
rect 7849 7293 7883 7327
rect 8585 7293 8619 7327
rect 8769 7293 8803 7327
rect 9045 7293 9079 7327
rect 10179 7293 10213 7327
rect 10333 7293 10367 7327
rect 10639 7293 10673 7327
rect 10793 7293 10827 7327
rect 11805 7293 11839 7327
rect 11897 7293 11931 7327
rect 13553 7293 13587 7327
rect 14565 7293 14599 7327
rect 14933 7293 14967 7327
rect 15026 7293 15060 7327
rect 15209 7293 15243 7327
rect 15439 7293 15473 7327
rect 15669 7293 15703 7327
rect 15853 7293 15887 7327
rect 15945 7293 15979 7327
rect 16037 7293 16071 7327
rect 16221 7293 16255 7327
rect 16773 7293 16807 7327
rect 17417 7293 17451 7327
rect 18337 7293 18371 7327
rect 18797 7293 18831 7327
rect 18889 7293 18923 7327
rect 20637 7293 20671 7327
rect 21833 7293 21867 7327
rect 22017 7293 22051 7327
rect 22569 7293 22603 7327
rect 26065 7293 26099 7327
rect 26709 7293 26743 7327
rect 29193 7293 29227 7327
rect 3617 7225 3651 7259
rect 3735 7225 3769 7259
rect 11069 7225 11103 7259
rect 12142 7225 12176 7259
rect 14381 7225 14415 7259
rect 15301 7225 15335 7259
rect 17141 7225 17175 7259
rect 17325 7225 17359 7259
rect 19073 7225 19107 7259
rect 19410 7225 19444 7259
rect 21925 7225 21959 7259
rect 22135 7225 22169 7259
rect 1225 7157 1259 7191
rect 4813 7157 4847 7191
rect 6929 7157 6963 7191
rect 9321 7157 9355 7191
rect 9965 7157 9999 7191
rect 10425 7157 10459 7191
rect 13645 7157 13679 7191
rect 15577 7157 15611 7191
rect 16405 7157 16439 7191
rect 16497 7157 16531 7191
rect 20545 7157 20579 7191
rect 22477 7157 22511 7191
rect 26249 7157 26283 7191
rect 26617 7157 26651 7191
rect 29101 7157 29135 7191
rect 6653 6953 6687 6987
rect 12081 6953 12115 6987
rect 15393 6953 15427 6987
rect 15485 6953 15519 6987
rect 25789 6953 25823 6987
rect 4445 6885 4479 6919
rect 4563 6885 4597 6919
rect 6745 6885 6779 6919
rect 7205 6885 7239 6919
rect 12357 6885 12391 6919
rect 15945 6885 15979 6919
rect 25881 6885 25915 6919
rect 26111 6851 26145 6885
rect 1133 6817 1167 6851
rect 1400 6817 1434 6851
rect 2605 6817 2639 6851
rect 2872 6817 2906 6851
rect 4261 6817 4295 6851
rect 4353 6817 4387 6851
rect 4721 6817 4755 6851
rect 6101 6817 6135 6851
rect 6377 6817 6411 6851
rect 6469 6817 6503 6851
rect 6561 6817 6595 6851
rect 6837 6817 6871 6851
rect 6929 6817 6963 6851
rect 7757 6817 7791 6851
rect 7850 6817 7884 6851
rect 8033 6817 8067 6851
rect 8125 6817 8159 6851
rect 8222 6817 8256 6851
rect 9229 6817 9263 6851
rect 9413 6817 9447 6851
rect 9597 6817 9631 6851
rect 9965 6817 9999 6851
rect 11069 6817 11103 6851
rect 12173 6817 12207 6851
rect 12541 6817 12575 6851
rect 12725 6817 12759 6851
rect 13001 6817 13035 6851
rect 13185 6817 13219 6851
rect 13277 6817 13311 6851
rect 13461 6817 13495 6851
rect 13645 6817 13679 6851
rect 13829 6817 13863 6851
rect 14197 6817 14231 6851
rect 14289 6817 14323 6851
rect 15025 6817 15059 6851
rect 15117 6817 15151 6851
rect 15239 6817 15273 6851
rect 15669 6817 15703 6851
rect 16405 6817 16439 6851
rect 16681 6817 16715 6851
rect 17877 6817 17911 6851
rect 17969 6817 18003 6851
rect 18245 6817 18279 6851
rect 18429 6817 18463 6851
rect 19634 6817 19668 6851
rect 20361 6817 20395 6851
rect 20637 6817 20671 6851
rect 20729 6817 20763 6851
rect 20913 6817 20947 6851
rect 21373 6817 21407 6851
rect 21557 6817 21591 6851
rect 21925 6817 21959 6851
rect 22109 6817 22143 6851
rect 22201 6817 22235 6851
rect 22457 6817 22491 6851
rect 25513 6817 25547 6851
rect 25697 6817 25731 6851
rect 25789 6817 25823 6851
rect 26433 6817 26467 6851
rect 26689 6817 26723 6851
rect 28089 6817 28123 6851
rect 28641 6817 28675 6851
rect 28908 6817 28942 6851
rect 30113 6817 30147 6851
rect 6193 6749 6227 6783
rect 7665 6749 7699 6783
rect 9873 6749 9907 6783
rect 10241 6749 10275 6783
rect 10333 6749 10367 6783
rect 12817 6749 12851 6783
rect 13553 6749 13587 6783
rect 14013 6749 14047 6783
rect 15393 6749 15427 6783
rect 15853 6749 15887 6783
rect 16313 6749 16347 6783
rect 16773 6749 16807 6783
rect 18061 6749 18095 6783
rect 19901 6749 19935 6783
rect 20545 6749 20579 6783
rect 21741 6749 21775 6783
rect 30665 6749 30699 6783
rect 4077 6681 4111 6715
rect 5917 6681 5951 6715
rect 7481 6681 7515 6715
rect 16129 6681 16163 6715
rect 26249 6681 26283 6715
rect 28365 6681 28399 6715
rect 2513 6613 2547 6647
rect 3985 6613 4019 6647
rect 6101 6613 6135 6647
rect 8401 6613 8435 6647
rect 8861 6613 8895 6647
rect 9137 6613 9171 6647
rect 9321 6613 9355 6647
rect 9689 6613 9723 6647
rect 13185 6613 13219 6647
rect 15945 6613 15979 6647
rect 18521 6613 18555 6647
rect 20913 6613 20947 6647
rect 21557 6613 21591 6647
rect 23581 6613 23615 6647
rect 26065 6613 26099 6647
rect 27813 6613 27847 6647
rect 28549 6613 28583 6647
rect 30021 6613 30055 6647
rect 1961 6409 1995 6443
rect 7665 6409 7699 6443
rect 9045 6409 9079 6443
rect 9965 6409 9999 6443
rect 18705 6409 18739 6443
rect 22201 6409 22235 6443
rect 28365 6409 28399 6443
rect 3249 6341 3283 6375
rect 6469 6341 6503 6375
rect 12173 6341 12207 6375
rect 29101 6341 29135 6375
rect 2329 6273 2363 6307
rect 3065 6273 3099 6307
rect 6653 6273 6687 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 8861 6273 8895 6307
rect 9597 6273 9631 6307
rect 9781 6273 9815 6307
rect 10057 6273 10091 6307
rect 19349 6273 19383 6307
rect 28181 6273 28215 6307
rect 2145 6205 2179 6239
rect 2605 6205 2639 6239
rect 2789 6205 2823 6239
rect 2927 6205 2961 6239
rect 3433 6205 3467 6239
rect 3525 6205 3559 6239
rect 3893 6205 3927 6239
rect 6193 6205 6227 6239
rect 6745 6205 6779 6239
rect 7573 6205 7607 6239
rect 8769 6205 8803 6239
rect 10333 6205 10367 6239
rect 12265 6205 12299 6239
rect 18889 6205 18923 6239
rect 18981 6205 19015 6239
rect 20361 6205 20395 6239
rect 21557 6205 21591 6239
rect 21715 6205 21749 6239
rect 22017 6205 22051 6239
rect 24685 6205 24719 6239
rect 24961 6205 24995 6239
rect 25053 6205 25087 6239
rect 25237 6205 25271 6239
rect 26709 6205 26743 6239
rect 27905 6205 27939 6239
rect 27997 6205 28031 6239
rect 28089 6205 28123 6239
rect 28549 6205 28583 6239
rect 28825 6205 28859 6239
rect 30481 6205 30515 6239
rect 2697 6137 2731 6171
rect 3617 6137 3651 6171
rect 3755 6137 3789 6171
rect 6837 6137 6871 6171
rect 9505 6137 9539 6171
rect 9689 6137 9723 6171
rect 19073 6137 19107 6171
rect 19191 6137 19225 6171
rect 19625 6137 19659 6171
rect 21833 6137 21867 6171
rect 21925 6137 21959 6171
rect 25504 6137 25538 6171
rect 27445 6137 27479 6171
rect 30214 6137 30248 6171
rect 2421 6069 2455 6103
rect 10241 6069 10275 6103
rect 26617 6069 26651 6103
rect 27721 6069 27755 6103
rect 28733 6069 28767 6103
rect 2789 5865 2823 5899
rect 9045 5865 9079 5899
rect 12449 5865 12483 5899
rect 14749 5865 14783 5899
rect 25605 5865 25639 5899
rect 25789 5865 25823 5899
rect 27813 5865 27847 5899
rect 29015 5865 29049 5899
rect 29929 5865 29963 5899
rect 30481 5865 30515 5899
rect 8677 5797 8711 5831
rect 8769 5797 8803 5831
rect 9137 5797 9171 5831
rect 9505 5797 9539 5831
rect 11437 5797 11471 5831
rect 13855 5797 13889 5831
rect 18705 5797 18739 5831
rect 18797 5797 18831 5831
rect 26433 5797 26467 5831
rect 27261 5797 27295 5831
rect 28825 5797 28859 5831
rect 28917 5797 28951 5831
rect 29101 5797 29135 5831
rect 1961 5729 1995 5763
rect 2237 5729 2271 5763
rect 2329 5729 2363 5763
rect 2973 5729 3007 5763
rect 3433 5729 3467 5763
rect 8401 5729 8435 5763
rect 8494 5729 8528 5763
rect 8907 5729 8941 5763
rect 9321 5729 9355 5763
rect 9597 5729 9631 5763
rect 9781 5729 9815 5763
rect 11345 5729 11379 5763
rect 11529 5729 11563 5763
rect 11667 5729 11701 5763
rect 12081 5729 12115 5763
rect 12909 5729 12943 5763
rect 13553 5729 13587 5763
rect 13645 5729 13679 5763
rect 13737 5729 13771 5763
rect 14013 5729 14047 5763
rect 14105 5729 14139 5763
rect 14243 5729 14277 5763
rect 14381 5729 14415 5763
rect 14473 5729 14507 5763
rect 14570 5729 14604 5763
rect 14841 5729 14875 5763
rect 14995 5729 15029 5763
rect 18613 5729 18647 5763
rect 18915 5729 18949 5763
rect 21557 5729 21591 5763
rect 22661 5729 22695 5763
rect 23121 5729 23155 5763
rect 25329 5729 25363 5763
rect 27629 5729 27663 5763
rect 27721 5729 27755 5763
rect 27997 5729 28031 5763
rect 28549 5729 28583 5763
rect 28641 5729 28675 5763
rect 29193 5729 29227 5763
rect 29377 5729 29411 5763
rect 30297 5729 30331 5763
rect 30389 5729 30423 5763
rect 3157 5661 3191 5695
rect 9689 5661 9723 5695
rect 11805 5661 11839 5695
rect 11989 5661 12023 5695
rect 13001 5661 13035 5695
rect 19073 5661 19107 5695
rect 22477 5661 22511 5695
rect 22937 5661 22971 5695
rect 28825 5661 28859 5695
rect 30021 5661 30055 5695
rect 13277 5593 13311 5627
rect 26157 5593 26191 5627
rect 30113 5593 30147 5627
rect 1869 5525 1903 5559
rect 2053 5525 2087 5559
rect 3341 5525 3375 5559
rect 11161 5525 11195 5559
rect 13369 5525 13403 5559
rect 15025 5525 15059 5559
rect 18429 5525 18463 5559
rect 21465 5525 21499 5559
rect 22845 5525 22879 5559
rect 23305 5525 23339 5559
rect 25789 5525 25823 5559
rect 27445 5525 27479 5559
rect 30205 5525 30239 5559
rect 3065 5321 3099 5355
rect 3525 5321 3559 5355
rect 4169 5321 4203 5355
rect 8125 5321 8159 5355
rect 8401 5321 8435 5355
rect 11805 5321 11839 5355
rect 12725 5321 12759 5355
rect 14197 5321 14231 5355
rect 17141 5321 17175 5355
rect 20085 5321 20119 5355
rect 22753 5321 22787 5355
rect 3893 5253 3927 5287
rect 3985 5253 4019 5287
rect 7573 5253 7607 5287
rect 30665 5253 30699 5287
rect 8861 5185 8895 5219
rect 13369 5185 13403 5219
rect 14565 5185 14599 5219
rect 16313 5185 16347 5219
rect 18153 5185 18187 5219
rect 18521 5185 18555 5219
rect 20821 5185 20855 5219
rect 21925 5185 21959 5219
rect 22661 5185 22695 5219
rect 23397 5185 23431 5219
rect 26065 5185 26099 5219
rect 26224 5185 26258 5219
rect 26341 5185 26375 5219
rect 26617 5185 26651 5219
rect 27077 5185 27111 5219
rect 27261 5185 27295 5219
rect 29929 5185 29963 5219
rect 1409 5117 1443 5151
rect 1501 5117 1535 5151
rect 1685 5117 1719 5151
rect 1952 5117 1986 5151
rect 7481 5117 7515 5151
rect 7665 5117 7699 5151
rect 8769 5117 8803 5151
rect 9321 5117 9355 5151
rect 10057 5117 10091 5151
rect 10149 5117 10183 5151
rect 10425 5117 10459 5151
rect 12909 5117 12943 5151
rect 13001 5117 13035 5151
rect 13093 5117 13127 5151
rect 13553 5117 13587 5151
rect 13737 5117 13771 5151
rect 14381 5117 14415 5151
rect 14657 5117 14691 5151
rect 14749 5117 14783 5151
rect 14933 5117 14967 5151
rect 15025 5117 15059 5151
rect 15853 5117 15887 5151
rect 16155 5117 16189 5151
rect 16589 5117 16623 5151
rect 17141 5117 17175 5151
rect 17325 5117 17359 5151
rect 18337 5117 18371 5151
rect 18712 5117 18746 5151
rect 18961 5117 18995 5151
rect 21005 5117 21039 5151
rect 21281 5117 21315 5151
rect 21465 5117 21499 5151
rect 21649 5117 21683 5151
rect 22017 5117 22051 5151
rect 22293 5117 22327 5151
rect 22477 5117 22511 5151
rect 22937 5117 22971 5151
rect 23121 5117 23155 5151
rect 23673 5117 23707 5151
rect 28089 5117 28123 5151
rect 28641 5117 28675 5151
rect 29377 5117 29411 5151
rect 29561 5117 29595 5151
rect 29653 5117 29687 5151
rect 30573 5117 30607 5151
rect 30665 5117 30699 5151
rect 30941 5117 30975 5151
rect 4353 5049 4387 5083
rect 7757 5049 7791 5083
rect 7941 5049 7975 5083
rect 10333 5049 10367 5083
rect 10670 5049 10704 5083
rect 13231 5049 13265 5083
rect 15945 5049 15979 5083
rect 16037 5049 16071 5083
rect 21557 5049 21591 5083
rect 21767 5049 21801 5083
rect 22155 5049 22189 5083
rect 22385 5049 22419 5083
rect 23029 5049 23063 5083
rect 23239 5049 23273 5083
rect 28181 5049 28215 5083
rect 30849 5049 30883 5083
rect 3341 4981 3375 5015
rect 3525 4981 3559 5015
rect 4153 4981 4187 5015
rect 9413 4981 9447 5015
rect 13921 4981 13955 5015
rect 15117 4981 15151 5015
rect 15669 4981 15703 5015
rect 16497 4981 16531 5015
rect 21189 4981 21223 5015
rect 23581 4981 23615 5015
rect 25421 4981 25455 5015
rect 28733 4981 28767 5015
rect 29193 4981 29227 5015
rect 3065 4777 3099 4811
rect 4629 4777 4663 4811
rect 4997 4777 5031 4811
rect 7389 4777 7423 4811
rect 10609 4777 10643 4811
rect 11069 4777 11103 4811
rect 13553 4777 13587 4811
rect 18889 4777 18923 4811
rect 25697 4777 25731 4811
rect 27905 4777 27939 4811
rect 29009 4777 29043 4811
rect 29193 4777 29227 4811
rect 30665 4777 30699 4811
rect 7665 4709 7699 4743
rect 7941 4709 7975 4743
rect 18429 4709 18463 4743
rect 18613 4709 18647 4743
rect 20545 4709 20579 4743
rect 21526 4709 21560 4743
rect 27997 4709 28031 4743
rect 29530 4709 29564 4743
rect 1685 4641 1719 4675
rect 1952 4641 1986 4675
rect 3157 4641 3191 4675
rect 3424 4641 3458 4675
rect 4813 4641 4847 4675
rect 5089 4641 5123 4675
rect 6193 4641 6227 4675
rect 7113 4641 7147 4675
rect 7297 4641 7331 4675
rect 7481 4641 7515 4675
rect 7849 4641 7883 4675
rect 10701 4641 10735 4675
rect 11161 4641 11195 4675
rect 13277 4641 13311 4675
rect 13461 4641 13495 4675
rect 14666 4641 14700 4675
rect 14933 4641 14967 4675
rect 15577 4641 15611 4675
rect 15761 4641 15795 4675
rect 16129 4641 16163 4675
rect 16385 4641 16419 4675
rect 17969 4641 18003 4675
rect 18981 4641 19015 4675
rect 20729 4641 20763 4675
rect 20821 4641 20855 4675
rect 21097 4641 21131 4675
rect 21281 4641 21315 4675
rect 23029 4641 23063 4675
rect 23285 4641 23319 4675
rect 28089 4641 28123 4675
rect 28365 4641 28399 4675
rect 28549 4641 28583 4675
rect 29285 4641 29319 4675
rect 13093 4573 13127 4607
rect 15945 4573 15979 4607
rect 17601 4573 17635 4607
rect 18061 4573 18095 4607
rect 25789 4573 25823 4607
rect 25881 4573 25915 4607
rect 27721 4573 27755 4607
rect 4537 4505 4571 4539
rect 28273 4505 28307 4539
rect 28641 4505 28675 4539
rect 6285 4437 6319 4471
rect 17509 4437 17543 4471
rect 18245 4437 18279 4471
rect 21005 4437 21039 4471
rect 22661 4437 22695 4471
rect 24409 4437 24443 4471
rect 25329 4437 25363 4471
rect 28549 4437 28583 4471
rect 29009 4437 29043 4471
rect 2697 4233 2731 4267
rect 2881 4233 2915 4267
rect 5089 4233 5123 4267
rect 6745 4233 6779 4267
rect 8217 4233 8251 4267
rect 8585 4233 8619 4267
rect 14933 4233 14967 4267
rect 16865 4233 16899 4267
rect 17785 4233 17819 4267
rect 20085 4233 20119 4267
rect 22017 4233 22051 4267
rect 26157 4233 26191 4267
rect 29009 4233 29043 4267
rect 29193 4233 29227 4267
rect 29469 4233 29503 4267
rect 17417 4165 17451 4199
rect 25421 4165 25455 4199
rect 27353 4165 27387 4199
rect 16405 4097 16439 4131
rect 21465 4097 21499 4131
rect 22661 4097 22695 4131
rect 25789 4097 25823 4131
rect 26801 4097 26835 4131
rect 27077 4097 27111 4131
rect 27997 4097 28031 4131
rect 28181 4097 28215 4131
rect 30849 4097 30883 4131
rect 31033 4097 31067 4131
rect 3433 4029 3467 4063
rect 3617 4029 3651 4063
rect 3709 4029 3743 4063
rect 5365 4029 5399 4063
rect 6837 4029 6871 4063
rect 8953 4029 8987 4063
rect 11253 4029 11287 4063
rect 13185 4029 13219 4063
rect 13277 4029 13311 4063
rect 13553 4029 13587 4063
rect 13820 4029 13854 4063
rect 16497 4029 16531 4063
rect 18337 4029 18371 4063
rect 18429 4029 18463 4063
rect 18705 4029 18739 4063
rect 21189 4029 21223 4063
rect 21372 4029 21406 4063
rect 21557 4029 21591 4063
rect 21741 4029 21775 4063
rect 22201 4029 22235 4063
rect 22293 4029 22327 4063
rect 23489 4029 23523 4063
rect 23581 4029 23615 4063
rect 23857 4029 23891 4063
rect 24113 4029 24147 4063
rect 26960 4029 26994 4063
rect 27813 4029 27847 4063
rect 30582 4029 30616 4063
rect 30941 4029 30975 4063
rect 3065 3961 3099 3995
rect 3249 3961 3283 3995
rect 3976 3961 4010 3995
rect 5632 3961 5666 3995
rect 7104 3961 7138 3995
rect 18950 3961 18984 3995
rect 29377 3961 29411 3995
rect 2865 3893 2899 3927
rect 8401 3893 8435 3927
rect 8585 3893 8619 3927
rect 11161 3893 11195 3927
rect 17785 3893 17819 3927
rect 17969 3893 18003 3927
rect 21833 3893 21867 3927
rect 25237 3893 25271 3927
rect 25329 3893 25363 3927
rect 28825 3893 28859 3927
rect 29177 3893 29211 3927
rect 3341 3689 3375 3723
rect 3801 3689 3835 3723
rect 3985 3689 4019 3723
rect 5549 3689 5583 3723
rect 5825 3689 5859 3723
rect 8217 3689 8251 3723
rect 12357 3689 12391 3723
rect 27537 3689 27571 3723
rect 29009 3689 29043 3723
rect 8401 3621 8435 3655
rect 8677 3621 8711 3655
rect 9965 3621 9999 3655
rect 10793 3621 10827 3655
rect 11222 3621 11256 3655
rect 21005 3621 21039 3655
rect 28650 3621 28684 3655
rect 3341 3553 3375 3587
rect 3525 3553 3559 3587
rect 3893 3553 3927 3587
rect 4261 3553 4295 3587
rect 4353 3553 4387 3587
rect 4445 3553 4479 3587
rect 4629 3553 4663 3587
rect 4721 3553 4755 3587
rect 4905 3553 4939 3587
rect 5641 3553 5675 3587
rect 6101 3553 6135 3587
rect 6193 3553 6227 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 7113 3553 7147 3587
rect 7573 3553 7607 3587
rect 7665 3553 7699 3587
rect 7757 3553 7791 3587
rect 7941 3553 7975 3587
rect 8033 3553 8067 3587
rect 8217 3553 8251 3587
rect 8309 3553 8343 3587
rect 8493 3553 8527 3587
rect 8585 3553 8619 3587
rect 8769 3553 8803 3587
rect 9873 3553 9907 3587
rect 10149 3553 10183 3587
rect 10333 3553 10367 3587
rect 10425 3553 10459 3587
rect 10517 3553 10551 3587
rect 10977 3553 11011 3587
rect 16497 3553 16531 3587
rect 19993 3553 20027 3587
rect 20453 3553 20487 3587
rect 20821 3553 20855 3587
rect 28917 3553 28951 3587
rect 29193 3553 29227 3587
rect 29285 3553 29319 3587
rect 4813 3485 4847 3519
rect 6561 3485 6595 3519
rect 20729 3485 20763 3519
rect 21281 3485 21315 3519
rect 21925 3485 21959 3519
rect 29009 3485 29043 3519
rect 7297 3349 7331 3383
rect 16405 3349 16439 3383
rect 19901 3349 19935 3383
rect 20269 3349 20303 3383
rect 20637 3349 20671 3383
rect 6653 3145 6687 3179
rect 8217 3145 8251 3179
rect 10609 3145 10643 3179
rect 11253 3145 11287 3179
rect 22845 3145 22879 3179
rect 24409 3145 24443 3179
rect 27077 3145 27111 3179
rect 27445 3145 27479 3179
rect 11805 3077 11839 3111
rect 16221 3077 16255 3111
rect 20913 3077 20947 3111
rect 21649 3077 21683 3111
rect 25605 3077 25639 3111
rect 6377 3009 6411 3043
rect 6837 3009 6871 3043
rect 11161 3009 11195 3043
rect 15853 3009 15887 3043
rect 21925 3009 21959 3043
rect 22201 3009 22235 3043
rect 25053 3009 25087 3043
rect 26065 3009 26099 3043
rect 26525 3009 26559 3043
rect 27353 3009 27387 3043
rect 28273 3009 28307 3043
rect 28457 3009 28491 3043
rect 6285 2941 6319 2975
rect 6561 2941 6595 2975
rect 7104 2941 7138 2975
rect 10149 2941 10183 2975
rect 10241 2941 10275 2975
rect 10333 2941 10367 2975
rect 10793 2941 10827 2975
rect 11529 2941 11563 2975
rect 13645 2941 13679 2975
rect 14197 2941 14231 2975
rect 16037 2941 16071 2975
rect 16129 2941 16163 2975
rect 16497 2941 16531 2975
rect 16865 2941 16899 2975
rect 17141 2941 17175 2975
rect 17325 2941 17359 2975
rect 19257 2941 19291 2975
rect 19349 2941 19383 2975
rect 19533 2941 19567 2975
rect 19800 2941 19834 2975
rect 21005 2941 21039 2975
rect 21189 2941 21223 2975
rect 22042 2941 22076 2975
rect 24041 2941 24075 2975
rect 25212 2941 25246 2975
rect 25329 2941 25363 2975
rect 26249 2941 26283 2975
rect 26709 2941 26743 2975
rect 26801 2941 26835 2975
rect 27537 2941 27571 2975
rect 27629 2941 27663 2975
rect 27721 2941 27755 2975
rect 28641 2941 28675 2975
rect 28825 2941 28859 2975
rect 29009 2941 29043 2975
rect 29193 2941 29227 2975
rect 29469 2941 29503 2975
rect 9965 2873 9999 2907
rect 15853 2873 15887 2907
rect 16221 2873 16255 2907
rect 16681 2873 16715 2907
rect 27261 2873 27295 2907
rect 10517 2805 10551 2839
rect 10885 2805 10919 2839
rect 10977 2805 11011 2839
rect 11437 2805 11471 2839
rect 11621 2805 11655 2839
rect 13829 2805 13863 2839
rect 14105 2805 14139 2839
rect 16405 2805 16439 2839
rect 17049 2805 17083 2839
rect 17509 2805 17543 2839
rect 23949 2805 23983 2839
rect 26525 2805 26559 2839
rect 26893 2805 26927 2839
rect 27061 2805 27095 2839
rect 29101 2805 29135 2839
rect 29377 2805 29411 2839
rect 15209 2601 15243 2635
rect 17693 2601 17727 2635
rect 10793 2533 10827 2567
rect 11145 2533 11179 2567
rect 11345 2533 11379 2567
rect 13093 2533 13127 2567
rect 15761 2533 15795 2567
rect 15945 2533 15979 2567
rect 26617 2533 26651 2567
rect 28488 2533 28522 2567
rect 10563 2499 10597 2533
rect 9597 2465 9631 2499
rect 9873 2465 9907 2499
rect 10149 2465 10183 2499
rect 11989 2465 12023 2499
rect 12449 2465 12483 2499
rect 13369 2465 13403 2499
rect 13625 2465 13659 2499
rect 15025 2465 15059 2499
rect 15301 2465 15335 2499
rect 16221 2465 16255 2499
rect 16477 2465 16511 2499
rect 18245 2465 18279 2499
rect 19717 2465 19751 2499
rect 19984 2465 20018 2499
rect 21557 2465 21591 2499
rect 21649 2465 21683 2499
rect 21925 2465 21959 2499
rect 22569 2465 22603 2499
rect 23765 2465 23799 2499
rect 24021 2465 24055 2499
rect 25513 2465 25547 2499
rect 25605 2465 25639 2499
rect 27169 2465 27203 2499
rect 28733 2465 28767 2499
rect 9965 2397 9999 2431
rect 11805 2397 11839 2431
rect 12173 2397 12207 2431
rect 12725 2397 12759 2431
rect 21465 2397 21499 2431
rect 21741 2397 21775 2431
rect 22293 2397 22327 2431
rect 25421 2397 25455 2431
rect 25697 2397 25731 2431
rect 10333 2329 10367 2363
rect 10977 2329 11011 2363
rect 12357 2329 12391 2363
rect 13277 2329 13311 2363
rect 14841 2329 14875 2363
rect 21097 2329 21131 2363
rect 25145 2329 25179 2363
rect 27353 2329 27387 2363
rect 9505 2261 9539 2295
rect 9781 2261 9815 2295
rect 10425 2261 10459 2295
rect 10609 2261 10643 2295
rect 11161 2261 11195 2295
rect 13093 2261 13127 2295
rect 14749 2261 14783 2295
rect 15577 2261 15611 2295
rect 17601 2261 17635 2295
rect 21281 2261 21315 2295
rect 22017 2261 22051 2295
rect 22385 2261 22419 2295
rect 22477 2261 22511 2295
rect 25237 2261 25271 2295
rect 11805 2057 11839 2091
rect 12449 2057 12483 2091
rect 12909 2057 12943 2091
rect 15025 2057 15059 2091
rect 15761 2057 15795 2091
rect 15945 2057 15979 2091
rect 17785 2057 17819 2091
rect 19993 2057 20027 2091
rect 20177 2057 20211 2091
rect 21557 2057 21591 2091
rect 22661 2057 22695 2091
rect 24041 2057 24075 2091
rect 25237 2057 25271 2091
rect 25421 2057 25455 2091
rect 26709 2057 26743 2091
rect 27077 2057 27111 2091
rect 10793 1989 10827 2023
rect 11621 1989 11655 2023
rect 12541 1989 12575 2023
rect 15209 1989 15243 2023
rect 15393 1989 15427 2023
rect 17417 1989 17451 2023
rect 18153 1989 18187 2023
rect 19901 1989 19935 2023
rect 20545 1989 20579 2023
rect 21373 1989 21407 2023
rect 21833 1989 21867 2023
rect 22385 1989 22419 2023
rect 22477 1989 22511 2023
rect 23673 1989 23707 2023
rect 23857 1989 23891 2023
rect 24501 1989 24535 2023
rect 26249 1989 26283 2023
rect 9229 1921 9263 1955
rect 9413 1921 9447 1955
rect 13553 1921 13587 1955
rect 22569 1921 22603 1955
rect 26433 1921 26467 1955
rect 26525 1921 26559 1955
rect 9321 1853 9355 1887
rect 11161 1853 11195 1887
rect 11253 1853 11287 1887
rect 11345 1853 11379 1887
rect 11529 1853 11563 1887
rect 12081 1853 12115 1887
rect 12265 1853 12299 1887
rect 13185 1853 13219 1887
rect 13829 1853 13863 1887
rect 16037 1853 16071 1887
rect 16304 1853 16338 1887
rect 18429 1853 18463 1887
rect 19349 1853 19383 1887
rect 19625 1853 19659 1887
rect 21189 1853 21223 1887
rect 22017 1855 22051 1889
rect 22109 1853 22143 1887
rect 22293 1853 22327 1887
rect 23213 1853 23247 1887
rect 23397 1853 23431 1887
rect 23673 1853 23707 1887
rect 24409 1853 24443 1887
rect 25145 1853 25179 1887
rect 25789 1853 25823 1887
rect 25881 1853 25915 1887
rect 26157 1853 26191 1887
rect 26801 1853 26835 1887
rect 28457 1853 28491 1887
rect 9680 1785 9714 1819
rect 10885 1785 10919 1819
rect 11989 1785 12023 1819
rect 12909 1785 12943 1819
rect 14841 1785 14875 1819
rect 15041 1785 15075 1819
rect 19901 1785 19935 1819
rect 20177 1785 20211 1819
rect 21525 1785 21559 1819
rect 21741 1785 21775 1819
rect 23489 1785 23523 1819
rect 24041 1785 24075 1819
rect 25605 1785 25639 1819
rect 26433 1785 26467 1819
rect 28190 1785 28224 1819
rect 11779 1717 11813 1751
rect 13093 1717 13127 1751
rect 13277 1717 13311 1751
rect 15761 1717 15795 1751
rect 17601 1717 17635 1751
rect 17785 1717 17819 1751
rect 18337 1717 18371 1751
rect 19441 1717 19475 1751
rect 19717 1717 19751 1751
rect 20637 1717 20671 1751
rect 25395 1717 25429 1751
rect 26065 1717 26099 1751
rect 26525 1717 26559 1751
rect 10701 1513 10735 1547
rect 11529 1513 11563 1547
rect 11713 1513 11747 1547
rect 13277 1513 13311 1547
rect 16221 1513 16255 1547
rect 16497 1513 16531 1547
rect 21097 1513 21131 1547
rect 22661 1513 22695 1547
rect 25329 1513 25363 1547
rect 27077 1513 27111 1547
rect 27537 1513 27571 1547
rect 12142 1445 12176 1479
rect 13614 1445 13648 1479
rect 17610 1445 17644 1479
rect 19962 1445 19996 1479
rect 24216 1445 24250 1479
rect 9321 1377 9355 1411
rect 9588 1377 9622 1411
rect 11161 1377 11195 1411
rect 11897 1377 11931 1411
rect 13369 1377 13403 1411
rect 16313 1377 16347 1411
rect 19717 1377 19751 1411
rect 21281 1377 21315 1411
rect 21548 1377 21582 1411
rect 23305 1377 23339 1411
rect 25421 1377 25455 1411
rect 25605 1377 25639 1411
rect 27169 1377 27203 1411
rect 27353 1377 27387 1411
rect 27445 1377 27479 1411
rect 17877 1309 17911 1343
rect 23213 1309 23247 1343
rect 23949 1309 23983 1343
rect 26433 1309 26467 1343
rect 27353 1241 27387 1275
rect 11529 1173 11563 1207
rect 14749 1173 14783 1207
rect 25605 1173 25639 1207
rect 10517 969 10551 1003
rect 11345 969 11379 1003
rect 21005 969 21039 1003
rect 25697 969 25731 1003
rect 10241 901 10275 935
rect 10425 833 10459 867
rect 10149 765 10183 799
rect 10517 765 10551 799
rect 10701 765 10735 799
rect 10977 765 11011 799
rect 11161 765 11195 799
rect 20821 765 20855 799
rect 21005 765 21039 799
rect 24041 765 24075 799
rect 24133 765 24167 799
rect 24317 765 24351 799
rect 24584 765 24618 799
rect 10425 697 10459 731
<< metal1 >>
rect 552 21786 31648 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 11436 21786
rect 11488 21734 11500 21786
rect 11552 21734 11564 21786
rect 11616 21734 11628 21786
rect 11680 21734 11692 21786
rect 11744 21734 19210 21786
rect 19262 21734 19274 21786
rect 19326 21734 19338 21786
rect 19390 21734 19402 21786
rect 19454 21734 19466 21786
rect 19518 21734 26984 21786
rect 27036 21734 27048 21786
rect 27100 21734 27112 21786
rect 27164 21734 27176 21786
rect 27228 21734 27240 21786
rect 27292 21734 31648 21786
rect 552 21712 31648 21734
rect 6454 21632 6460 21684
rect 6512 21632 6518 21684
rect 7282 21632 7288 21684
rect 7340 21632 7346 21684
rect 8386 21632 8392 21684
rect 8444 21632 8450 21684
rect 8662 21632 8668 21684
rect 8720 21632 8726 21684
rect 9401 21675 9459 21681
rect 9401 21641 9413 21675
rect 9447 21672 9459 21675
rect 9950 21672 9956 21684
rect 9447 21644 9956 21672
rect 9447 21641 9459 21644
rect 9401 21635 9459 21641
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 10318 21632 10324 21684
rect 10376 21632 10382 21684
rect 11790 21632 11796 21684
rect 11848 21632 11854 21684
rect 12250 21632 12256 21684
rect 12308 21632 12314 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 27522 21632 27528 21684
rect 27580 21672 27586 21684
rect 27580 21644 28028 21672
rect 27580 21632 27586 21644
rect 3326 21564 3332 21616
rect 3384 21604 3390 21616
rect 4062 21604 4068 21616
rect 3384 21576 4068 21604
rect 3384 21564 3390 21576
rect 4062 21564 4068 21576
rect 4120 21564 4126 21616
rect 25685 21607 25743 21613
rect 25685 21573 25697 21607
rect 25731 21604 25743 21607
rect 26878 21604 26884 21616
rect 25731 21576 26884 21604
rect 25731 21573 25743 21576
rect 25685 21567 25743 21573
rect 26878 21564 26884 21576
rect 26936 21564 26942 21616
rect 3068 21508 3464 21536
rect 2682 21428 2688 21480
rect 2740 21468 2746 21480
rect 3068 21477 3096 21508
rect 2777 21471 2835 21477
rect 2777 21468 2789 21471
rect 2740 21440 2789 21468
rect 2740 21428 2746 21440
rect 2777 21437 2789 21440
rect 2823 21468 2835 21471
rect 3053 21471 3111 21477
rect 3053 21468 3065 21471
rect 2823 21440 3065 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 3053 21437 3065 21440
rect 3099 21437 3111 21471
rect 3053 21431 3111 21437
rect 3234 21428 3240 21480
rect 3292 21428 3298 21480
rect 3326 21428 3332 21480
rect 3384 21428 3390 21480
rect 3436 21468 3464 21508
rect 3510 21496 3516 21548
rect 3568 21496 3574 21548
rect 8018 21536 8024 21548
rect 3988 21508 8024 21536
rect 3988 21477 4016 21508
rect 3973 21471 4031 21477
rect 3973 21468 3985 21471
rect 3436 21440 3985 21468
rect 3973 21437 3985 21440
rect 4019 21437 4031 21471
rect 3973 21431 4031 21437
rect 4062 21428 4068 21480
rect 4120 21428 4126 21480
rect 4246 21428 4252 21480
rect 4304 21428 4310 21480
rect 6104 21477 6132 21508
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 26510 21536 26516 21548
rect 11195 21508 11560 21536
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 6089 21471 6147 21477
rect 6089 21437 6101 21471
rect 6135 21437 6147 21471
rect 6089 21431 6147 21437
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 6641 21471 6699 21477
rect 6641 21468 6653 21471
rect 6512 21440 6653 21468
rect 6512 21428 6518 21440
rect 6641 21437 6653 21440
rect 6687 21468 6699 21471
rect 8205 21471 8263 21477
rect 8205 21468 8217 21471
rect 6687 21440 8217 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 8205 21437 8217 21440
rect 8251 21468 8263 21471
rect 8294 21468 8300 21480
rect 8251 21440 8300 21468
rect 8251 21437 8263 21440
rect 8205 21431 8263 21437
rect 8294 21428 8300 21440
rect 8352 21468 8358 21480
rect 9217 21471 9275 21477
rect 9217 21468 9229 21471
rect 8352 21440 9229 21468
rect 8352 21428 8358 21440
rect 9217 21437 9229 21440
rect 9263 21437 9275 21471
rect 9217 21431 9275 21437
rect 9585 21471 9643 21477
rect 9585 21437 9597 21471
rect 9631 21437 9643 21471
rect 9585 21431 9643 21437
rect 9677 21471 9735 21477
rect 9677 21437 9689 21471
rect 9723 21437 9735 21471
rect 9677 21431 9735 21437
rect 2406 21360 2412 21412
rect 2464 21400 2470 21412
rect 2961 21403 3019 21409
rect 2961 21400 2973 21403
rect 2464 21372 2973 21400
rect 2464 21360 2470 21372
rect 2961 21369 2973 21372
rect 3007 21369 3019 21403
rect 2961 21363 3019 21369
rect 3418 21360 3424 21412
rect 3476 21400 3482 21412
rect 3881 21403 3939 21409
rect 3881 21400 3893 21403
rect 3476 21372 3893 21400
rect 3476 21360 3482 21372
rect 3881 21369 3893 21372
rect 3927 21369 3939 21403
rect 3881 21363 3939 21369
rect 6917 21403 6975 21409
rect 6917 21369 6929 21403
rect 6963 21369 6975 21403
rect 6917 21363 6975 21369
rect 7101 21403 7159 21409
rect 7101 21369 7113 21403
rect 7147 21400 7159 21403
rect 7561 21403 7619 21409
rect 7561 21400 7573 21403
rect 7147 21372 7573 21400
rect 7147 21369 7159 21372
rect 7101 21363 7159 21369
rect 7561 21369 7573 21372
rect 7607 21369 7619 21403
rect 7561 21363 7619 21369
rect 2498 21292 2504 21344
rect 2556 21332 2562 21344
rect 2685 21335 2743 21341
rect 2685 21332 2697 21335
rect 2556 21304 2697 21332
rect 2556 21292 2562 21304
rect 2685 21301 2697 21304
rect 2731 21301 2743 21335
rect 2685 21295 2743 21301
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 3513 21335 3571 21341
rect 3513 21332 3525 21335
rect 2832 21304 3525 21332
rect 2832 21292 2838 21304
rect 3513 21301 3525 21304
rect 3559 21301 3571 21335
rect 3513 21295 3571 21301
rect 4062 21292 4068 21344
rect 4120 21292 4126 21344
rect 6178 21292 6184 21344
rect 6236 21292 6242 21344
rect 6733 21335 6791 21341
rect 6733 21301 6745 21335
rect 6779 21332 6791 21335
rect 6822 21332 6828 21344
rect 6779 21304 6828 21332
rect 6779 21301 6791 21304
rect 6733 21295 6791 21301
rect 6822 21292 6828 21304
rect 6880 21292 6886 21344
rect 6932 21332 6960 21363
rect 7006 21332 7012 21344
rect 6932 21304 7012 21332
rect 7006 21292 7012 21304
rect 7064 21332 7070 21344
rect 9600 21332 9628 21431
rect 7064 21304 9628 21332
rect 9692 21332 9720 21431
rect 9858 21428 9864 21480
rect 9916 21428 9922 21480
rect 9953 21471 10011 21477
rect 9953 21437 9965 21471
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 9766 21360 9772 21412
rect 9824 21400 9830 21412
rect 9968 21400 9996 21431
rect 10502 21428 10508 21480
rect 10560 21428 10566 21480
rect 11241 21471 11299 21477
rect 11241 21437 11253 21471
rect 11287 21437 11299 21471
rect 11241 21431 11299 21437
rect 9824 21372 9996 21400
rect 11256 21400 11284 21431
rect 11330 21428 11336 21480
rect 11388 21428 11394 21480
rect 11532 21477 11560 21508
rect 12406 21508 13768 21536
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 12406 21400 12434 21508
rect 13740 21480 13768 21508
rect 15672 21508 16988 21536
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 15672 21477 15700 21508
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 13780 21440 15669 21468
rect 13780 21428 13786 21440
rect 15657 21437 15669 21440
rect 15703 21437 15715 21471
rect 15657 21431 15715 21437
rect 16393 21471 16451 21477
rect 16393 21437 16405 21471
rect 16439 21468 16451 21471
rect 16574 21468 16580 21480
rect 16439 21440 16580 21468
rect 16439 21437 16451 21440
rect 16393 21431 16451 21437
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 16666 21428 16672 21480
rect 16724 21428 16730 21480
rect 16960 21477 16988 21508
rect 25792 21508 26516 21536
rect 16945 21471 17003 21477
rect 16945 21437 16957 21471
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 18598 21428 18604 21480
rect 18656 21468 18662 21480
rect 19153 21471 19211 21477
rect 19153 21468 19165 21471
rect 18656 21440 19165 21468
rect 18656 21428 18662 21440
rect 19153 21437 19165 21440
rect 19199 21437 19211 21471
rect 19153 21431 19211 21437
rect 19426 21428 19432 21480
rect 19484 21468 19490 21480
rect 19521 21471 19579 21477
rect 19521 21468 19533 21471
rect 19484 21440 19533 21468
rect 19484 21428 19490 21440
rect 19521 21437 19533 21440
rect 19567 21437 19579 21471
rect 19521 21431 19579 21437
rect 11256 21372 12434 21400
rect 16853 21403 16911 21409
rect 9824 21360 9830 21372
rect 16853 21369 16865 21403
rect 16899 21400 16911 21403
rect 17586 21400 17592 21412
rect 16899 21372 17592 21400
rect 16899 21369 16911 21372
rect 16853 21363 16911 21369
rect 17586 21360 17592 21372
rect 17644 21360 17650 21412
rect 19242 21360 19248 21412
rect 19300 21360 19306 21412
rect 19337 21403 19395 21409
rect 19337 21369 19349 21403
rect 19383 21369 19395 21403
rect 19536 21400 19564 21431
rect 19794 21428 19800 21480
rect 19852 21468 19858 21480
rect 21542 21468 21548 21480
rect 19852 21440 21548 21468
rect 19852 21428 19858 21440
rect 21542 21428 21548 21440
rect 21600 21428 21606 21480
rect 21634 21428 21640 21480
rect 21692 21428 21698 21480
rect 23842 21428 23848 21480
rect 23900 21428 23906 21480
rect 24394 21428 24400 21480
rect 24452 21428 24458 21480
rect 24946 21428 24952 21480
rect 25004 21428 25010 21480
rect 25498 21428 25504 21480
rect 25556 21428 25562 21480
rect 25792 21477 25820 21508
rect 26510 21496 26516 21508
rect 26568 21496 26574 21548
rect 25777 21471 25835 21477
rect 25777 21437 25789 21471
rect 25823 21437 25835 21471
rect 25777 21431 25835 21437
rect 26050 21428 26056 21480
rect 26108 21428 26114 21480
rect 28000 21477 28028 21644
rect 28994 21496 29000 21548
rect 29052 21496 29058 21548
rect 27893 21471 27951 21477
rect 27893 21437 27905 21471
rect 27939 21437 27951 21471
rect 27893 21431 27951 21437
rect 27985 21471 28043 21477
rect 27985 21437 27997 21471
rect 28031 21437 28043 21471
rect 27985 21431 28043 21437
rect 20254 21400 20260 21412
rect 19536 21372 20260 21400
rect 19337 21363 19395 21369
rect 9950 21332 9956 21344
rect 9692 21304 9956 21332
rect 7064 21292 7070 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10134 21292 10140 21344
rect 10192 21292 10198 21344
rect 11609 21335 11667 21341
rect 11609 21301 11621 21335
rect 11655 21332 11667 21335
rect 12802 21332 12808 21344
rect 11655 21304 12808 21332
rect 11655 21301 11667 21304
rect 11609 21295 11667 21301
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 15562 21292 15568 21344
rect 15620 21292 15626 21344
rect 15746 21292 15752 21344
rect 15804 21332 15810 21344
rect 16485 21335 16543 21341
rect 16485 21332 16497 21335
rect 15804 21304 16497 21332
rect 15804 21292 15810 21304
rect 16485 21301 16497 21304
rect 16531 21332 16543 21335
rect 16758 21332 16764 21344
rect 16531 21304 16764 21332
rect 16531 21301 16543 21304
rect 16485 21295 16543 21301
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 17770 21332 17776 21344
rect 17083 21304 17776 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 17770 21292 17776 21304
rect 17828 21292 17834 21344
rect 18506 21292 18512 21344
rect 18564 21332 18570 21344
rect 18969 21335 19027 21341
rect 18969 21332 18981 21335
rect 18564 21304 18981 21332
rect 18564 21292 18570 21304
rect 18969 21301 18981 21304
rect 19015 21301 19027 21335
rect 19352 21332 19380 21363
rect 20254 21360 20260 21372
rect 20312 21360 20318 21412
rect 27626 21403 27684 21409
rect 27626 21400 27638 21403
rect 25976 21372 27638 21400
rect 19610 21332 19616 21344
rect 19352 21304 19616 21332
rect 18969 21295 19027 21301
rect 19610 21292 19616 21304
rect 19668 21292 19674 21344
rect 19702 21292 19708 21344
rect 19760 21292 19766 21344
rect 21818 21292 21824 21344
rect 21876 21292 21882 21344
rect 24026 21292 24032 21344
rect 24084 21292 24090 21344
rect 24578 21292 24584 21344
rect 24636 21292 24642 21344
rect 25130 21292 25136 21344
rect 25188 21292 25194 21344
rect 25976 21341 26004 21372
rect 27626 21369 27638 21372
rect 27672 21369 27684 21403
rect 27908 21400 27936 21431
rect 28258 21428 28264 21480
rect 28316 21428 28322 21480
rect 29178 21428 29184 21480
rect 29236 21468 29242 21480
rect 29273 21471 29331 21477
rect 29273 21468 29285 21471
rect 29236 21440 29285 21468
rect 29236 21428 29242 21440
rect 29273 21437 29285 21440
rect 29319 21437 29331 21471
rect 29273 21431 29331 21437
rect 27908 21372 28028 21400
rect 27626 21363 27684 21369
rect 28000 21344 28028 21372
rect 25961 21335 26019 21341
rect 25961 21301 25973 21335
rect 26007 21301 26019 21335
rect 25961 21295 26019 21301
rect 26234 21292 26240 21344
rect 26292 21292 26298 21344
rect 26510 21292 26516 21344
rect 26568 21292 26574 21344
rect 27982 21292 27988 21344
rect 28040 21292 28046 21344
rect 28166 21292 28172 21344
rect 28224 21292 28230 21344
rect 28445 21335 28503 21341
rect 28445 21301 28457 21335
rect 28491 21332 28503 21335
rect 30466 21332 30472 21344
rect 28491 21304 30472 21332
rect 28491 21301 28503 21304
rect 28445 21295 28503 21301
rect 30466 21292 30472 21304
rect 30524 21292 30530 21344
rect 552 21242 31648 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 12096 21242
rect 12148 21190 12160 21242
rect 12212 21190 12224 21242
rect 12276 21190 12288 21242
rect 12340 21190 12352 21242
rect 12404 21190 19870 21242
rect 19922 21190 19934 21242
rect 19986 21190 19998 21242
rect 20050 21190 20062 21242
rect 20114 21190 20126 21242
rect 20178 21190 27644 21242
rect 27696 21190 27708 21242
rect 27760 21190 27772 21242
rect 27824 21190 27836 21242
rect 27888 21190 27900 21242
rect 27952 21190 31648 21242
rect 552 21168 31648 21190
rect 1029 21131 1087 21137
rect 1029 21097 1041 21131
rect 1075 21128 1087 21131
rect 3234 21128 3240 21140
rect 1075 21100 3240 21128
rect 1075 21097 1087 21100
rect 1029 21091 1087 21097
rect 3234 21088 3240 21100
rect 3292 21088 3298 21140
rect 3970 21088 3976 21140
rect 4028 21128 4034 21140
rect 4249 21131 4307 21137
rect 4249 21128 4261 21131
rect 4028 21100 4261 21128
rect 4028 21088 4034 21100
rect 4249 21097 4261 21100
rect 4295 21097 4307 21131
rect 4249 21091 4307 21097
rect 6270 21088 6276 21140
rect 6328 21088 6334 21140
rect 7929 21131 7987 21137
rect 7929 21097 7941 21131
rect 7975 21128 7987 21131
rect 8294 21128 8300 21140
rect 7975 21100 8300 21128
rect 7975 21097 7987 21100
rect 7929 21091 7987 21097
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 8478 21088 8484 21140
rect 8536 21088 8542 21140
rect 9858 21088 9864 21140
rect 9916 21128 9922 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 9916 21100 10149 21128
rect 9916 21088 9922 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 12621 21131 12679 21137
rect 12621 21097 12633 21131
rect 12667 21128 12679 21131
rect 13814 21128 13820 21140
rect 12667 21100 13820 21128
rect 12667 21097 12679 21100
rect 12621 21091 12679 21097
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 16393 21131 16451 21137
rect 16393 21097 16405 21131
rect 16439 21128 16451 21131
rect 16666 21128 16672 21140
rect 16439 21100 16672 21128
rect 16439 21097 16451 21100
rect 16393 21091 16451 21097
rect 16666 21088 16672 21100
rect 16724 21128 16730 21140
rect 16724 21100 18368 21128
rect 16724 21088 16730 21100
rect 3510 21020 3516 21072
rect 3568 21060 3574 21072
rect 5350 21060 5356 21072
rect 3568 21032 5356 21060
rect 3568 21020 3574 21032
rect 5350 21020 5356 21032
rect 5408 21060 5414 21072
rect 5408 21032 6132 21060
rect 5408 21020 5414 21032
rect 2153 20995 2211 21001
rect 2153 20961 2165 20995
rect 2199 20992 2211 20995
rect 2314 20992 2320 21004
rect 2199 20964 2320 20992
rect 2199 20961 2211 20964
rect 2153 20955 2211 20961
rect 2314 20952 2320 20964
rect 2372 20952 2378 21004
rect 2406 20952 2412 21004
rect 2464 20952 2470 21004
rect 2498 20952 2504 21004
rect 2556 20952 2562 21004
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 4062 20992 4068 21004
rect 2823 20964 4068 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 4157 20995 4215 21001
rect 4157 20961 4169 20995
rect 4203 20992 4215 20995
rect 4430 20992 4436 21004
rect 4203 20964 4436 20992
rect 4203 20961 4215 20964
rect 4157 20955 4215 20961
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 4614 20952 4620 21004
rect 4672 20952 4678 21004
rect 6104 21001 6132 21032
rect 6178 21020 6184 21072
rect 6236 21060 6242 21072
rect 6236 21032 6592 21060
rect 6236 21020 6242 21032
rect 5537 20995 5595 21001
rect 5537 20961 5549 20995
rect 5583 20961 5595 20995
rect 5537 20955 5595 20961
rect 6089 20995 6147 21001
rect 6089 20961 6101 20995
rect 6135 20961 6147 20995
rect 6089 20955 6147 20961
rect 5552 20856 5580 20955
rect 6454 20952 6460 21004
rect 6512 20952 6518 21004
rect 6564 21001 6592 21032
rect 11698 21020 11704 21072
rect 11756 21020 11762 21072
rect 17678 21020 17684 21072
rect 17736 21060 17742 21072
rect 18141 21063 18199 21069
rect 18141 21060 18153 21063
rect 17736 21032 18153 21060
rect 17736 21020 17742 21032
rect 18141 21029 18153 21032
rect 18187 21029 18199 21063
rect 18141 21023 18199 21029
rect 6822 21001 6828 21004
rect 6549 20995 6607 21001
rect 6549 20961 6561 20995
rect 6595 20961 6607 20995
rect 6816 20992 6828 21001
rect 6783 20964 6828 20992
rect 6549 20955 6607 20961
rect 6816 20955 6828 20964
rect 6822 20952 6828 20955
rect 6880 20952 6886 21004
rect 8294 20952 8300 21004
rect 8352 20952 8358 21004
rect 8386 20952 8392 21004
rect 8444 20992 8450 21004
rect 8849 20995 8907 21001
rect 8849 20992 8861 20995
rect 8444 20964 8861 20992
rect 8444 20952 8450 20964
rect 8849 20961 8861 20964
rect 8895 20961 8907 20995
rect 8849 20955 8907 20961
rect 9125 20995 9183 21001
rect 9125 20961 9137 20995
rect 9171 20961 9183 20995
rect 9125 20955 9183 20961
rect 9309 20995 9367 21001
rect 9309 20961 9321 20995
rect 9355 20992 9367 20995
rect 9401 20995 9459 21001
rect 9401 20992 9413 20995
rect 9355 20964 9413 20992
rect 9355 20961 9367 20964
rect 9309 20955 9367 20961
rect 9401 20961 9413 20964
rect 9447 20961 9459 20995
rect 9401 20955 9459 20961
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 10226 20992 10232 21004
rect 10091 20964 10232 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 8202 20884 8208 20936
rect 8260 20924 8266 20936
rect 9140 20924 9168 20955
rect 10226 20952 10232 20964
rect 10284 20992 10290 21004
rect 11241 20995 11299 21001
rect 11241 20992 11253 20995
rect 10284 20964 11253 20992
rect 10284 20952 10290 20964
rect 11241 20961 11253 20964
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 12066 20952 12072 21004
rect 12124 20952 12130 21004
rect 12345 20995 12403 21001
rect 12345 20961 12357 20995
rect 12391 20961 12403 20995
rect 12345 20955 12403 20961
rect 8260 20896 9168 20924
rect 8260 20884 8266 20896
rect 10318 20884 10324 20936
rect 10376 20924 10382 20936
rect 10689 20927 10747 20933
rect 10689 20924 10701 20927
rect 10376 20896 10701 20924
rect 10376 20884 10382 20896
rect 10689 20893 10701 20896
rect 10735 20924 10747 20927
rect 11330 20924 11336 20936
rect 10735 20896 11336 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 11330 20884 11336 20896
rect 11388 20924 11394 20936
rect 12360 20924 12388 20955
rect 12802 20952 12808 21004
rect 12860 20952 12866 21004
rect 13722 20952 13728 21004
rect 13780 20992 13786 21004
rect 13817 20995 13875 21001
rect 13817 20992 13829 20995
rect 13780 20964 13829 20992
rect 13780 20952 13786 20964
rect 13817 20961 13829 20964
rect 13863 20961 13875 20995
rect 13817 20955 13875 20961
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20961 15255 20995
rect 15197 20955 15255 20961
rect 11388 20896 12388 20924
rect 15212 20924 15240 20955
rect 15286 20952 15292 21004
rect 15344 20952 15350 21004
rect 15470 20952 15476 21004
rect 15528 20952 15534 21004
rect 15746 20952 15752 21004
rect 15804 20952 15810 21004
rect 15933 20995 15991 21001
rect 15933 20961 15945 20995
rect 15979 20992 15991 20995
rect 16574 20992 16580 21004
rect 15979 20964 16580 20992
rect 15979 20961 15991 20964
rect 15933 20955 15991 20961
rect 16574 20952 16580 20964
rect 16632 20952 16638 21004
rect 17770 20952 17776 21004
rect 17828 20952 17834 21004
rect 17954 20952 17960 21004
rect 18012 21001 18018 21004
rect 18012 20995 18061 21001
rect 18012 20961 18015 20995
rect 18049 20961 18061 20995
rect 18012 20955 18061 20961
rect 18012 20952 18018 20955
rect 18230 20952 18236 21004
rect 18288 20952 18294 21004
rect 18340 21001 18368 21100
rect 19242 21088 19248 21140
rect 19300 21128 19306 21140
rect 19886 21128 19892 21140
rect 19300 21100 19892 21128
rect 19300 21088 19306 21100
rect 19886 21088 19892 21100
rect 19944 21128 19950 21140
rect 20073 21131 20131 21137
rect 20073 21128 20085 21131
rect 19944 21100 20085 21128
rect 19944 21088 19950 21100
rect 20073 21097 20085 21100
rect 20119 21097 20131 21131
rect 20073 21091 20131 21097
rect 21542 21020 21548 21072
rect 21600 21060 21606 21072
rect 23876 21063 23934 21069
rect 21600 21032 22692 21060
rect 21600 21020 21606 21032
rect 18340 20995 18419 21001
rect 18340 20964 18373 20995
rect 18361 20961 18373 20964
rect 18407 20961 18419 20995
rect 18361 20955 18419 20961
rect 18506 20952 18512 21004
rect 18564 20952 18570 21004
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20992 18751 20995
rect 19702 20992 19708 21004
rect 18739 20964 19708 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 21818 20952 21824 21004
rect 21876 20992 21882 21004
rect 22664 21001 22692 21032
rect 23876 21029 23888 21063
rect 23922 21060 23934 21063
rect 24026 21060 24032 21072
rect 23922 21032 24032 21060
rect 23922 21029 23934 21032
rect 23876 21023 23934 21029
rect 24026 21020 24032 21032
rect 24084 21020 24090 21072
rect 24136 21032 25636 21060
rect 24136 21001 24164 21032
rect 22382 20995 22440 21001
rect 22382 20992 22394 20995
rect 21876 20964 22394 20992
rect 21876 20952 21882 20964
rect 22382 20961 22394 20964
rect 22428 20961 22440 20995
rect 22382 20955 22440 20961
rect 22649 20995 22707 21001
rect 22649 20961 22661 20995
rect 22695 20961 22707 20995
rect 22649 20955 22707 20961
rect 24121 20995 24179 21001
rect 24121 20961 24133 20995
rect 24167 20961 24179 20995
rect 24121 20955 24179 20961
rect 24578 20952 24584 21004
rect 24636 20992 24642 21004
rect 25326 20995 25384 21001
rect 25326 20992 25338 20995
rect 24636 20964 25338 20992
rect 24636 20952 24642 20964
rect 25326 20961 25338 20964
rect 25372 20961 25384 20995
rect 25326 20955 25384 20961
rect 15764 20924 15792 20952
rect 15212 20896 15792 20924
rect 11388 20884 11394 20896
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 18966 20884 18972 20936
rect 19024 20884 19030 20936
rect 25608 20933 25636 21032
rect 26234 21020 26240 21072
rect 26292 21060 26298 21072
rect 27534 21063 27592 21069
rect 27534 21060 27546 21063
rect 26292 21032 27546 21060
rect 26292 21020 26298 21032
rect 27534 21029 27546 21032
rect 27580 21029 27592 21063
rect 27534 21023 27592 21029
rect 28166 21020 28172 21072
rect 28224 21060 28230 21072
rect 29006 21063 29064 21069
rect 29006 21060 29018 21063
rect 28224 21032 29018 21060
rect 28224 21020 28230 21032
rect 29006 21029 29018 21032
rect 29052 21029 29064 21063
rect 29006 21023 29064 21029
rect 29288 21032 30788 21060
rect 29288 20936 29316 21032
rect 30466 20952 30472 21004
rect 30524 21001 30530 21004
rect 30760 21001 30788 21032
rect 30524 20992 30536 21001
rect 30745 20995 30803 21001
rect 30524 20964 30569 20992
rect 30524 20955 30536 20964
rect 30745 20961 30757 20995
rect 30791 20961 30803 20995
rect 30745 20955 30803 20961
rect 30524 20952 30530 20955
rect 25593 20927 25651 20933
rect 25593 20893 25605 20927
rect 25639 20924 25651 20927
rect 25774 20924 25780 20936
rect 25639 20896 25780 20924
rect 25639 20893 25651 20896
rect 25593 20887 25651 20893
rect 25774 20884 25780 20896
rect 25832 20884 25838 20936
rect 27798 20884 27804 20936
rect 27856 20884 27862 20936
rect 29270 20884 29276 20936
rect 29328 20884 29334 20936
rect 4172 20828 5580 20856
rect 11517 20859 11575 20865
rect 2222 20748 2228 20800
rect 2280 20788 2286 20800
rect 2682 20788 2688 20800
rect 2280 20760 2688 20788
rect 2280 20748 2286 20760
rect 2682 20748 2688 20760
rect 2740 20788 2746 20800
rect 4172 20788 4200 20828
rect 11517 20825 11529 20859
rect 11563 20856 11575 20859
rect 12894 20856 12900 20868
rect 11563 20828 12900 20856
rect 11563 20825 11575 20828
rect 11517 20819 11575 20825
rect 12894 20816 12900 20828
rect 12952 20816 12958 20868
rect 12989 20859 13047 20865
rect 12989 20825 13001 20859
rect 13035 20856 13047 20859
rect 13814 20856 13820 20868
rect 13035 20828 13820 20856
rect 13035 20825 13047 20828
rect 12989 20819 13047 20825
rect 13814 20816 13820 20828
rect 13872 20816 13878 20868
rect 2740 20760 4200 20788
rect 2740 20748 2746 20760
rect 5442 20748 5448 20800
rect 5500 20748 5506 20800
rect 5905 20791 5963 20797
rect 5905 20757 5917 20791
rect 5951 20788 5963 20791
rect 6270 20788 6276 20800
rect 5951 20760 6276 20788
rect 5951 20757 5963 20760
rect 5905 20751 5963 20757
rect 6270 20748 6276 20760
rect 6328 20748 6334 20800
rect 8662 20748 8668 20800
rect 8720 20748 8726 20800
rect 13722 20748 13728 20800
rect 13780 20748 13786 20800
rect 15657 20791 15715 20797
rect 15657 20757 15669 20791
rect 15703 20788 15715 20791
rect 15746 20788 15752 20800
rect 15703 20760 15752 20788
rect 15703 20757 15715 20760
rect 15657 20751 15715 20757
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 15838 20748 15844 20800
rect 15896 20748 15902 20800
rect 17862 20748 17868 20800
rect 17920 20748 17926 20800
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 21269 20791 21327 20797
rect 21269 20788 21281 20791
rect 20864 20760 21281 20788
rect 20864 20748 20870 20760
rect 21269 20757 21281 20760
rect 21315 20757 21327 20791
rect 21269 20751 21327 20757
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 22741 20791 22799 20797
rect 22741 20788 22753 20791
rect 22704 20760 22753 20788
rect 22704 20748 22710 20760
rect 22741 20757 22753 20760
rect 22787 20757 22799 20791
rect 22741 20751 22799 20757
rect 24210 20748 24216 20800
rect 24268 20748 24274 20800
rect 26418 20748 26424 20800
rect 26476 20748 26482 20800
rect 27893 20791 27951 20797
rect 27893 20757 27905 20791
rect 27939 20788 27951 20791
rect 28074 20788 28080 20800
rect 27939 20760 28080 20788
rect 27939 20757 27951 20760
rect 27893 20751 27951 20757
rect 28074 20748 28080 20760
rect 28132 20748 28138 20800
rect 29362 20748 29368 20800
rect 29420 20748 29426 20800
rect 552 20698 31648 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 11436 20698
rect 11488 20646 11500 20698
rect 11552 20646 11564 20698
rect 11616 20646 11628 20698
rect 11680 20646 11692 20698
rect 11744 20646 19210 20698
rect 19262 20646 19274 20698
rect 19326 20646 19338 20698
rect 19390 20646 19402 20698
rect 19454 20646 19466 20698
rect 19518 20646 26984 20698
rect 27036 20646 27048 20698
rect 27100 20646 27112 20698
rect 27164 20646 27176 20698
rect 27228 20646 27240 20698
rect 27292 20646 31648 20698
rect 552 20624 31648 20646
rect 2314 20544 2320 20596
rect 2372 20584 2378 20596
rect 2593 20587 2651 20593
rect 2593 20584 2605 20587
rect 2372 20556 2605 20584
rect 2372 20544 2378 20556
rect 2593 20553 2605 20556
rect 2639 20553 2651 20587
rect 2593 20547 2651 20553
rect 4246 20544 4252 20596
rect 4304 20584 4310 20596
rect 4341 20587 4399 20593
rect 4341 20584 4353 20587
rect 4304 20556 4353 20584
rect 4304 20544 4310 20556
rect 4341 20553 4353 20556
rect 4387 20553 4399 20587
rect 4341 20547 4399 20553
rect 8570 20544 8576 20596
rect 8628 20544 8634 20596
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 12066 20584 12072 20596
rect 12023 20556 12072 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 16942 20544 16948 20596
rect 17000 20544 17006 20596
rect 17129 20587 17187 20593
rect 17129 20553 17141 20587
rect 17175 20584 17187 20587
rect 17494 20584 17500 20596
rect 17175 20556 17500 20584
rect 17175 20553 17187 20556
rect 17129 20547 17187 20553
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 20254 20544 20260 20596
rect 20312 20544 20318 20596
rect 29362 20584 29368 20596
rect 21928 20556 29368 20584
rect 17865 20519 17923 20525
rect 17865 20485 17877 20519
rect 17911 20516 17923 20519
rect 18046 20516 18052 20528
rect 17911 20488 18052 20516
rect 17911 20485 17923 20488
rect 17865 20479 17923 20485
rect 18046 20476 18052 20488
rect 18104 20476 18110 20528
rect 18598 20516 18604 20528
rect 18156 20488 18604 20516
rect 4430 20408 4436 20460
rect 4488 20448 4494 20460
rect 5074 20448 5080 20460
rect 4488 20420 5080 20448
rect 4488 20408 4494 20420
rect 2222 20340 2228 20392
rect 2280 20340 2286 20392
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20380 3111 20383
rect 3326 20380 3332 20392
rect 3099 20352 3332 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 3326 20340 3332 20352
rect 3384 20340 3390 20392
rect 4062 20340 4068 20392
rect 4120 20340 4126 20392
rect 4540 20389 4568 20420
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 5261 20451 5319 20457
rect 5261 20417 5273 20451
rect 5307 20448 5319 20451
rect 5442 20448 5448 20460
rect 5307 20420 5448 20448
rect 5307 20417 5319 20420
rect 5261 20411 5319 20417
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 5994 20408 6000 20460
rect 6052 20448 6058 20460
rect 6641 20451 6699 20457
rect 6641 20448 6653 20451
rect 6052 20420 6653 20448
rect 6052 20408 6058 20420
rect 6641 20417 6653 20420
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20448 13599 20451
rect 13722 20448 13728 20460
rect 13587 20420 13728 20448
rect 13587 20417 13599 20420
rect 13541 20411 13599 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20448 15439 20451
rect 15562 20448 15568 20460
rect 15427 20420 15568 20448
rect 15427 20417 15439 20420
rect 15381 20411 15439 20417
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 18156 20448 18184 20488
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 18693 20451 18751 20457
rect 18693 20448 18705 20451
rect 15896 20420 17540 20448
rect 15896 20408 15902 20420
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20349 4583 20383
rect 4525 20343 4583 20349
rect 4614 20340 4620 20392
rect 4672 20340 4678 20392
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 4798 20380 4804 20392
rect 4755 20352 4804 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 4982 20340 4988 20392
rect 5040 20340 5046 20392
rect 5169 20383 5227 20389
rect 5169 20349 5181 20383
rect 5215 20380 5227 20383
rect 5537 20383 5595 20389
rect 5537 20380 5549 20383
rect 5215 20352 5549 20380
rect 5215 20349 5227 20352
rect 5169 20343 5227 20349
rect 5537 20349 5549 20352
rect 5583 20349 5595 20383
rect 5537 20343 5595 20349
rect 8018 20340 8024 20392
rect 8076 20340 8082 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 8389 20383 8447 20389
rect 8389 20380 8401 20383
rect 8352 20352 8401 20380
rect 8352 20340 8358 20352
rect 8389 20349 8401 20352
rect 8435 20349 8447 20383
rect 8389 20343 8447 20349
rect 8938 20340 8944 20392
rect 8996 20340 9002 20392
rect 9208 20383 9266 20389
rect 9208 20349 9220 20383
rect 9254 20380 9266 20383
rect 10134 20380 10140 20392
rect 9254 20352 10140 20380
rect 9254 20349 9266 20352
rect 9208 20343 9266 20349
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 10597 20383 10655 20389
rect 10597 20349 10609 20383
rect 10643 20380 10655 20383
rect 12161 20383 12219 20389
rect 12161 20380 12173 20383
rect 10643 20352 12173 20380
rect 10643 20349 10655 20352
rect 10597 20343 10655 20349
rect 12161 20349 12173 20352
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12618 20380 12624 20392
rect 12299 20352 12624 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12618 20340 12624 20352
rect 12676 20380 12682 20392
rect 13173 20383 13231 20389
rect 13173 20380 13185 20383
rect 12676 20352 13185 20380
rect 12676 20340 12682 20352
rect 13173 20349 13185 20352
rect 13219 20380 13231 20383
rect 13630 20380 13636 20392
rect 13219 20352 13636 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 13814 20340 13820 20392
rect 13872 20340 13878 20392
rect 15654 20340 15660 20392
rect 15712 20340 15718 20392
rect 16758 20340 16764 20392
rect 16816 20380 16822 20392
rect 17512 20389 17540 20420
rect 17696 20420 18184 20448
rect 17405 20383 17463 20389
rect 17405 20380 17417 20383
rect 16816 20352 17417 20380
rect 16816 20340 16822 20352
rect 17405 20349 17417 20352
rect 17451 20349 17463 20383
rect 17405 20343 17463 20349
rect 17497 20383 17555 20389
rect 17497 20349 17509 20383
rect 17543 20349 17555 20383
rect 17497 20343 17555 20349
rect 2961 20315 3019 20321
rect 2961 20281 2973 20315
rect 3007 20312 3019 20315
rect 3234 20312 3240 20324
rect 3007 20284 3240 20312
rect 3007 20281 3019 20284
rect 2961 20275 3019 20281
rect 3234 20272 3240 20284
rect 3292 20272 3298 20324
rect 4341 20315 4399 20321
rect 4341 20281 4353 20315
rect 4387 20312 4399 20315
rect 7006 20312 7012 20324
rect 4387 20284 5396 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 1946 20204 1952 20256
rect 2004 20244 2010 20256
rect 2133 20247 2191 20253
rect 2133 20244 2145 20247
rect 2004 20216 2145 20244
rect 2004 20204 2010 20216
rect 2133 20213 2145 20216
rect 2179 20213 2191 20247
rect 2133 20207 2191 20213
rect 3326 20204 3332 20256
rect 3384 20244 3390 20256
rect 3421 20247 3479 20253
rect 3421 20244 3433 20247
rect 3384 20216 3433 20244
rect 3384 20204 3390 20216
rect 3421 20213 3433 20216
rect 3467 20213 3479 20247
rect 3421 20207 3479 20213
rect 4801 20247 4859 20253
rect 4801 20213 4813 20247
rect 4847 20244 4859 20247
rect 4890 20244 4896 20256
rect 4847 20216 4896 20244
rect 4847 20213 4859 20216
rect 4801 20207 4859 20213
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 5368 20244 5396 20284
rect 6196 20284 7012 20312
rect 6196 20244 6224 20284
rect 7006 20272 7012 20284
rect 7064 20272 7070 20324
rect 10864 20315 10922 20321
rect 10864 20281 10876 20315
rect 10910 20312 10922 20315
rect 11054 20312 11060 20324
rect 10910 20284 11060 20312
rect 10910 20281 10922 20284
rect 10864 20275 10922 20281
rect 11054 20272 11060 20284
rect 11112 20272 11118 20324
rect 17420 20312 17448 20343
rect 17586 20340 17592 20392
rect 17644 20340 17650 20392
rect 17696 20312 17724 20420
rect 18156 20389 18184 20420
rect 18432 20420 18705 20448
rect 18432 20392 18460 20420
rect 18693 20417 18705 20420
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 20441 20451 20499 20457
rect 20441 20448 20453 20451
rect 18932 20420 20453 20448
rect 18932 20408 18938 20420
rect 20441 20417 20453 20420
rect 20487 20417 20499 20451
rect 20441 20411 20499 20417
rect 17773 20383 17831 20389
rect 17773 20349 17785 20383
rect 17819 20349 17831 20383
rect 17773 20343 17831 20349
rect 18141 20383 18199 20389
rect 18141 20349 18153 20383
rect 18187 20349 18199 20383
rect 18141 20343 18199 20349
rect 17420 20284 17724 20312
rect 17788 20256 17816 20343
rect 18230 20340 18236 20392
rect 18288 20340 18294 20392
rect 18322 20340 18328 20392
rect 18380 20340 18386 20392
rect 18414 20340 18420 20392
rect 18472 20340 18478 20392
rect 18509 20383 18567 20389
rect 18509 20349 18521 20383
rect 18555 20380 18567 20383
rect 18969 20383 19027 20389
rect 18616 20380 18828 20382
rect 18555 20354 18828 20380
rect 18555 20352 18644 20354
rect 18555 20349 18567 20352
rect 18509 20343 18567 20349
rect 5368 20216 6224 20244
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8478 20244 8484 20256
rect 8159 20216 8484 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 13265 20247 13323 20253
rect 13265 20213 13277 20247
rect 13311 20244 13323 20247
rect 13354 20244 13360 20256
rect 13311 20216 13360 20244
rect 13311 20213 13323 20216
rect 13265 20207 13323 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 15105 20247 15163 20253
rect 15105 20213 15117 20247
rect 15151 20244 15163 20247
rect 15194 20244 15200 20256
rect 15151 20216 15200 20244
rect 15151 20213 15163 20216
rect 15105 20207 15163 20213
rect 15194 20204 15200 20216
rect 15252 20244 15258 20256
rect 16022 20244 16028 20256
rect 15252 20216 16028 20244
rect 15252 20204 15258 20216
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 17034 20204 17040 20256
rect 17092 20244 17098 20256
rect 17770 20244 17776 20256
rect 17092 20216 17776 20244
rect 17092 20204 17098 20216
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 18800 20244 18828 20354
rect 18969 20349 18981 20383
rect 19015 20380 19027 20383
rect 19058 20380 19064 20392
rect 19015 20352 19064 20380
rect 19015 20349 19027 20352
rect 18969 20343 19027 20349
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 19426 20340 19432 20392
rect 19484 20380 19490 20392
rect 19794 20380 19800 20392
rect 19484 20352 19800 20380
rect 19484 20340 19490 20352
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 20254 20340 20260 20392
rect 20312 20380 20318 20392
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 20312 20352 20637 20380
rect 20312 20340 20318 20352
rect 20625 20349 20637 20352
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 20898 20340 20904 20392
rect 20956 20340 20962 20392
rect 21928 20389 21956 20556
rect 29362 20544 29368 20556
rect 29420 20544 29426 20596
rect 22462 20408 22468 20460
rect 22520 20448 22526 20460
rect 22738 20448 22744 20460
rect 22520 20420 22744 20448
rect 22520 20408 22526 20420
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 29089 20451 29147 20457
rect 29089 20417 29101 20451
rect 29135 20448 29147 20451
rect 29549 20451 29607 20457
rect 29549 20448 29561 20451
rect 29135 20420 29561 20448
rect 29135 20417 29147 20420
rect 29089 20411 29147 20417
rect 29549 20417 29561 20420
rect 29595 20417 29607 20451
rect 29549 20411 29607 20417
rect 21913 20383 21971 20389
rect 21913 20349 21925 20383
rect 21959 20349 21971 20383
rect 21913 20343 21971 20349
rect 22281 20383 22339 20389
rect 22281 20349 22293 20383
rect 22327 20380 22339 20383
rect 22370 20380 22376 20392
rect 22327 20352 22376 20380
rect 22327 20349 22339 20352
rect 22281 20343 22339 20349
rect 22370 20340 22376 20352
rect 22428 20340 22434 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20349 22707 20383
rect 22649 20343 22707 20349
rect 22833 20383 22891 20389
rect 22833 20349 22845 20383
rect 22879 20349 22891 20383
rect 22833 20343 22891 20349
rect 19702 20272 19708 20324
rect 19760 20312 19766 20324
rect 20809 20315 20867 20321
rect 20809 20312 20821 20315
rect 19760 20284 20821 20312
rect 19760 20272 19766 20284
rect 20809 20281 20821 20284
rect 20855 20312 20867 20315
rect 22094 20312 22100 20324
rect 20855 20284 22100 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 22094 20272 22100 20284
rect 22152 20272 22158 20324
rect 22186 20272 22192 20324
rect 22244 20272 22250 20324
rect 22572 20312 22600 20343
rect 22296 20284 22600 20312
rect 19334 20244 19340 20256
rect 18800 20216 19340 20244
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 19886 20244 19892 20256
rect 19668 20216 19892 20244
rect 19668 20204 19674 20216
rect 19886 20204 19892 20216
rect 19944 20204 19950 20256
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 22296 20244 22324 20284
rect 20312 20216 22324 20244
rect 20312 20204 20318 20216
rect 22462 20204 22468 20256
rect 22520 20204 22526 20256
rect 22664 20244 22692 20343
rect 22848 20312 22876 20343
rect 22922 20340 22928 20392
rect 22980 20380 22986 20392
rect 23750 20380 23756 20392
rect 22980 20352 23756 20380
rect 22980 20340 22986 20352
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 25510 20383 25568 20389
rect 25510 20380 25522 20383
rect 25188 20352 25522 20380
rect 25188 20340 25194 20352
rect 25510 20349 25522 20352
rect 25556 20349 25568 20383
rect 25510 20343 25568 20349
rect 25774 20340 25780 20392
rect 25832 20380 25838 20392
rect 27249 20383 27307 20389
rect 27249 20380 27261 20383
rect 25832 20352 27261 20380
rect 25832 20340 25838 20352
rect 27249 20349 27261 20352
rect 27295 20380 27307 20383
rect 27798 20380 27804 20392
rect 27295 20352 27804 20380
rect 27295 20349 27307 20352
rect 27249 20343 27307 20349
rect 27798 20340 27804 20352
rect 27856 20380 27862 20392
rect 28997 20383 29055 20389
rect 28997 20380 29009 20383
rect 27856 20352 29009 20380
rect 27856 20340 27862 20352
rect 28997 20349 29009 20352
rect 29043 20380 29055 20383
rect 29270 20380 29276 20392
rect 29043 20352 29276 20380
rect 29043 20349 29055 20352
rect 28997 20343 29055 20349
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 26510 20312 26516 20324
rect 22848 20284 26516 20312
rect 26510 20272 26516 20284
rect 26568 20272 26574 20324
rect 26878 20272 26884 20324
rect 26936 20312 26942 20324
rect 26982 20315 27040 20321
rect 26982 20312 26994 20315
rect 26936 20284 26994 20312
rect 26936 20272 26942 20284
rect 26982 20281 26994 20284
rect 27028 20281 27040 20315
rect 26982 20275 27040 20281
rect 29454 20272 29460 20324
rect 29512 20312 29518 20324
rect 29794 20315 29852 20321
rect 29794 20312 29806 20315
rect 29512 20284 29806 20312
rect 29512 20272 29518 20284
rect 29794 20281 29806 20284
rect 29840 20281 29852 20315
rect 29794 20275 29852 20281
rect 22922 20244 22928 20256
rect 22664 20216 22928 20244
rect 22922 20204 22928 20216
rect 22980 20204 22986 20256
rect 23109 20247 23167 20253
rect 23109 20213 23121 20247
rect 23155 20244 23167 20247
rect 23474 20244 23480 20256
rect 23155 20216 23480 20244
rect 23155 20213 23167 20216
rect 23109 20207 23167 20213
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 24118 20204 24124 20256
rect 24176 20244 24182 20256
rect 24397 20247 24455 20253
rect 24397 20244 24409 20247
rect 24176 20216 24409 20244
rect 24176 20204 24182 20216
rect 24397 20213 24409 20216
rect 24443 20213 24455 20247
rect 24397 20207 24455 20213
rect 25866 20204 25872 20256
rect 25924 20204 25930 20256
rect 29365 20247 29423 20253
rect 29365 20213 29377 20247
rect 29411 20244 29423 20247
rect 29546 20244 29552 20256
rect 29411 20216 29552 20244
rect 29411 20213 29423 20216
rect 29365 20207 29423 20213
rect 29546 20204 29552 20216
rect 29604 20204 29610 20256
rect 29638 20204 29644 20256
rect 29696 20244 29702 20256
rect 30929 20247 30987 20253
rect 30929 20244 30941 20247
rect 29696 20216 30941 20244
rect 29696 20204 29702 20216
rect 30929 20213 30941 20216
rect 30975 20213 30987 20247
rect 30929 20207 30987 20213
rect 552 20154 31648 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 12096 20154
rect 12148 20102 12160 20154
rect 12212 20102 12224 20154
rect 12276 20102 12288 20154
rect 12340 20102 12352 20154
rect 12404 20102 19870 20154
rect 19922 20102 19934 20154
rect 19986 20102 19998 20154
rect 20050 20102 20062 20154
rect 20114 20102 20126 20154
rect 20178 20102 27644 20154
rect 27696 20102 27708 20154
rect 27760 20102 27772 20154
rect 27824 20102 27836 20154
rect 27888 20102 27900 20154
rect 27952 20102 31648 20154
rect 552 20080 31648 20102
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 5261 20043 5319 20049
rect 5261 20040 5273 20043
rect 5040 20012 5273 20040
rect 5040 20000 5046 20012
rect 5261 20009 5273 20012
rect 5307 20009 5319 20043
rect 5261 20003 5319 20009
rect 5350 20000 5356 20052
rect 5408 20040 5414 20052
rect 7098 20040 7104 20052
rect 5408 20012 7104 20040
rect 5408 20000 5414 20012
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20040 7619 20043
rect 8386 20040 8392 20052
rect 7607 20012 8392 20040
rect 7607 20009 7619 20012
rect 7561 20003 7619 20009
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 8481 20043 8539 20049
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 8938 20040 8944 20052
rect 8527 20012 8944 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 10226 20040 10232 20052
rect 10183 20012 10232 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 10226 20000 10232 20012
rect 10284 20000 10290 20052
rect 11054 20000 11060 20052
rect 11112 20000 11118 20052
rect 14734 20000 14740 20052
rect 14792 20040 14798 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 14792 20012 14933 20040
rect 14792 20000 14798 20012
rect 14921 20009 14933 20012
rect 14967 20040 14979 20043
rect 15470 20040 15476 20052
rect 14967 20012 15476 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 15470 20000 15476 20012
rect 15528 20040 15534 20052
rect 15528 20012 16252 20040
rect 15528 20000 15534 20012
rect 2216 19975 2274 19981
rect 2216 19941 2228 19975
rect 2262 19972 2274 19975
rect 2406 19972 2412 19984
rect 2262 19944 2412 19972
rect 2262 19941 2274 19944
rect 2216 19935 2274 19941
rect 2406 19932 2412 19944
rect 2464 19932 2470 19984
rect 4706 19932 4712 19984
rect 4764 19972 4770 19984
rect 5813 19975 5871 19981
rect 5813 19972 5825 19975
rect 4764 19944 5825 19972
rect 4764 19932 4770 19944
rect 1946 19864 1952 19916
rect 2004 19864 2010 19916
rect 3418 19864 3424 19916
rect 3476 19864 3482 19916
rect 3510 19864 3516 19916
rect 3568 19904 3574 19916
rect 3677 19907 3735 19913
rect 3677 19904 3689 19907
rect 3568 19876 3689 19904
rect 3568 19864 3574 19876
rect 3677 19873 3689 19876
rect 3723 19873 3735 19907
rect 3677 19867 3735 19873
rect 5261 19907 5319 19913
rect 5261 19873 5273 19907
rect 5307 19904 5319 19907
rect 5350 19904 5356 19916
rect 5307 19876 5356 19904
rect 5307 19873 5319 19876
rect 5261 19867 5319 19873
rect 5350 19864 5356 19876
rect 5408 19864 5414 19916
rect 5460 19913 5488 19944
rect 5813 19941 5825 19944
rect 5859 19941 5871 19975
rect 5813 19935 5871 19941
rect 7190 19932 7196 19984
rect 7248 19972 7254 19984
rect 8202 19972 8208 19984
rect 7248 19944 8208 19972
rect 7248 19932 7254 19944
rect 8202 19932 8208 19944
rect 8260 19932 8266 19984
rect 8662 19932 8668 19984
rect 8720 19972 8726 19984
rect 9024 19975 9082 19981
rect 9024 19972 9036 19975
rect 8720 19944 9036 19972
rect 8720 19932 8726 19944
rect 9024 19941 9036 19944
rect 9070 19941 9082 19975
rect 11882 19972 11888 19984
rect 9024 19935 9082 19941
rect 11440 19944 11888 19972
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 5994 19864 6000 19916
rect 6052 19864 6058 19916
rect 6181 19907 6239 19913
rect 6181 19873 6193 19907
rect 6227 19873 6239 19907
rect 6181 19867 6239 19873
rect 4798 19796 4804 19848
rect 4856 19836 4862 19848
rect 6196 19836 6224 19867
rect 6270 19864 6276 19916
rect 6328 19864 6334 19916
rect 6454 19864 6460 19916
rect 6512 19904 6518 19916
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 6512 19876 7389 19904
rect 6512 19864 6518 19876
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 7650 19864 7656 19916
rect 7708 19904 7714 19916
rect 8018 19904 8024 19916
rect 7708 19876 8024 19904
rect 7708 19864 7714 19876
rect 8018 19864 8024 19876
rect 8076 19904 8082 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 8076 19876 8401 19904
rect 8076 19864 8082 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 8478 19864 8484 19916
rect 8536 19904 8542 19916
rect 8757 19907 8815 19913
rect 8757 19904 8769 19907
rect 8536 19876 8769 19904
rect 8536 19864 8542 19876
rect 8757 19873 8769 19876
rect 8803 19873 8815 19907
rect 8757 19867 8815 19873
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11440 19913 11468 19944
rect 11882 19932 11888 19944
rect 11940 19932 11946 19984
rect 15286 19932 15292 19984
rect 15344 19972 15350 19984
rect 15562 19972 15568 19984
rect 15344 19944 15568 19972
rect 15344 19932 15350 19944
rect 15562 19932 15568 19944
rect 15620 19932 15626 19984
rect 15930 19932 15936 19984
rect 15988 19972 15994 19984
rect 16224 19972 16252 20012
rect 16574 20000 16580 20052
rect 16632 20000 16638 20052
rect 17221 20043 17279 20049
rect 17221 20009 17233 20043
rect 17267 20040 17279 20043
rect 17678 20040 17684 20052
rect 17267 20012 17684 20040
rect 17267 20009 17279 20012
rect 17221 20003 17279 20009
rect 17678 20000 17684 20012
rect 17736 20040 17742 20052
rect 17954 20040 17960 20052
rect 17736 20012 17960 20040
rect 17736 20000 17742 20012
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 18233 20043 18291 20049
rect 18233 20009 18245 20043
rect 18279 20040 18291 20043
rect 18414 20040 18420 20052
rect 18279 20012 18420 20040
rect 18279 20009 18291 20012
rect 18233 20003 18291 20009
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 18966 20040 18972 20052
rect 18739 20012 18972 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 19426 20040 19432 20052
rect 19306 20012 19432 20040
rect 16485 19975 16543 19981
rect 16485 19972 16497 19975
rect 15988 19944 16160 19972
rect 16224 19944 16497 19972
rect 15988 19932 15994 19944
rect 11333 19907 11391 19913
rect 11333 19904 11345 19907
rect 11112 19876 11345 19904
rect 11112 19864 11118 19876
rect 11333 19873 11345 19876
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 11425 19907 11483 19913
rect 11425 19873 11437 19907
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 11517 19907 11575 19913
rect 11517 19873 11529 19907
rect 11563 19873 11575 19907
rect 11517 19867 11575 19873
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19873 11759 19907
rect 11701 19867 11759 19873
rect 6365 19839 6423 19845
rect 4856 19808 6316 19836
rect 4856 19796 4862 19808
rect 4890 19728 4896 19780
rect 4948 19768 4954 19780
rect 5994 19768 6000 19780
rect 4948 19740 6000 19768
rect 4948 19728 4954 19740
rect 5994 19728 6000 19740
rect 6052 19728 6058 19780
rect 3329 19703 3387 19709
rect 3329 19669 3341 19703
rect 3375 19700 3387 19703
rect 4062 19700 4068 19712
rect 3375 19672 4068 19700
rect 3375 19669 3387 19672
rect 3329 19663 3387 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 4801 19703 4859 19709
rect 4801 19700 4813 19703
rect 4212 19672 4813 19700
rect 4212 19660 4218 19672
rect 4801 19669 4813 19672
rect 4847 19669 4859 19703
rect 6288 19700 6316 19808
rect 6365 19805 6377 19839
rect 6411 19836 6423 19839
rect 7006 19836 7012 19848
rect 6411 19808 7012 19836
rect 6411 19805 6423 19808
rect 6365 19799 6423 19805
rect 7006 19796 7012 19808
rect 7064 19836 7070 19848
rect 7101 19839 7159 19845
rect 7101 19836 7113 19839
rect 7064 19808 7113 19836
rect 7064 19796 7070 19808
rect 7101 19805 7113 19808
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 7190 19796 7196 19848
rect 7248 19796 7254 19848
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 6546 19728 6552 19780
rect 6604 19768 6610 19780
rect 7300 19768 7328 19799
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11532 19836 11560 19867
rect 11296 19808 11560 19836
rect 11296 19796 11302 19808
rect 6604 19740 7328 19768
rect 6604 19728 6610 19740
rect 11146 19728 11152 19780
rect 11204 19768 11210 19780
rect 11716 19768 11744 19867
rect 13354 19864 13360 19916
rect 13412 19864 13418 19916
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 13556 19876 15393 19904
rect 13556 19836 13584 19876
rect 15381 19873 15393 19876
rect 15427 19873 15439 19907
rect 15381 19867 15439 19873
rect 12406 19808 13584 19836
rect 13633 19839 13691 19845
rect 12406 19768 12434 19808
rect 13633 19805 13645 19839
rect 13679 19836 13691 19839
rect 14550 19836 14556 19848
rect 13679 19808 14556 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 15396 19836 15424 19867
rect 15470 19864 15476 19916
rect 15528 19864 15534 19916
rect 15749 19907 15807 19913
rect 15749 19873 15761 19907
rect 15795 19904 15807 19907
rect 16022 19904 16028 19916
rect 15795 19876 16028 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16132 19913 16160 19944
rect 16485 19941 16497 19944
rect 16531 19941 16543 19975
rect 16592 19972 16620 20000
rect 17126 19972 17132 19984
rect 16592 19944 17132 19972
rect 16485 19935 16543 19941
rect 17126 19932 17132 19944
rect 17184 19972 17190 19984
rect 17184 19944 17356 19972
rect 17184 19932 17190 19944
rect 16298 19913 16304 19916
rect 16117 19907 16175 19913
rect 16117 19873 16129 19907
rect 16163 19873 16175 19907
rect 16117 19867 16175 19873
rect 16265 19907 16304 19913
rect 16265 19873 16277 19907
rect 16265 19867 16304 19873
rect 16298 19864 16304 19867
rect 16356 19864 16362 19916
rect 16390 19864 16396 19916
rect 16448 19864 16454 19916
rect 16666 19913 16672 19916
rect 16623 19907 16672 19913
rect 16623 19873 16635 19907
rect 16669 19873 16672 19907
rect 16623 19867 16672 19873
rect 16666 19864 16672 19867
rect 16724 19864 16730 19916
rect 16942 19864 16948 19916
rect 17000 19904 17006 19916
rect 17328 19913 17356 19944
rect 17586 19932 17592 19984
rect 17644 19932 17650 19984
rect 19306 19972 19334 20012
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 19797 20043 19855 20049
rect 19797 20009 19809 20043
rect 19843 20040 19855 20043
rect 20346 20040 20352 20052
rect 19843 20012 20352 20040
rect 19843 20009 19855 20012
rect 19797 20003 19855 20009
rect 18156 19944 19334 19972
rect 18156 19916 18184 19944
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 17000 19876 17049 19904
rect 17000 19864 17006 19876
rect 17037 19873 17049 19876
rect 17083 19873 17095 19907
rect 17037 19867 17095 19873
rect 17313 19907 17371 19913
rect 17313 19873 17325 19907
rect 17359 19904 17371 19907
rect 17359 19876 18092 19904
rect 17359 19873 17371 19876
rect 17313 19867 17371 19873
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 15396 19808 17417 19836
rect 17405 19805 17417 19808
rect 17451 19805 17463 19839
rect 18064 19836 18092 19876
rect 18138 19864 18144 19916
rect 18196 19864 18202 19916
rect 18417 19907 18475 19913
rect 18417 19873 18429 19907
rect 18463 19873 18475 19907
rect 18417 19867 18475 19873
rect 18432 19836 18460 19867
rect 18506 19864 18512 19916
rect 18564 19904 18570 19916
rect 18601 19907 18659 19913
rect 18601 19904 18613 19907
rect 18564 19876 18613 19904
rect 18564 19864 18570 19876
rect 18601 19873 18613 19876
rect 18647 19873 18659 19907
rect 18601 19867 18659 19873
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 18969 19907 19027 19913
rect 18969 19904 18981 19907
rect 18748 19876 18981 19904
rect 18748 19864 18754 19876
rect 18969 19873 18981 19876
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 19061 19907 19119 19913
rect 19061 19873 19073 19907
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 19153 19907 19211 19913
rect 19153 19873 19165 19907
rect 19199 19873 19211 19907
rect 19153 19867 19211 19873
rect 19076 19836 19104 19867
rect 18064 19808 18460 19836
rect 17405 19799 17463 19805
rect 11204 19740 12434 19768
rect 15933 19771 15991 19777
rect 11204 19728 11210 19740
rect 15933 19737 15945 19771
rect 15979 19768 15991 19771
rect 16574 19768 16580 19780
rect 15979 19740 16580 19768
rect 15979 19737 15991 19740
rect 15933 19731 15991 19737
rect 16574 19728 16580 19740
rect 16632 19728 16638 19780
rect 16761 19771 16819 19777
rect 16761 19737 16773 19771
rect 16807 19768 16819 19771
rect 17586 19768 17592 19780
rect 16807 19740 17592 19768
rect 16807 19737 16819 19740
rect 16761 19731 16819 19737
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 9766 19700 9772 19712
rect 6288 19672 9772 19700
rect 4801 19663 4859 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 15197 19703 15255 19709
rect 15197 19669 15209 19703
rect 15243 19700 15255 19703
rect 15286 19700 15292 19712
rect 15243 19672 15292 19700
rect 15243 19669 15255 19672
rect 15197 19663 15255 19669
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 16390 19700 16396 19712
rect 15528 19672 16396 19700
rect 15528 19660 15534 19672
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 16482 19660 16488 19712
rect 16540 19700 16546 19712
rect 16853 19703 16911 19709
rect 16853 19700 16865 19703
rect 16540 19672 16865 19700
rect 16540 19660 16546 19672
rect 16853 19669 16865 19672
rect 16899 19669 16911 19703
rect 18432 19700 18460 19808
rect 18708 19808 19104 19836
rect 19168 19836 19196 19867
rect 19334 19864 19340 19916
rect 19392 19864 19398 19916
rect 19610 19864 19616 19916
rect 19668 19864 19674 19916
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 19168 19808 19441 19836
rect 18509 19771 18567 19777
rect 18509 19737 18521 19771
rect 18555 19768 18567 19771
rect 18708 19768 18736 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 18555 19740 18736 19768
rect 18555 19737 18567 19740
rect 18509 19731 18567 19737
rect 19058 19728 19064 19780
rect 19116 19768 19122 19780
rect 19812 19768 19840 20003
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 22186 20000 22192 20052
rect 22244 20040 22250 20052
rect 26418 20040 26424 20052
rect 22244 20012 26424 20040
rect 22244 20000 22250 20012
rect 26418 20000 26424 20012
rect 26476 20000 26482 20052
rect 29178 20040 29184 20052
rect 27908 20012 29184 20040
rect 22830 19932 22836 19984
rect 22888 19972 22894 19984
rect 23845 19975 23903 19981
rect 22888 19944 23428 19972
rect 22888 19932 22894 19944
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19902 19947 19907
rect 20898 19904 20904 19916
rect 19996 19902 20904 19904
rect 19935 19876 20904 19902
rect 19935 19874 20024 19876
rect 19935 19873 19947 19874
rect 19889 19867 19947 19873
rect 19116 19740 19840 19768
rect 19116 19728 19122 19740
rect 19996 19700 20024 19874
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 21542 19864 21548 19916
rect 21600 19864 21606 19916
rect 22186 19864 22192 19916
rect 22244 19904 22250 19916
rect 22649 19913 22707 19919
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 22244 19876 22293 19904
rect 22244 19864 22250 19876
rect 22281 19873 22293 19876
rect 22327 19873 22339 19907
rect 22281 19867 22339 19873
rect 22373 19907 22431 19913
rect 22373 19873 22385 19907
rect 22419 19873 22431 19907
rect 22373 19867 22431 19873
rect 22484 19907 22542 19913
rect 22484 19873 22496 19907
rect 22530 19873 22542 19907
rect 22649 19879 22661 19913
rect 22695 19910 22707 19913
rect 22695 19882 22784 19910
rect 22695 19879 22707 19882
rect 22649 19873 22707 19879
rect 22484 19867 22542 19873
rect 22278 19728 22284 19780
rect 22336 19768 22342 19780
rect 22376 19768 22404 19867
rect 22336 19740 22404 19768
rect 22499 19768 22527 19867
rect 22756 19848 22784 19882
rect 23106 19864 23112 19916
rect 23164 19864 23170 19916
rect 23198 19864 23204 19916
rect 23256 19864 23262 19916
rect 23400 19913 23428 19944
rect 23845 19941 23857 19975
rect 23891 19972 23903 19975
rect 24210 19972 24216 19984
rect 23891 19944 24216 19972
rect 23891 19941 23903 19944
rect 23845 19935 23903 19941
rect 24210 19932 24216 19944
rect 24268 19932 24274 19984
rect 27522 19932 27528 19984
rect 27580 19972 27586 19984
rect 27908 19981 27936 20012
rect 29178 20000 29184 20012
rect 29236 20000 29242 20052
rect 29454 20000 29460 20052
rect 29512 20000 29518 20052
rect 27893 19975 27951 19981
rect 27893 19972 27905 19975
rect 27580 19944 27905 19972
rect 27580 19932 27586 19944
rect 27893 19941 27905 19944
rect 27939 19941 27951 19975
rect 29638 19972 29644 19984
rect 27893 19935 27951 19941
rect 29196 19944 29644 19972
rect 23385 19907 23443 19913
rect 23385 19873 23397 19907
rect 23431 19873 23443 19907
rect 23385 19867 23443 19873
rect 23474 19864 23480 19916
rect 23532 19864 23538 19916
rect 23750 19864 23756 19916
rect 23808 19864 23814 19916
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19873 23995 19907
rect 23937 19867 23995 19873
rect 22738 19796 22744 19848
rect 22796 19796 22802 19848
rect 22830 19796 22836 19848
rect 22888 19836 22894 19848
rect 22925 19839 22983 19845
rect 22925 19836 22937 19839
rect 22888 19808 22937 19836
rect 22888 19796 22894 19808
rect 22925 19805 22937 19808
rect 22971 19805 22983 19839
rect 23124 19836 23152 19864
rect 23952 19836 23980 19867
rect 24118 19864 24124 19916
rect 24176 19864 24182 19916
rect 25774 19864 25780 19916
rect 25832 19904 25838 19916
rect 27709 19907 27767 19913
rect 27709 19904 27721 19907
rect 25832 19876 27721 19904
rect 25832 19864 25838 19876
rect 27709 19873 27721 19876
rect 27755 19873 27767 19907
rect 27709 19867 27767 19873
rect 27982 19864 27988 19916
rect 28040 19904 28046 19916
rect 28810 19904 28816 19916
rect 28040 19876 28816 19904
rect 28040 19864 28046 19876
rect 28810 19864 28816 19876
rect 28868 19864 28874 19916
rect 29196 19913 29224 19944
rect 29638 19932 29644 19944
rect 29696 19932 29702 19984
rect 28997 19907 29055 19913
rect 28997 19873 29009 19907
rect 29043 19873 29055 19907
rect 28997 19867 29055 19873
rect 29089 19907 29147 19913
rect 29089 19873 29101 19907
rect 29135 19873 29147 19907
rect 29089 19867 29147 19873
rect 29181 19907 29239 19913
rect 29181 19873 29193 19907
rect 29227 19873 29239 19907
rect 29181 19867 29239 19873
rect 23124 19808 23980 19836
rect 22925 19799 22983 19805
rect 25590 19796 25596 19848
rect 25648 19836 25654 19848
rect 25685 19839 25743 19845
rect 25685 19836 25697 19839
rect 25648 19808 25697 19836
rect 25648 19796 25654 19808
rect 25685 19805 25697 19808
rect 25731 19805 25743 19839
rect 25685 19799 25743 19805
rect 25866 19768 25872 19780
rect 22499 19740 25872 19768
rect 22336 19728 22342 19740
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 18432 19672 20024 19700
rect 16853 19663 16911 19669
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 21453 19703 21511 19709
rect 21453 19700 21465 19703
rect 21324 19672 21465 19700
rect 21324 19660 21330 19672
rect 21453 19669 21465 19672
rect 21499 19669 21511 19703
rect 21453 19663 21511 19669
rect 22738 19660 22744 19712
rect 22796 19700 22802 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 22796 19672 22845 19700
rect 22796 19660 22802 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 22833 19663 22891 19669
rect 23014 19660 23020 19712
rect 23072 19700 23078 19712
rect 23569 19703 23627 19709
rect 23569 19700 23581 19703
rect 23072 19672 23581 19700
rect 23072 19660 23078 19672
rect 23569 19669 23581 19672
rect 23615 19669 23627 19703
rect 23569 19663 23627 19669
rect 25130 19660 25136 19712
rect 25188 19660 25194 19712
rect 27430 19660 27436 19712
rect 27488 19700 27494 19712
rect 27617 19703 27675 19709
rect 27617 19700 27629 19703
rect 27488 19672 27629 19700
rect 27488 19660 27494 19672
rect 27617 19669 27629 19672
rect 27663 19669 27675 19703
rect 27617 19663 27675 19669
rect 27982 19660 27988 19712
rect 28040 19660 28046 19712
rect 29012 19700 29040 19867
rect 29104 19836 29132 19867
rect 29546 19864 29552 19916
rect 29604 19864 29610 19916
rect 29822 19913 29828 19916
rect 29816 19867 29828 19913
rect 29822 19864 29828 19867
rect 29880 19864 29886 19916
rect 29362 19836 29368 19848
rect 29104 19808 29368 19836
rect 29362 19796 29368 19808
rect 29420 19796 29426 19848
rect 29730 19700 29736 19712
rect 29012 19672 29736 19700
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 29914 19660 29920 19712
rect 29972 19700 29978 19712
rect 30929 19703 30987 19709
rect 30929 19700 30941 19703
rect 29972 19672 30941 19700
rect 29972 19660 29978 19672
rect 30929 19669 30941 19672
rect 30975 19669 30987 19703
rect 30929 19663 30987 19669
rect 552 19610 31648 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 11436 19610
rect 11488 19558 11500 19610
rect 11552 19558 11564 19610
rect 11616 19558 11628 19610
rect 11680 19558 11692 19610
rect 11744 19558 19210 19610
rect 19262 19558 19274 19610
rect 19326 19558 19338 19610
rect 19390 19558 19402 19610
rect 19454 19558 19466 19610
rect 19518 19558 26984 19610
rect 27036 19558 27048 19610
rect 27100 19558 27112 19610
rect 27164 19558 27176 19610
rect 27228 19558 27240 19610
rect 27292 19558 31648 19610
rect 552 19536 31648 19558
rect 2406 19456 2412 19508
rect 2464 19456 2470 19508
rect 6270 19496 6276 19508
rect 3068 19468 6276 19496
rect 3068 19360 3096 19468
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 6454 19456 6460 19508
rect 6512 19456 6518 19508
rect 9033 19499 9091 19505
rect 9033 19465 9045 19499
rect 9079 19496 9091 19499
rect 9766 19496 9772 19508
rect 9079 19468 9772 19496
rect 9079 19465 9091 19468
rect 9033 19459 9091 19465
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 15654 19456 15660 19508
rect 15712 19496 15718 19508
rect 16117 19499 16175 19505
rect 16117 19496 16129 19499
rect 15712 19468 16129 19496
rect 15712 19456 15718 19468
rect 16117 19465 16129 19468
rect 16163 19465 16175 19499
rect 16117 19459 16175 19465
rect 16301 19499 16359 19505
rect 16301 19465 16313 19499
rect 16347 19496 16359 19499
rect 16577 19499 16635 19505
rect 16577 19496 16589 19499
rect 16347 19468 16589 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 16577 19465 16589 19468
rect 16623 19465 16635 19499
rect 16577 19459 16635 19465
rect 16758 19456 16764 19508
rect 16816 19456 16822 19508
rect 17218 19496 17224 19508
rect 16859 19468 17224 19496
rect 3234 19388 3240 19440
rect 3292 19428 3298 19440
rect 3292 19400 5764 19428
rect 3292 19388 3298 19400
rect 2424 19332 3096 19360
rect 2424 19304 2452 19332
rect 3068 19304 3096 19332
rect 3142 19320 3148 19372
rect 3200 19360 3206 19372
rect 3973 19363 4031 19369
rect 3200 19332 3556 19360
rect 3200 19320 3206 19332
rect 1946 19252 1952 19304
rect 2004 19252 2010 19304
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19261 2099 19295
rect 2041 19255 2099 19261
rect 2056 19224 2084 19255
rect 2130 19252 2136 19304
rect 2188 19252 2194 19304
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 2406 19292 2412 19304
rect 2363 19264 2412 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2406 19252 2412 19264
rect 2464 19252 2470 19304
rect 2498 19252 2504 19304
rect 2556 19292 2562 19304
rect 2685 19295 2743 19301
rect 2685 19292 2697 19295
rect 2556 19264 2697 19292
rect 2556 19252 2562 19264
rect 2685 19261 2697 19264
rect 2731 19261 2743 19295
rect 2685 19255 2743 19261
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19261 2835 19295
rect 2777 19255 2835 19261
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19261 2927 19295
rect 2869 19255 2927 19261
rect 2590 19224 2596 19236
rect 2056 19196 2596 19224
rect 2590 19184 2596 19196
rect 2648 19224 2654 19236
rect 2792 19224 2820 19255
rect 2648 19196 2820 19224
rect 2884 19224 2912 19255
rect 3050 19252 3056 19304
rect 3108 19252 3114 19304
rect 3326 19252 3332 19304
rect 3384 19292 3390 19304
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 3384 19264 3433 19292
rect 3384 19252 3390 19264
rect 3421 19261 3433 19264
rect 3467 19261 3479 19295
rect 3528 19292 3556 19332
rect 3973 19329 3985 19363
rect 4019 19360 4031 19363
rect 4246 19360 4252 19372
rect 4019 19332 4252 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4246 19320 4252 19332
rect 4304 19360 4310 19372
rect 4890 19360 4896 19372
rect 4304 19332 4896 19360
rect 4304 19320 4310 19332
rect 4890 19320 4896 19332
rect 4948 19320 4954 19372
rect 3528 19264 3740 19292
rect 3421 19255 3479 19261
rect 3237 19227 3295 19233
rect 3237 19224 3249 19227
rect 2884 19196 3249 19224
rect 2648 19184 2654 19196
rect 3237 19193 3249 19196
rect 3283 19193 3295 19227
rect 3237 19187 3295 19193
rect 3602 19184 3608 19236
rect 3660 19184 3666 19236
rect 3712 19224 3740 19264
rect 4062 19252 4068 19304
rect 4120 19292 4126 19304
rect 4157 19295 4215 19301
rect 4157 19292 4169 19295
rect 4120 19264 4169 19292
rect 4120 19252 4126 19264
rect 4157 19261 4169 19264
rect 4203 19261 4215 19295
rect 5736 19292 5764 19400
rect 15562 19388 15568 19440
rect 15620 19428 15626 19440
rect 16482 19428 16488 19440
rect 15620 19400 16488 19428
rect 15620 19388 15626 19400
rect 16482 19388 16488 19400
rect 16540 19428 16546 19440
rect 16859 19428 16887 19468
rect 17218 19456 17224 19468
rect 17276 19496 17282 19508
rect 17276 19468 17540 19496
rect 17276 19456 17282 19468
rect 16540 19400 16887 19428
rect 16540 19388 16546 19400
rect 15013 19363 15071 19369
rect 6196 19332 6684 19360
rect 5810 19292 5816 19304
rect 5736 19264 5816 19292
rect 4157 19255 4215 19261
rect 5810 19252 5816 19264
rect 5868 19252 5874 19304
rect 5961 19295 6019 19301
rect 5961 19261 5973 19295
rect 6007 19292 6019 19295
rect 6196 19292 6224 19332
rect 6362 19301 6368 19304
rect 6007 19264 6224 19292
rect 6319 19295 6368 19301
rect 6007 19261 6019 19264
rect 5961 19255 6019 19261
rect 6319 19261 6331 19295
rect 6365 19261 6368 19295
rect 6319 19255 6368 19261
rect 6362 19252 6368 19255
rect 6420 19252 6426 19304
rect 6454 19252 6460 19304
rect 6512 19294 6518 19304
rect 6656 19302 6684 19332
rect 15013 19329 15025 19363
rect 15059 19360 15071 19363
rect 16114 19360 16120 19372
rect 15059 19332 16120 19360
rect 15059 19329 15071 19332
rect 15013 19323 15071 19329
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 17512 19360 17540 19468
rect 17586 19456 17592 19508
rect 17644 19456 17650 19508
rect 17681 19499 17739 19505
rect 17681 19465 17693 19499
rect 17727 19496 17739 19499
rect 18046 19496 18052 19508
rect 17727 19468 18052 19496
rect 17727 19465 17739 19468
rect 17681 19459 17739 19465
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 18230 19456 18236 19508
rect 18288 19496 18294 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 18288 19468 19073 19496
rect 18288 19456 18294 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 21174 19456 21180 19508
rect 21232 19496 21238 19508
rect 22830 19496 22836 19508
rect 21232 19468 22836 19496
rect 21232 19456 21238 19468
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 23198 19456 23204 19508
rect 23256 19496 23262 19508
rect 28074 19496 28080 19508
rect 23256 19468 28080 19496
rect 23256 19456 23262 19468
rect 28074 19456 28080 19468
rect 28132 19456 28138 19508
rect 29733 19499 29791 19505
rect 29733 19465 29745 19499
rect 29779 19496 29791 19499
rect 29822 19496 29828 19508
rect 29779 19468 29828 19496
rect 29779 19465 29791 19468
rect 29733 19459 29791 19465
rect 29822 19456 29828 19468
rect 29880 19456 29886 19508
rect 20254 19428 20260 19440
rect 18064 19400 20260 19428
rect 17681 19363 17739 19369
rect 17681 19360 17693 19363
rect 17512 19332 17693 19360
rect 17681 19329 17693 19332
rect 17727 19360 17739 19363
rect 18064 19360 18092 19400
rect 20254 19388 20260 19400
rect 20312 19388 20318 19440
rect 20530 19388 20536 19440
rect 20588 19428 20594 19440
rect 22005 19431 22063 19437
rect 22005 19428 22017 19431
rect 20588 19400 22017 19428
rect 20588 19388 20594 19400
rect 22005 19397 22017 19400
rect 22051 19397 22063 19431
rect 29454 19428 29460 19440
rect 22005 19391 22063 19397
rect 28736 19400 29460 19428
rect 19702 19360 19708 19372
rect 17727 19332 18092 19360
rect 19076 19332 19708 19360
rect 17727 19329 17739 19332
rect 17681 19323 17739 19329
rect 6741 19305 6799 19311
rect 6741 19302 6753 19305
rect 6549 19295 6607 19301
rect 6549 19294 6561 19295
rect 6512 19266 6561 19294
rect 6512 19252 6518 19266
rect 6549 19261 6561 19266
rect 6595 19261 6607 19295
rect 6656 19274 6753 19302
rect 6741 19271 6753 19274
rect 6787 19302 6799 19305
rect 6787 19292 6868 19302
rect 6914 19292 6920 19304
rect 6787 19274 6920 19292
rect 6787 19271 6799 19274
rect 6741 19265 6799 19271
rect 6840 19264 6920 19274
rect 6549 19255 6607 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 8202 19252 8208 19304
rect 8260 19292 8266 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8260 19264 9045 19292
rect 8260 19252 8266 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19292 9275 19295
rect 10226 19292 10232 19304
rect 9263 19264 10232 19292
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 10226 19252 10232 19264
rect 10284 19252 10290 19304
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 11112 19264 11161 19292
rect 11112 19252 11118 19264
rect 11149 19261 11161 19264
rect 11195 19261 11207 19295
rect 11149 19255 11207 19261
rect 14550 19252 14556 19304
rect 14608 19252 14614 19304
rect 14734 19252 14740 19304
rect 14792 19252 14798 19304
rect 14826 19252 14832 19304
rect 14884 19292 14890 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14884 19264 14933 19292
rect 14884 19252 14890 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19261 15163 19295
rect 15105 19255 15163 19261
rect 4706 19224 4712 19236
rect 3712 19196 4712 19224
rect 1673 19159 1731 19165
rect 1673 19125 1685 19159
rect 1719 19156 1731 19159
rect 3510 19156 3516 19168
rect 1719 19128 3516 19156
rect 1719 19125 1731 19128
rect 1673 19119 1731 19125
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 4080 19165 4108 19196
rect 4706 19184 4712 19196
rect 4764 19184 4770 19236
rect 5074 19184 5080 19236
rect 5132 19224 5138 19236
rect 6089 19227 6147 19233
rect 6089 19224 6101 19227
rect 5132 19196 6101 19224
rect 5132 19184 5138 19196
rect 6089 19193 6101 19196
rect 6135 19193 6147 19227
rect 6089 19187 6147 19193
rect 6178 19184 6184 19236
rect 6236 19184 6242 19236
rect 6638 19184 6644 19236
rect 6696 19184 6702 19236
rect 15120 19224 15148 19255
rect 15286 19252 15292 19304
rect 15344 19252 15350 19304
rect 15657 19295 15715 19301
rect 15657 19261 15669 19295
rect 15703 19261 15715 19295
rect 15657 19255 15715 19261
rect 15381 19227 15439 19233
rect 15381 19224 15393 19227
rect 15120 19196 15393 19224
rect 15381 19193 15393 19196
rect 15427 19193 15439 19227
rect 15672 19224 15700 19255
rect 15746 19252 15752 19304
rect 15804 19252 15810 19304
rect 15838 19252 15844 19304
rect 15896 19252 15902 19304
rect 16022 19252 16028 19304
rect 16080 19252 16086 19304
rect 16758 19292 16764 19304
rect 16132 19264 16764 19292
rect 16132 19224 16160 19264
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 16850 19252 16856 19304
rect 16908 19252 16914 19304
rect 17126 19252 17132 19304
rect 17184 19252 17190 19304
rect 17218 19252 17224 19304
rect 17276 19252 17282 19304
rect 17586 19301 17592 19304
rect 17415 19295 17473 19301
rect 17415 19261 17427 19295
rect 17461 19261 17473 19295
rect 17415 19255 17473 19261
rect 17543 19295 17592 19301
rect 17543 19261 17555 19295
rect 17589 19261 17592 19295
rect 17543 19255 17592 19261
rect 15672 19196 16160 19224
rect 16285 19227 16343 19233
rect 15381 19187 15439 19193
rect 16285 19193 16297 19227
rect 16331 19224 16343 19227
rect 16390 19224 16396 19236
rect 16331 19196 16396 19224
rect 16331 19193 16343 19196
rect 16285 19187 16343 19193
rect 16390 19184 16396 19196
rect 16448 19184 16454 19236
rect 16485 19227 16543 19233
rect 16485 19193 16497 19227
rect 16531 19224 16543 19227
rect 16942 19224 16948 19236
rect 16531 19196 16948 19224
rect 16531 19193 16543 19196
rect 16485 19187 16543 19193
rect 16942 19184 16948 19196
rect 17000 19184 17006 19236
rect 17034 19184 17040 19236
rect 17092 19224 17098 19236
rect 17420 19224 17448 19255
rect 17586 19252 17592 19255
rect 17644 19252 17650 19304
rect 17862 19252 17868 19304
rect 17920 19252 17926 19304
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19076 19292 19104 19332
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 21140 19332 22293 19360
rect 21140 19320 21146 19332
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 22281 19323 22339 19329
rect 22370 19320 22376 19372
rect 22428 19360 22434 19372
rect 25774 19360 25780 19372
rect 22428 19332 22508 19360
rect 22428 19320 22434 19332
rect 19024 19264 19104 19292
rect 19024 19252 19030 19264
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19208 19264 19334 19292
rect 19208 19252 19214 19264
rect 17092 19196 17448 19224
rect 19306 19224 19334 19264
rect 19610 19252 19616 19304
rect 19668 19292 19674 19304
rect 21818 19292 21824 19304
rect 19668 19264 21824 19292
rect 19668 19252 19674 19264
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 22480 19301 22508 19332
rect 24780 19332 25780 19360
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 22443 19264 22477 19292
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19292 22615 19295
rect 22646 19292 22652 19304
rect 22603 19264 22652 19292
rect 22603 19261 22615 19264
rect 22557 19255 22615 19261
rect 22646 19252 22652 19264
rect 22704 19252 22710 19304
rect 22738 19252 22744 19304
rect 22796 19252 22802 19304
rect 22833 19295 22891 19301
rect 22833 19261 22845 19295
rect 22879 19292 22891 19295
rect 23014 19292 23020 19304
rect 22879 19264 23020 19292
rect 22879 19261 22891 19264
rect 22833 19255 22891 19261
rect 23014 19252 23020 19264
rect 23072 19252 23078 19304
rect 24397 19295 24455 19301
rect 24397 19261 24409 19295
rect 24443 19292 24455 19295
rect 24780 19292 24808 19332
rect 25774 19320 25780 19332
rect 25832 19320 25838 19372
rect 25866 19320 25872 19372
rect 25924 19320 25930 19372
rect 26436 19332 27568 19360
rect 24443 19264 24808 19292
rect 24443 19261 24455 19264
rect 24397 19255 24455 19261
rect 25314 19252 25320 19304
rect 25372 19252 25378 19304
rect 25498 19301 25504 19304
rect 25476 19295 25504 19301
rect 25476 19261 25488 19295
rect 25476 19255 25504 19261
rect 25498 19252 25504 19255
rect 25556 19252 25562 19304
rect 25590 19252 25596 19304
rect 25648 19252 25654 19304
rect 26329 19295 26387 19301
rect 26329 19261 26341 19295
rect 26375 19292 26387 19295
rect 26436 19292 26464 19332
rect 26375 19264 26464 19292
rect 26513 19295 26571 19301
rect 26375 19261 26387 19264
rect 26329 19255 26387 19261
rect 26513 19261 26525 19295
rect 26559 19261 26571 19295
rect 26513 19255 26571 19261
rect 19794 19224 19800 19236
rect 19306 19196 19800 19224
rect 17092 19184 17098 19196
rect 19794 19184 19800 19196
rect 19852 19184 19858 19236
rect 21085 19227 21143 19233
rect 21085 19193 21097 19227
rect 21131 19193 21143 19227
rect 21085 19187 21143 19193
rect 21637 19227 21695 19233
rect 21637 19193 21649 19227
rect 21683 19224 21695 19227
rect 22370 19224 22376 19236
rect 21683 19196 22376 19224
rect 21683 19193 21695 19196
rect 21637 19187 21695 19193
rect 4065 19159 4123 19165
rect 4065 19125 4077 19159
rect 4111 19156 4123 19159
rect 4154 19156 4160 19168
rect 4111 19128 4160 19156
rect 4111 19125 4123 19128
rect 4065 19119 4123 19125
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4525 19159 4583 19165
rect 4525 19125 4537 19159
rect 4571 19156 4583 19159
rect 6270 19156 6276 19168
rect 4571 19128 6276 19156
rect 4571 19125 4583 19128
rect 4525 19119 4583 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 11241 19159 11299 19165
rect 11241 19125 11253 19159
rect 11287 19156 11299 19159
rect 11422 19156 11428 19168
rect 11287 19128 11428 19156
rect 11287 19125 11299 19128
rect 11241 19119 11299 19125
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 17221 19159 17279 19165
rect 17221 19156 17233 19159
rect 15804 19128 17233 19156
rect 15804 19116 15810 19128
rect 17221 19125 17233 19128
rect 17267 19125 17279 19159
rect 17221 19119 17279 19125
rect 20990 19116 20996 19168
rect 21048 19116 21054 19168
rect 21100 19156 21128 19187
rect 22370 19184 22376 19196
rect 22428 19184 22434 19236
rect 23109 19227 23167 19233
rect 23109 19224 23121 19227
rect 22572 19196 23121 19224
rect 21358 19156 21364 19168
rect 21100 19128 21364 19156
rect 21358 19116 21364 19128
rect 21416 19156 21422 19168
rect 22572 19156 22600 19196
rect 23109 19193 23121 19196
rect 23155 19193 23167 19227
rect 26528 19224 26556 19255
rect 26694 19252 26700 19304
rect 26752 19252 26758 19304
rect 26878 19252 26884 19304
rect 26936 19252 26942 19304
rect 26970 19252 26976 19304
rect 27028 19252 27034 19304
rect 27065 19295 27123 19301
rect 27065 19261 27077 19295
rect 27111 19261 27123 19295
rect 27065 19255 27123 19261
rect 26786 19224 26792 19236
rect 26528 19196 26792 19224
rect 23109 19187 23167 19193
rect 26786 19184 26792 19196
rect 26844 19184 26850 19236
rect 21416 19128 22600 19156
rect 21416 19116 21422 19128
rect 23014 19116 23020 19168
rect 23072 19116 23078 19168
rect 24489 19159 24547 19165
rect 24489 19125 24501 19159
rect 24535 19156 24547 19159
rect 24578 19156 24584 19168
rect 24535 19128 24584 19156
rect 24535 19125 24547 19128
rect 24489 19119 24547 19125
rect 24578 19116 24584 19128
rect 24636 19116 24642 19168
rect 24670 19116 24676 19168
rect 24728 19116 24734 19168
rect 25038 19116 25044 19168
rect 25096 19156 25102 19168
rect 25498 19156 25504 19168
rect 25096 19128 25504 19156
rect 25096 19116 25102 19128
rect 25498 19116 25504 19128
rect 25556 19156 25562 19168
rect 27080 19156 27108 19255
rect 27430 19252 27436 19304
rect 27488 19252 27494 19304
rect 27540 19292 27568 19332
rect 28736 19292 28764 19400
rect 29454 19388 29460 19400
rect 29512 19428 29518 19440
rect 29914 19428 29920 19440
rect 29512 19400 29920 19428
rect 29512 19388 29518 19400
rect 29914 19388 29920 19400
rect 29972 19388 29978 19440
rect 28810 19320 28816 19372
rect 28868 19360 28874 19372
rect 28868 19332 30512 19360
rect 28868 19320 28874 19332
rect 27540 19264 28764 19292
rect 29086 19252 29092 19304
rect 29144 19252 29150 19304
rect 29273 19295 29331 19301
rect 29273 19261 29285 19295
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 27341 19227 27399 19233
rect 27341 19193 27353 19227
rect 27387 19224 27399 19227
rect 27678 19227 27736 19233
rect 27678 19224 27690 19227
rect 27387 19196 27690 19224
rect 27387 19193 27399 19196
rect 27341 19187 27399 19193
rect 27678 19193 27690 19196
rect 27724 19193 27736 19227
rect 29288 19224 29316 19255
rect 29362 19252 29368 19304
rect 29420 19252 29426 19304
rect 29454 19252 29460 19304
rect 29512 19252 29518 19304
rect 29822 19252 29828 19304
rect 29880 19292 29886 19304
rect 30009 19295 30067 19301
rect 30009 19292 30021 19295
rect 29880 19264 30021 19292
rect 29880 19252 29886 19264
rect 30009 19261 30021 19264
rect 30055 19261 30067 19295
rect 30009 19255 30067 19261
rect 30101 19295 30159 19301
rect 30101 19261 30113 19295
rect 30147 19292 30159 19295
rect 30190 19292 30196 19304
rect 30147 19264 30196 19292
rect 30147 19261 30159 19264
rect 30101 19255 30159 19261
rect 30190 19252 30196 19264
rect 30248 19252 30254 19304
rect 30282 19252 30288 19304
rect 30340 19252 30346 19304
rect 30374 19252 30380 19304
rect 30432 19252 30438 19304
rect 30484 19301 30512 19332
rect 30469 19295 30527 19301
rect 30469 19261 30481 19295
rect 30515 19261 30527 19295
rect 30469 19255 30527 19261
rect 29914 19224 29920 19236
rect 29288 19196 29920 19224
rect 27678 19187 27736 19193
rect 29914 19184 29920 19196
rect 29972 19184 29978 19236
rect 28813 19159 28871 19165
rect 28813 19156 28825 19159
rect 25556 19128 28825 19156
rect 25556 19116 25562 19128
rect 28813 19125 28825 19128
rect 28859 19156 28871 19159
rect 29362 19156 29368 19168
rect 28859 19128 29368 19156
rect 28859 19125 28871 19128
rect 28813 19119 28871 19125
rect 29362 19116 29368 19128
rect 29420 19116 29426 19168
rect 29730 19116 29736 19168
rect 29788 19156 29794 19168
rect 29825 19159 29883 19165
rect 29825 19156 29837 19159
rect 29788 19128 29837 19156
rect 29788 19116 29794 19128
rect 29825 19125 29837 19128
rect 29871 19125 29883 19159
rect 29825 19119 29883 19125
rect 30650 19116 30656 19168
rect 30708 19116 30714 19168
rect 552 19066 31648 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 12096 19066
rect 12148 19014 12160 19066
rect 12212 19014 12224 19066
rect 12276 19014 12288 19066
rect 12340 19014 12352 19066
rect 12404 19014 19870 19066
rect 19922 19014 19934 19066
rect 19986 19014 19998 19066
rect 20050 19014 20062 19066
rect 20114 19014 20126 19066
rect 20178 19014 27644 19066
rect 27696 19014 27708 19066
rect 27760 19014 27772 19066
rect 27824 19014 27836 19066
rect 27888 19014 27900 19066
rect 27952 19014 31648 19066
rect 552 18992 31648 19014
rect 2130 18912 2136 18964
rect 2188 18952 2194 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 2188 18924 2329 18952
rect 2188 18912 2194 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 5074 18912 5080 18964
rect 5132 18912 5138 18964
rect 5166 18912 5172 18964
rect 5224 18952 5230 18964
rect 6178 18952 6184 18964
rect 5224 18924 6184 18952
rect 5224 18912 5230 18924
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 6546 18952 6552 18964
rect 6503 18924 6552 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 7190 18912 7196 18964
rect 7248 18912 7254 18964
rect 11238 18912 11244 18964
rect 11296 18912 11302 18964
rect 13814 18912 13820 18964
rect 13872 18952 13878 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 13872 18924 14473 18952
rect 13872 18912 13878 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 14461 18915 14519 18921
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 16540 18912 16574 18952
rect 17310 18912 17316 18964
rect 17368 18912 17374 18964
rect 17497 18955 17555 18961
rect 17497 18921 17509 18955
rect 17543 18952 17555 18955
rect 17586 18952 17592 18964
rect 17543 18924 17592 18952
rect 17543 18921 17555 18924
rect 17497 18915 17555 18921
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 17828 18924 20484 18952
rect 17828 18912 17834 18924
rect 2958 18884 2964 18896
rect 2148 18856 2964 18884
rect 2148 18825 2176 18856
rect 2958 18844 2964 18856
rect 3016 18844 3022 18896
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 6086 18884 6092 18896
rect 5868 18856 6092 18884
rect 5868 18844 5874 18856
rect 6086 18844 6092 18856
rect 6144 18884 6150 18896
rect 6365 18887 6423 18893
rect 6144 18856 6316 18884
rect 6144 18844 6150 18856
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18816 2007 18819
rect 2133 18819 2191 18825
rect 1995 18788 2084 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 2056 18760 2084 18788
rect 2133 18785 2145 18819
rect 2179 18785 2191 18819
rect 2133 18779 2191 18785
rect 2406 18776 2412 18828
rect 2464 18776 2470 18828
rect 2590 18776 2596 18828
rect 2648 18776 2654 18828
rect 2682 18776 2688 18828
rect 2740 18776 2746 18828
rect 2777 18819 2835 18825
rect 2777 18785 2789 18819
rect 2823 18816 2835 18819
rect 3418 18816 3424 18828
rect 2823 18788 3424 18816
rect 2823 18785 2835 18788
rect 2777 18779 2835 18785
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18785 4307 18819
rect 4985 18819 5043 18825
rect 4985 18816 4997 18819
rect 4249 18779 4307 18785
rect 4632 18788 4997 18816
rect 2038 18708 2044 18760
rect 2096 18748 2102 18760
rect 3602 18748 3608 18760
rect 2096 18720 3608 18748
rect 2096 18708 2102 18720
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 3789 18751 3847 18757
rect 3789 18717 3801 18751
rect 3835 18717 3847 18751
rect 3789 18711 3847 18717
rect 3145 18683 3203 18689
rect 3145 18680 3157 18683
rect 2746 18652 3157 18680
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 2746 18612 2774 18652
rect 3145 18649 3157 18652
rect 3191 18649 3203 18683
rect 3145 18643 3203 18649
rect 3510 18640 3516 18692
rect 3568 18680 3574 18692
rect 3804 18680 3832 18711
rect 3970 18708 3976 18760
rect 4028 18708 4034 18760
rect 4154 18708 4160 18760
rect 4212 18708 4218 18760
rect 4264 18680 4292 18779
rect 4632 18689 4660 18788
rect 4985 18785 4997 18788
rect 5031 18785 5043 18819
rect 4985 18779 5043 18785
rect 5166 18776 5172 18828
rect 5224 18776 5230 18828
rect 6178 18776 6184 18828
rect 6236 18776 6242 18828
rect 6288 18816 6316 18856
rect 6365 18853 6377 18887
rect 6411 18884 6423 18887
rect 6411 18856 6960 18884
rect 6411 18853 6423 18856
rect 6365 18847 6423 18853
rect 6932 18828 6960 18856
rect 11422 18844 11428 18896
rect 11480 18844 11486 18896
rect 15194 18884 15200 18896
rect 14752 18856 15200 18884
rect 6457 18819 6515 18825
rect 6457 18816 6469 18819
rect 6288 18788 6469 18816
rect 6457 18785 6469 18788
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 6472 18748 6500 18779
rect 6914 18776 6920 18828
rect 6972 18816 6978 18828
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 6972 18788 7389 18816
rect 6972 18776 6978 18788
rect 7377 18785 7389 18788
rect 7423 18785 7435 18819
rect 7377 18779 7435 18785
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18816 7619 18819
rect 8110 18816 8116 18828
rect 7607 18788 8116 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 8110 18776 8116 18788
rect 8168 18776 8174 18828
rect 11054 18816 11060 18828
rect 9416 18788 11060 18816
rect 9416 18760 9444 18788
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 11790 18816 11796 18828
rect 11655 18788 11796 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 14752 18825 14780 18856
rect 15194 18844 15200 18856
rect 15252 18844 15258 18896
rect 16546 18884 16574 18912
rect 17328 18884 17356 18912
rect 19702 18884 19708 18896
rect 16546 18856 16712 18884
rect 17328 18856 19708 18884
rect 11885 18819 11943 18825
rect 11885 18785 11897 18819
rect 11931 18785 11943 18819
rect 11885 18779 11943 18785
rect 14737 18819 14795 18825
rect 14737 18785 14749 18819
rect 14783 18785 14795 18819
rect 14737 18779 14795 18785
rect 9398 18748 9404 18760
rect 6472 18720 9404 18748
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 10962 18708 10968 18760
rect 11020 18748 11026 18760
rect 11900 18748 11928 18779
rect 14826 18776 14832 18828
rect 14884 18776 14890 18828
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18785 14979 18819
rect 14921 18779 14979 18785
rect 15105 18819 15163 18825
rect 15105 18785 15117 18819
rect 15151 18816 15163 18819
rect 15286 18816 15292 18828
rect 15151 18788 15292 18816
rect 15151 18785 15163 18788
rect 15105 18779 15163 18785
rect 11020 18720 11928 18748
rect 14936 18748 14964 18779
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 15381 18819 15439 18825
rect 15381 18785 15393 18819
rect 15427 18785 15439 18819
rect 15381 18779 15439 18785
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18816 15531 18819
rect 15562 18816 15568 18828
rect 15519 18788 15568 18816
rect 15519 18785 15531 18788
rect 15473 18779 15531 18785
rect 15197 18751 15255 18757
rect 15197 18748 15209 18751
rect 14936 18720 15209 18748
rect 11020 18708 11026 18720
rect 15197 18717 15209 18720
rect 15243 18717 15255 18751
rect 15197 18711 15255 18717
rect 3568 18652 4292 18680
rect 4617 18683 4675 18689
rect 3568 18640 3574 18652
rect 4617 18649 4629 18683
rect 4663 18649 4675 18683
rect 4617 18643 4675 18649
rect 11330 18640 11336 18692
rect 11388 18680 11394 18692
rect 11701 18683 11759 18689
rect 11701 18680 11713 18683
rect 11388 18652 11713 18680
rect 11388 18640 11394 18652
rect 11701 18649 11713 18652
rect 11747 18649 11759 18683
rect 15396 18680 15424 18779
rect 15562 18776 15568 18788
rect 15620 18776 15626 18828
rect 15657 18819 15715 18825
rect 15657 18785 15669 18819
rect 15703 18785 15715 18819
rect 15657 18779 15715 18785
rect 15672 18748 15700 18779
rect 15746 18776 15752 18828
rect 15804 18776 15810 18828
rect 16114 18776 16120 18828
rect 16172 18776 16178 18828
rect 16684 18825 16712 18856
rect 19702 18844 19708 18856
rect 19760 18844 19766 18896
rect 16301 18819 16359 18825
rect 16301 18785 16313 18819
rect 16347 18785 16359 18819
rect 16577 18819 16635 18825
rect 16577 18806 16589 18819
rect 16301 18779 16359 18785
rect 16480 18785 16589 18806
rect 16623 18785 16635 18819
rect 16480 18779 16635 18785
rect 16669 18819 16727 18825
rect 16669 18785 16681 18819
rect 16715 18785 16727 18819
rect 16669 18779 16727 18785
rect 16853 18819 16911 18825
rect 16853 18785 16865 18819
rect 16899 18785 16911 18819
rect 16853 18779 16911 18785
rect 16206 18748 16212 18760
rect 15672 18720 16212 18748
rect 16206 18708 16212 18720
rect 16264 18748 16270 18760
rect 16316 18748 16344 18779
rect 16264 18720 16344 18748
rect 16480 18778 16620 18779
rect 16264 18708 16270 18720
rect 15838 18680 15844 18692
rect 15396 18652 15844 18680
rect 11701 18643 11759 18649
rect 15838 18640 15844 18652
rect 15896 18680 15902 18692
rect 16480 18680 16508 18778
rect 16868 18748 16896 18779
rect 16942 18776 16948 18828
rect 17000 18776 17006 18828
rect 17034 18776 17040 18828
rect 17092 18816 17098 18828
rect 17129 18819 17187 18825
rect 17129 18816 17141 18819
rect 17092 18788 17141 18816
rect 17092 18776 17098 18788
rect 17129 18785 17141 18788
rect 17175 18785 17187 18819
rect 17129 18779 17187 18785
rect 17218 18776 17224 18828
rect 17276 18776 17282 18828
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18816 17371 18819
rect 17678 18816 17684 18828
rect 17359 18788 17684 18816
rect 17359 18785 17371 18788
rect 17313 18779 17371 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18782 18816 18788 18828
rect 18104 18788 18788 18816
rect 18104 18776 18110 18788
rect 18782 18776 18788 18788
rect 18840 18816 18846 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 18840 18788 20085 18816
rect 18840 18776 18846 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 20073 18779 20131 18785
rect 20254 18776 20260 18828
rect 20312 18776 20318 18828
rect 20456 18825 20484 18924
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 22278 18952 22284 18964
rect 20956 18924 22284 18952
rect 20956 18912 20962 18924
rect 22278 18912 22284 18924
rect 22336 18912 22342 18964
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 22649 18955 22707 18961
rect 22649 18952 22661 18955
rect 22428 18924 22661 18952
rect 22428 18912 22434 18924
rect 22649 18921 22661 18924
rect 22695 18921 22707 18955
rect 25130 18952 25136 18964
rect 22649 18915 22707 18921
rect 24412 18924 25136 18952
rect 21542 18893 21548 18896
rect 21536 18884 21548 18893
rect 21503 18856 21548 18884
rect 21536 18847 21548 18856
rect 21542 18844 21548 18847
rect 21600 18844 21606 18896
rect 21818 18844 21824 18896
rect 21876 18884 21882 18896
rect 21876 18856 23888 18884
rect 21876 18844 21882 18856
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18816 20499 18819
rect 20530 18816 20536 18828
rect 20487 18788 20536 18816
rect 20487 18785 20499 18788
rect 20441 18779 20499 18785
rect 20530 18776 20536 18788
rect 20588 18776 20594 18828
rect 20622 18776 20628 18828
rect 20680 18776 20686 18828
rect 20714 18776 20720 18828
rect 20772 18776 20778 18828
rect 20809 18819 20867 18825
rect 20809 18785 20821 18819
rect 20855 18816 20867 18819
rect 20990 18816 20996 18828
rect 20855 18788 20996 18816
rect 20855 18785 20867 18788
rect 20809 18779 20867 18785
rect 17494 18748 17500 18760
rect 16868 18720 17500 18748
rect 17494 18708 17500 18720
rect 17552 18748 17558 18760
rect 18966 18748 18972 18760
rect 17552 18720 18972 18748
rect 17552 18708 17558 18720
rect 18966 18708 18972 18720
rect 19024 18708 19030 18760
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 20824 18748 20852 18779
rect 20990 18776 20996 18788
rect 21048 18776 21054 18828
rect 21266 18776 21272 18828
rect 21324 18776 21330 18828
rect 22922 18776 22928 18828
rect 22980 18776 22986 18828
rect 23860 18825 23888 18856
rect 23845 18819 23903 18825
rect 23845 18785 23857 18819
rect 23891 18785 23903 18819
rect 23845 18779 23903 18785
rect 19668 18720 20852 18748
rect 23860 18748 23888 18779
rect 24026 18776 24032 18828
rect 24084 18776 24090 18828
rect 24118 18776 24124 18828
rect 24176 18776 24182 18828
rect 24213 18819 24271 18825
rect 24213 18785 24225 18819
rect 24259 18816 24271 18819
rect 24412 18816 24440 18924
rect 25130 18912 25136 18924
rect 25188 18912 25194 18964
rect 25590 18912 25596 18964
rect 25648 18952 25654 18964
rect 25961 18955 26019 18961
rect 25961 18952 25973 18955
rect 25648 18924 25973 18952
rect 25648 18912 25654 18924
rect 25961 18921 25973 18924
rect 26007 18952 26019 18955
rect 26050 18952 26056 18964
rect 26007 18924 26056 18952
rect 26007 18921 26019 18924
rect 25961 18915 26019 18921
rect 26050 18912 26056 18924
rect 26108 18952 26114 18964
rect 26697 18955 26755 18961
rect 26697 18952 26709 18955
rect 26108 18924 26709 18952
rect 26108 18912 26114 18924
rect 26697 18921 26709 18924
rect 26743 18921 26755 18955
rect 26697 18915 26755 18921
rect 26878 18912 26884 18964
rect 26936 18952 26942 18964
rect 27249 18955 27307 18961
rect 27249 18952 27261 18955
rect 26936 18924 27261 18952
rect 26936 18912 26942 18924
rect 27249 18921 27261 18924
rect 27295 18921 27307 18955
rect 27249 18915 27307 18921
rect 27430 18912 27436 18964
rect 27488 18952 27494 18964
rect 27488 18924 28580 18952
rect 27488 18912 27494 18924
rect 24489 18887 24547 18893
rect 24489 18853 24501 18887
rect 24535 18884 24547 18887
rect 24826 18887 24884 18893
rect 24826 18884 24838 18887
rect 24535 18856 24838 18884
rect 24535 18853 24547 18856
rect 24489 18847 24547 18853
rect 24826 18853 24838 18856
rect 24872 18853 24884 18887
rect 27982 18884 27988 18896
rect 24826 18847 24884 18853
rect 26712 18856 27988 18884
rect 26712 18828 26740 18856
rect 27982 18844 27988 18856
rect 28040 18844 28046 18896
rect 24259 18788 24440 18816
rect 24259 18785 24271 18788
rect 24213 18779 24271 18785
rect 24578 18776 24584 18828
rect 24636 18776 24642 18828
rect 26694 18816 26700 18828
rect 24688 18788 26700 18816
rect 24688 18748 24716 18788
rect 26694 18776 26700 18788
rect 26752 18776 26758 18828
rect 26786 18776 26792 18828
rect 26844 18776 26850 18828
rect 27433 18819 27491 18825
rect 27433 18816 27445 18819
rect 27172 18788 27445 18816
rect 23860 18720 24716 18748
rect 26513 18751 26571 18757
rect 19668 18708 19674 18720
rect 26513 18717 26525 18751
rect 26559 18717 26571 18751
rect 26513 18711 26571 18717
rect 17310 18680 17316 18692
rect 15896 18652 17316 18680
rect 15896 18640 15902 18652
rect 17310 18640 17316 18652
rect 17368 18640 17374 18692
rect 17678 18640 17684 18692
rect 17736 18680 17742 18692
rect 20898 18680 20904 18692
rect 17736 18652 20904 18680
rect 17736 18640 17742 18652
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 26528 18680 26556 18711
rect 27172 18689 27200 18788
rect 27433 18785 27445 18788
rect 27479 18785 27491 18819
rect 27433 18779 27491 18785
rect 27522 18776 27528 18828
rect 27580 18776 27586 18828
rect 27706 18776 27712 18828
rect 27764 18776 27770 18828
rect 27798 18776 27804 18828
rect 27856 18776 27862 18828
rect 28074 18776 28080 18828
rect 28132 18816 28138 18828
rect 28552 18825 28580 18924
rect 29362 18912 29368 18964
rect 29420 18912 29426 18964
rect 29454 18912 29460 18964
rect 29512 18912 29518 18964
rect 29546 18912 29552 18964
rect 29604 18952 29610 18964
rect 29730 18952 29736 18964
rect 29604 18924 29736 18952
rect 29604 18912 29610 18924
rect 29730 18912 29736 18924
rect 29788 18912 29794 18964
rect 29822 18912 29828 18964
rect 29880 18912 29886 18964
rect 29914 18912 29920 18964
rect 29972 18912 29978 18964
rect 30374 18912 30380 18964
rect 30432 18952 30438 18964
rect 30432 18924 30512 18952
rect 30432 18912 30438 18924
rect 28997 18887 29055 18893
rect 28997 18853 29009 18887
rect 29043 18884 29055 18887
rect 30282 18884 30288 18896
rect 29043 18856 30288 18884
rect 29043 18853 29055 18856
rect 28997 18847 29055 18853
rect 30282 18844 30288 18856
rect 30340 18844 30346 18896
rect 28353 18819 28411 18825
rect 28353 18816 28365 18819
rect 28132 18788 28365 18816
rect 28132 18776 28138 18788
rect 28353 18785 28365 18788
rect 28399 18785 28411 18819
rect 28353 18779 28411 18785
rect 28537 18819 28595 18825
rect 28537 18785 28549 18819
rect 28583 18785 28595 18819
rect 28537 18779 28595 18785
rect 28626 18776 28632 18828
rect 28684 18776 28690 18828
rect 28721 18819 28779 18825
rect 28721 18785 28733 18819
rect 28767 18816 28779 18819
rect 29454 18816 29460 18828
rect 28767 18788 29460 18816
rect 28767 18785 28779 18788
rect 28721 18779 28779 18785
rect 29454 18776 29460 18788
rect 29512 18776 29518 18828
rect 30098 18776 30104 18828
rect 30156 18776 30162 18828
rect 30190 18776 30196 18828
rect 30248 18776 30254 18828
rect 30484 18825 30512 18924
rect 30377 18819 30435 18825
rect 30377 18785 30389 18819
rect 30423 18785 30435 18819
rect 30377 18779 30435 18785
rect 30469 18819 30527 18825
rect 30469 18785 30481 18819
rect 30515 18816 30527 18819
rect 30515 18788 30788 18816
rect 30515 18785 30527 18788
rect 30469 18779 30527 18785
rect 29178 18748 29184 18760
rect 27540 18720 29184 18748
rect 25516 18652 26556 18680
rect 25516 18624 25544 18652
rect 2188 18584 2774 18612
rect 3053 18615 3111 18621
rect 2188 18572 2194 18584
rect 3053 18581 3065 18615
rect 3099 18612 3111 18615
rect 4338 18612 4344 18624
rect 3099 18584 4344 18612
rect 3099 18581 3111 18584
rect 3053 18575 3111 18581
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 8202 18612 8208 18624
rect 7156 18584 8208 18612
rect 7156 18572 7162 18584
rect 8202 18572 8208 18584
rect 8260 18612 8266 18624
rect 15378 18612 15384 18624
rect 8260 18584 15384 18612
rect 8260 18572 8266 18584
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16482 18612 16488 18624
rect 16080 18584 16488 18612
rect 16080 18572 16086 18584
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 16761 18615 16819 18621
rect 16761 18612 16773 18615
rect 16724 18584 16773 18612
rect 16724 18572 16730 18584
rect 16761 18581 16773 18584
rect 16807 18581 16819 18615
rect 16761 18575 16819 18581
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 17862 18612 17868 18624
rect 17460 18584 17868 18612
rect 17460 18572 17466 18584
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 20165 18615 20223 18621
rect 20165 18581 20177 18615
rect 20211 18612 20223 18615
rect 20990 18612 20996 18624
rect 20211 18584 20996 18612
rect 20211 18581 20223 18584
rect 20165 18575 20223 18581
rect 20990 18572 20996 18584
rect 21048 18572 21054 18624
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 21542 18612 21548 18624
rect 21131 18584 21548 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 22830 18572 22836 18624
rect 22888 18572 22894 18624
rect 25498 18572 25504 18624
rect 25556 18572 25562 18624
rect 26528 18612 26556 18652
rect 27157 18683 27215 18689
rect 27157 18649 27169 18683
rect 27203 18649 27215 18683
rect 27157 18643 27215 18649
rect 27540 18612 27568 18720
rect 29178 18708 29184 18720
rect 29236 18708 29242 18760
rect 29546 18708 29552 18760
rect 29604 18748 29610 18760
rect 30392 18748 30420 18779
rect 29604 18720 30420 18748
rect 29604 18708 29610 18720
rect 29086 18640 29092 18692
rect 29144 18680 29150 18692
rect 30466 18680 30472 18692
rect 29144 18652 30472 18680
rect 29144 18640 29150 18652
rect 30466 18640 30472 18652
rect 30524 18680 30530 18692
rect 30650 18680 30656 18692
rect 30524 18652 30656 18680
rect 30524 18640 30530 18652
rect 30650 18640 30656 18652
rect 30708 18640 30714 18692
rect 26528 18584 27568 18612
rect 27798 18572 27804 18624
rect 27856 18612 27862 18624
rect 28810 18612 28816 18624
rect 27856 18584 28816 18612
rect 27856 18572 27862 18584
rect 28810 18572 28816 18584
rect 28868 18612 28874 18624
rect 30760 18612 30788 18788
rect 28868 18584 30788 18612
rect 28868 18572 28874 18584
rect 552 18522 31648 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 11436 18522
rect 11488 18470 11500 18522
rect 11552 18470 11564 18522
rect 11616 18470 11628 18522
rect 11680 18470 11692 18522
rect 11744 18470 19210 18522
rect 19262 18470 19274 18522
rect 19326 18470 19338 18522
rect 19390 18470 19402 18522
rect 19454 18470 19466 18522
rect 19518 18470 26984 18522
rect 27036 18470 27048 18522
rect 27100 18470 27112 18522
rect 27164 18470 27176 18522
rect 27228 18470 27240 18522
rect 27292 18470 31648 18522
rect 552 18448 31648 18470
rect 1489 18411 1547 18417
rect 1489 18377 1501 18411
rect 1535 18408 1547 18411
rect 2590 18408 2596 18420
rect 1535 18380 2596 18408
rect 1535 18377 1547 18380
rect 1489 18371 1547 18377
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 10502 18408 10508 18420
rect 5960 18380 10508 18408
rect 5960 18368 5966 18380
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 10962 18368 10968 18420
rect 11020 18368 11026 18420
rect 15286 18368 15292 18420
rect 15344 18368 15350 18420
rect 17402 18408 17408 18420
rect 15948 18380 17408 18408
rect 6914 18300 6920 18352
rect 6972 18300 6978 18352
rect 7116 18312 10088 18340
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 2222 18204 2228 18216
rect 1443 18176 2228 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2222 18164 2228 18176
rect 2280 18204 2286 18216
rect 2682 18204 2688 18216
rect 2280 18176 2688 18204
rect 2280 18164 2286 18176
rect 2682 18164 2688 18176
rect 2740 18164 2746 18216
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18204 3019 18207
rect 4617 18207 4675 18213
rect 4617 18204 4629 18207
rect 3007 18176 3280 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 1673 18139 1731 18145
rect 1673 18105 1685 18139
rect 1719 18105 1731 18139
rect 1673 18099 1731 18105
rect 1302 18028 1308 18080
rect 1360 18028 1366 18080
rect 1688 18068 1716 18099
rect 1854 18096 1860 18148
rect 1912 18136 1918 18148
rect 1949 18139 2007 18145
rect 1949 18136 1961 18139
rect 1912 18108 1961 18136
rect 1912 18096 1918 18108
rect 1949 18105 1961 18108
rect 1995 18136 2007 18139
rect 2038 18136 2044 18148
rect 1995 18108 2044 18136
rect 1995 18105 2007 18108
rect 1949 18099 2007 18105
rect 2038 18096 2044 18108
rect 2096 18096 2102 18148
rect 2130 18096 2136 18148
rect 2188 18096 2194 18148
rect 2317 18139 2375 18145
rect 2317 18105 2329 18139
rect 2363 18136 2375 18139
rect 2866 18136 2872 18148
rect 2363 18108 2872 18136
rect 2363 18105 2375 18108
rect 2317 18099 2375 18105
rect 2866 18096 2872 18108
rect 2924 18096 2930 18148
rect 3252 18077 3280 18176
rect 4264 18176 4629 18204
rect 4264 18148 4292 18176
rect 4617 18173 4629 18176
rect 4663 18173 4675 18207
rect 4617 18167 4675 18173
rect 6270 18164 6276 18216
rect 6328 18204 6334 18216
rect 7116 18204 7144 18312
rect 10060 18216 10088 18312
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 6328 18176 7144 18204
rect 7193 18207 7251 18213
rect 6328 18164 6334 18176
rect 7193 18173 7205 18207
rect 7239 18204 7251 18207
rect 7650 18204 7656 18216
rect 7239 18176 7656 18204
rect 7239 18173 7251 18176
rect 7193 18167 7251 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7742 18164 7748 18216
rect 7800 18164 7806 18216
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 7929 18207 7987 18213
rect 7929 18173 7941 18207
rect 7975 18173 7987 18207
rect 7929 18167 7987 18173
rect 8113 18207 8171 18213
rect 8113 18173 8125 18207
rect 8159 18204 8171 18207
rect 8202 18204 8208 18216
rect 8159 18176 8208 18204
rect 8159 18173 8171 18176
rect 8113 18167 8171 18173
rect 4246 18096 4252 18148
rect 4304 18096 4310 18148
rect 4338 18096 4344 18148
rect 4396 18145 4402 18148
rect 4396 18136 4408 18145
rect 6549 18139 6607 18145
rect 4396 18108 4441 18136
rect 4396 18099 4408 18108
rect 6549 18105 6561 18139
rect 6595 18136 6607 18139
rect 6638 18136 6644 18148
rect 6595 18108 6644 18136
rect 6595 18105 6607 18108
rect 6549 18099 6607 18105
rect 4396 18096 4402 18099
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 7374 18136 7380 18148
rect 7024 18108 7380 18136
rect 2409 18071 2467 18077
rect 2409 18068 2421 18071
rect 1688 18040 2421 18068
rect 2409 18037 2421 18040
rect 2455 18037 2467 18071
rect 2409 18031 2467 18037
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 3786 18068 3792 18080
rect 3283 18040 3792 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 3786 18028 3792 18040
rect 3844 18068 3850 18080
rect 4154 18068 4160 18080
rect 3844 18040 4160 18068
rect 3844 18028 3850 18040
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 7024 18077 7052 18108
rect 7374 18096 7380 18108
rect 7432 18096 7438 18148
rect 7009 18071 7067 18077
rect 7009 18037 7021 18071
rect 7055 18037 7067 18071
rect 7009 18031 7067 18037
rect 7282 18028 7288 18080
rect 7340 18028 7346 18080
rect 7469 18071 7527 18077
rect 7469 18037 7481 18071
rect 7515 18068 7527 18071
rect 7558 18068 7564 18080
rect 7515 18040 7564 18068
rect 7515 18037 7527 18040
rect 7469 18031 7527 18037
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 7852 18068 7880 18167
rect 7944 18136 7972 18167
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 9398 18164 9404 18216
rect 9456 18164 9462 18216
rect 10042 18164 10048 18216
rect 10100 18164 10106 18216
rect 9490 18136 9496 18148
rect 7944 18108 9496 18136
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 10152 18136 10180 18235
rect 10502 18164 10508 18216
rect 10560 18164 10566 18216
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18204 12403 18207
rect 12529 18207 12587 18213
rect 12529 18204 12541 18207
rect 12391 18176 12541 18204
rect 12391 18173 12403 18176
rect 12345 18167 12403 18173
rect 12529 18173 12541 18176
rect 12575 18173 12587 18207
rect 12529 18167 12587 18173
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 13630 18204 13636 18216
rect 12676 18176 13636 18204
rect 12676 18164 12682 18176
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 13725 18207 13783 18213
rect 13725 18173 13737 18207
rect 13771 18204 13783 18207
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 13771 18176 13921 18204
rect 13771 18173 13783 18176
rect 13725 18167 13783 18173
rect 13909 18173 13921 18176
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 14182 18164 14188 18216
rect 14240 18164 14246 18216
rect 15838 18164 15844 18216
rect 15896 18164 15902 18216
rect 15948 18213 15976 18380
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 17696 18380 17816 18408
rect 16577 18343 16635 18349
rect 16577 18309 16589 18343
rect 16623 18340 16635 18343
rect 16850 18340 16856 18352
rect 16623 18312 16856 18340
rect 16623 18309 16635 18312
rect 16577 18303 16635 18309
rect 16850 18300 16856 18312
rect 16908 18340 16914 18352
rect 17696 18340 17724 18380
rect 17788 18349 17816 18380
rect 17862 18368 17868 18420
rect 17920 18408 17926 18420
rect 20254 18408 20260 18420
rect 17920 18380 20260 18408
rect 17920 18368 17926 18380
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 20533 18411 20591 18417
rect 20533 18377 20545 18411
rect 20579 18408 20591 18411
rect 20714 18408 20720 18420
rect 20579 18380 20720 18408
rect 20579 18377 20591 18380
rect 20533 18371 20591 18377
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 22186 18408 22192 18420
rect 20916 18380 22192 18408
rect 16908 18312 17724 18340
rect 17773 18343 17831 18349
rect 16908 18300 16914 18312
rect 17773 18309 17785 18343
rect 17819 18309 17831 18343
rect 17773 18303 17831 18309
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 16132 18244 16313 18272
rect 16132 18213 16160 18244
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16448 18244 16681 18272
rect 16448 18232 16454 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 16669 18235 16727 18241
rect 16868 18244 17049 18272
rect 15933 18207 15991 18213
rect 15933 18173 15945 18207
rect 15979 18173 15991 18207
rect 15933 18167 15991 18173
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18173 16175 18207
rect 16117 18167 16175 18173
rect 16206 18164 16212 18216
rect 16264 18164 16270 18216
rect 16485 18207 16543 18213
rect 16485 18204 16497 18207
rect 16316 18176 16497 18204
rect 10870 18136 10876 18148
rect 10060 18108 10876 18136
rect 10060 18080 10088 18108
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 11606 18096 11612 18148
rect 11664 18136 11670 18148
rect 12078 18139 12136 18145
rect 12078 18136 12090 18139
rect 11664 18108 12090 18136
rect 11664 18096 11670 18108
rect 12078 18105 12090 18108
rect 12124 18105 12136 18139
rect 12078 18099 12136 18105
rect 15194 18096 15200 18148
rect 15252 18136 15258 18148
rect 15657 18139 15715 18145
rect 15657 18136 15669 18139
rect 15252 18108 15669 18136
rect 15252 18096 15258 18108
rect 15657 18105 15669 18108
rect 15703 18105 15715 18139
rect 16224 18136 16252 18164
rect 16316 18148 16344 18176
rect 16485 18173 16497 18176
rect 16531 18173 16543 18207
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 16485 18167 16543 18173
rect 16592 18176 16773 18204
rect 15657 18099 15715 18105
rect 15856 18108 16252 18136
rect 10042 18068 10048 18080
rect 7852 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 15856 18068 15884 18108
rect 16298 18096 16304 18148
rect 16356 18096 16362 18148
rect 16592 18136 16620 18176
rect 16761 18173 16773 18176
rect 16807 18173 16819 18207
rect 16868 18204 16896 18244
rect 17037 18241 17049 18244
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 17402 18232 17408 18284
rect 17460 18232 17466 18284
rect 17494 18232 17500 18284
rect 17552 18232 17558 18284
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 20916 18272 20944 18380
rect 22186 18368 22192 18380
rect 22244 18408 22250 18420
rect 22830 18408 22836 18420
rect 22244 18380 22836 18408
rect 22244 18368 22250 18380
rect 22830 18368 22836 18380
rect 22888 18368 22894 18420
rect 24026 18368 24032 18420
rect 24084 18408 24090 18420
rect 24121 18411 24179 18417
rect 24121 18408 24133 18411
rect 24084 18380 24133 18408
rect 24084 18368 24090 18380
rect 24121 18377 24133 18380
rect 24167 18377 24179 18411
rect 24121 18371 24179 18377
rect 26973 18411 27031 18417
rect 26973 18377 26985 18411
rect 27019 18408 27031 18411
rect 27706 18408 27712 18420
rect 27019 18380 27712 18408
rect 27019 18377 27031 18380
rect 26973 18371 27031 18377
rect 27706 18368 27712 18380
rect 27764 18368 27770 18420
rect 28074 18368 28080 18420
rect 28132 18368 28138 18420
rect 28813 18411 28871 18417
rect 28813 18377 28825 18411
rect 28859 18408 28871 18411
rect 29546 18408 29552 18420
rect 28859 18380 29552 18408
rect 28859 18377 28871 18380
rect 28813 18371 28871 18377
rect 29546 18368 29552 18380
rect 29604 18368 29610 18420
rect 30098 18368 30104 18420
rect 30156 18408 30162 18420
rect 30193 18411 30251 18417
rect 30193 18408 30205 18411
rect 30156 18380 30205 18408
rect 30156 18368 30162 18380
rect 30193 18377 30205 18380
rect 30239 18377 30251 18411
rect 30193 18371 30251 18377
rect 23290 18300 23296 18352
rect 23348 18340 23354 18352
rect 27614 18340 27620 18352
rect 23348 18312 27620 18340
rect 23348 18300 23354 18312
rect 18288 18244 20944 18272
rect 18288 18232 18294 18244
rect 17865 18217 17923 18223
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 16868 18176 16957 18204
rect 16761 18167 16819 18173
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17221 18207 17279 18213
rect 17221 18204 17233 18207
rect 17184 18176 17233 18204
rect 17184 18164 17190 18176
rect 17221 18173 17233 18176
rect 17267 18173 17279 18207
rect 17221 18167 17279 18173
rect 17313 18207 17371 18213
rect 17313 18173 17325 18207
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 17681 18207 17739 18213
rect 17681 18173 17693 18207
rect 17727 18173 17739 18207
rect 17865 18183 17877 18217
rect 17911 18214 17923 18217
rect 17911 18186 18000 18214
rect 17911 18183 17923 18186
rect 17865 18177 17923 18183
rect 17681 18167 17739 18173
rect 16500 18108 16620 18136
rect 15344 18040 15884 18068
rect 15344 18028 15350 18040
rect 15930 18028 15936 18080
rect 15988 18068 15994 18080
rect 16316 18068 16344 18096
rect 16500 18080 16528 18108
rect 15988 18040 16344 18068
rect 15988 18028 15994 18040
rect 16482 18028 16488 18080
rect 16540 18028 16546 18080
rect 17236 18068 17264 18167
rect 17328 18136 17356 18167
rect 17696 18136 17724 18167
rect 17862 18136 17868 18148
rect 17328 18108 17868 18136
rect 17862 18096 17868 18108
rect 17920 18096 17926 18148
rect 17972 18068 18000 18186
rect 19794 18164 19800 18216
rect 19852 18204 19858 18216
rect 19889 18207 19947 18213
rect 19889 18204 19901 18207
rect 19852 18176 19901 18204
rect 19852 18164 19858 18176
rect 19889 18173 19901 18176
rect 19935 18173 19947 18207
rect 19889 18167 19947 18173
rect 20070 18164 20076 18216
rect 20128 18164 20134 18216
rect 20438 18164 20444 18216
rect 20496 18164 20502 18216
rect 20640 18213 20668 18244
rect 20990 18232 20996 18284
rect 21048 18232 21054 18284
rect 21082 18232 21088 18284
rect 21140 18232 21146 18284
rect 21174 18232 21180 18284
rect 21232 18232 21238 18284
rect 25222 18272 25228 18284
rect 24596 18244 25228 18272
rect 20625 18207 20683 18213
rect 20625 18173 20637 18207
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 20901 18207 20959 18213
rect 20901 18173 20913 18207
rect 20947 18204 20959 18207
rect 21358 18204 21364 18216
rect 20947 18176 21364 18204
rect 20947 18173 20959 18176
rect 20901 18167 20959 18173
rect 18874 18096 18880 18148
rect 18932 18136 18938 18148
rect 19337 18139 19395 18145
rect 19337 18136 19349 18139
rect 18932 18108 19349 18136
rect 18932 18096 18938 18108
rect 19337 18105 19349 18108
rect 19383 18105 19395 18139
rect 19337 18099 19395 18105
rect 19521 18139 19579 18145
rect 19521 18105 19533 18139
rect 19567 18136 19579 18139
rect 20916 18136 20944 18167
rect 21358 18164 21364 18176
rect 21416 18164 21422 18216
rect 23014 18164 23020 18216
rect 23072 18204 23078 18216
rect 23477 18207 23535 18213
rect 23477 18204 23489 18207
rect 23072 18176 23489 18204
rect 23072 18164 23078 18176
rect 23477 18173 23489 18176
rect 23523 18173 23535 18207
rect 23477 18167 23535 18173
rect 24305 18207 24363 18213
rect 24305 18173 24317 18207
rect 24351 18173 24363 18207
rect 24305 18167 24363 18173
rect 24397 18207 24455 18213
rect 24397 18173 24409 18207
rect 24443 18204 24455 18207
rect 24486 18204 24492 18216
rect 24443 18176 24492 18204
rect 24443 18173 24455 18176
rect 24397 18167 24455 18173
rect 19567 18108 20944 18136
rect 19567 18105 19579 18108
rect 19521 18099 19579 18105
rect 23290 18096 23296 18148
rect 23348 18096 23354 18148
rect 24320 18136 24348 18167
rect 24486 18164 24492 18176
rect 24544 18164 24550 18216
rect 24596 18213 24624 18244
rect 25222 18232 25228 18244
rect 25280 18232 25286 18284
rect 25317 18275 25375 18281
rect 25317 18241 25329 18275
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 24581 18207 24639 18213
rect 24581 18173 24593 18207
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 24673 18207 24731 18213
rect 24673 18173 24685 18207
rect 24719 18204 24731 18207
rect 25038 18204 25044 18216
rect 24719 18176 25044 18204
rect 24719 18173 24731 18176
rect 24673 18167 24731 18173
rect 25038 18164 25044 18176
rect 25096 18164 25102 18216
rect 25130 18164 25136 18216
rect 25188 18204 25194 18216
rect 25332 18204 25360 18235
rect 25188 18176 25360 18204
rect 25700 18204 25728 18312
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 28350 18300 28356 18352
rect 28408 18340 28414 18352
rect 29086 18340 29092 18352
rect 28408 18312 29092 18340
rect 28408 18300 28414 18312
rect 29086 18300 29092 18312
rect 29144 18300 29150 18352
rect 29178 18300 29184 18352
rect 29236 18340 29242 18352
rect 29236 18312 29592 18340
rect 29236 18300 29242 18312
rect 29564 18284 29592 18312
rect 29365 18275 29423 18281
rect 29365 18272 29377 18275
rect 26620 18244 28120 18272
rect 26620 18216 26648 18244
rect 25869 18207 25927 18213
rect 25869 18204 25881 18207
rect 25700 18176 25881 18204
rect 25188 18164 25194 18176
rect 25869 18173 25881 18176
rect 25915 18173 25927 18207
rect 25869 18167 25927 18173
rect 26050 18164 26056 18216
rect 26108 18164 26114 18216
rect 26237 18207 26295 18213
rect 26237 18173 26249 18207
rect 26283 18204 26295 18207
rect 26329 18207 26387 18213
rect 26329 18204 26341 18207
rect 26283 18176 26341 18204
rect 26283 18173 26295 18176
rect 26237 18167 26295 18173
rect 26329 18173 26341 18176
rect 26375 18173 26387 18207
rect 26329 18167 26387 18173
rect 26513 18207 26571 18213
rect 26513 18173 26525 18207
rect 26559 18173 26571 18207
rect 26513 18167 26571 18173
rect 24320 18108 24808 18136
rect 17236 18040 18000 18068
rect 19429 18071 19487 18077
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 19610 18068 19616 18080
rect 19475 18040 19616 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 21361 18071 21419 18077
rect 21361 18068 21373 18071
rect 20956 18040 21373 18068
rect 20956 18028 20962 18040
rect 21361 18037 21373 18040
rect 21407 18037 21419 18071
rect 21361 18031 21419 18037
rect 23661 18071 23719 18077
rect 23661 18037 23673 18071
rect 23707 18068 23719 18071
rect 24578 18068 24584 18080
rect 23707 18040 24584 18068
rect 23707 18037 23719 18040
rect 23661 18031 23719 18037
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 24780 18077 24808 18108
rect 25148 18108 25820 18136
rect 24765 18071 24823 18077
rect 24765 18037 24777 18071
rect 24811 18037 24823 18071
rect 24765 18031 24823 18037
rect 24946 18028 24952 18080
rect 25004 18068 25010 18080
rect 25148 18077 25176 18108
rect 25133 18071 25191 18077
rect 25133 18068 25145 18071
rect 25004 18040 25145 18068
rect 25004 18028 25010 18040
rect 25133 18037 25145 18040
rect 25179 18037 25191 18071
rect 25133 18031 25191 18037
rect 25225 18071 25283 18077
rect 25225 18037 25237 18071
rect 25271 18068 25283 18071
rect 25314 18068 25320 18080
rect 25271 18040 25320 18068
rect 25271 18037 25283 18040
rect 25225 18031 25283 18037
rect 25314 18028 25320 18040
rect 25372 18028 25378 18080
rect 25792 18068 25820 18108
rect 26142 18096 26148 18148
rect 26200 18136 26206 18148
rect 26528 18136 26556 18167
rect 26602 18164 26608 18216
rect 26660 18164 26666 18216
rect 26697 18207 26755 18213
rect 26697 18173 26709 18207
rect 26743 18204 26755 18207
rect 26786 18204 26792 18216
rect 26743 18176 26792 18204
rect 26743 18173 26755 18176
rect 26697 18167 26755 18173
rect 26786 18164 26792 18176
rect 26844 18204 26850 18216
rect 26844 18176 28028 18204
rect 26844 18164 26850 18176
rect 27430 18136 27436 18148
rect 26200 18108 27436 18136
rect 26200 18096 26206 18108
rect 27430 18096 27436 18108
rect 27488 18096 27494 18148
rect 27614 18096 27620 18148
rect 27672 18136 27678 18148
rect 27709 18139 27767 18145
rect 27709 18136 27721 18139
rect 27672 18108 27721 18136
rect 27672 18096 27678 18108
rect 27709 18105 27721 18108
rect 27755 18105 27767 18139
rect 27709 18099 27767 18105
rect 27893 18139 27951 18145
rect 27893 18105 27905 18139
rect 27939 18105 27951 18139
rect 27893 18099 27951 18105
rect 27908 18068 27936 18099
rect 25792 18040 27936 18068
rect 28000 18068 28028 18176
rect 28092 18136 28120 18244
rect 28184 18244 29377 18272
rect 28184 18213 28212 18244
rect 29365 18241 29377 18244
rect 29411 18241 29423 18275
rect 29365 18235 29423 18241
rect 29546 18232 29552 18284
rect 29604 18232 29610 18284
rect 29638 18232 29644 18284
rect 29696 18272 29702 18284
rect 29733 18275 29791 18281
rect 29733 18272 29745 18275
rect 29696 18244 29745 18272
rect 29696 18232 29702 18244
rect 29733 18241 29745 18244
rect 29779 18241 29791 18275
rect 29733 18235 29791 18241
rect 28169 18207 28227 18213
rect 28169 18173 28181 18207
rect 28215 18173 28227 18207
rect 28169 18167 28227 18173
rect 28350 18164 28356 18216
rect 28408 18164 28414 18216
rect 28445 18207 28503 18213
rect 28445 18173 28457 18207
rect 28491 18173 28503 18207
rect 28445 18167 28503 18173
rect 28537 18207 28595 18213
rect 28537 18173 28549 18207
rect 28583 18204 28595 18207
rect 29454 18204 29460 18216
rect 28583 18176 29460 18204
rect 28583 18173 28595 18176
rect 28537 18167 28595 18173
rect 28460 18136 28488 18167
rect 29454 18164 29460 18176
rect 29512 18204 29518 18216
rect 29825 18207 29883 18213
rect 29825 18204 29837 18207
rect 29512 18176 29837 18204
rect 29512 18164 29518 18176
rect 29825 18173 29837 18176
rect 29871 18173 29883 18207
rect 29825 18167 29883 18173
rect 28626 18136 28632 18148
rect 28092 18108 28632 18136
rect 28626 18096 28632 18108
rect 28684 18096 28690 18148
rect 28902 18096 28908 18148
rect 28960 18136 28966 18148
rect 28997 18139 29055 18145
rect 28997 18136 29009 18139
rect 28960 18108 29009 18136
rect 28960 18096 28966 18108
rect 28997 18105 29009 18108
rect 29043 18105 29055 18139
rect 28997 18099 29055 18105
rect 29181 18139 29239 18145
rect 29181 18105 29193 18139
rect 29227 18136 29239 18139
rect 29638 18136 29644 18148
rect 29227 18108 29644 18136
rect 29227 18105 29239 18108
rect 29181 18099 29239 18105
rect 29196 18068 29224 18099
rect 29638 18096 29644 18108
rect 29696 18096 29702 18148
rect 28000 18040 29224 18068
rect 552 17978 31648 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 12096 17978
rect 12148 17926 12160 17978
rect 12212 17926 12224 17978
rect 12276 17926 12288 17978
rect 12340 17926 12352 17978
rect 12404 17926 19870 17978
rect 19922 17926 19934 17978
rect 19986 17926 19998 17978
rect 20050 17926 20062 17978
rect 20114 17926 20126 17978
rect 20178 17926 27644 17978
rect 27696 17926 27708 17978
rect 27760 17926 27772 17978
rect 27824 17926 27836 17978
rect 27888 17926 27900 17978
rect 27952 17926 31648 17978
rect 552 17904 31648 17926
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 3510 17864 3516 17876
rect 3375 17836 3516 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 4246 17824 4252 17876
rect 4304 17824 4310 17876
rect 7834 17864 7840 17876
rect 6748 17836 7840 17864
rect 2682 17756 2688 17808
rect 2740 17796 2746 17808
rect 2740 17768 4200 17796
rect 2740 17756 2746 17768
rect 1302 17688 1308 17740
rect 1360 17728 1366 17740
rect 2222 17737 2228 17740
rect 1949 17731 2007 17737
rect 1949 17728 1961 17731
rect 1360 17700 1961 17728
rect 1360 17688 1366 17700
rect 1949 17697 1961 17700
rect 1995 17697 2007 17731
rect 1949 17691 2007 17697
rect 2216 17691 2228 17737
rect 2222 17688 2228 17691
rect 2280 17688 2286 17740
rect 3510 17688 3516 17740
rect 3568 17728 3574 17740
rect 3605 17731 3663 17737
rect 3605 17728 3617 17731
rect 3568 17700 3617 17728
rect 3568 17688 3574 17700
rect 3605 17697 3617 17700
rect 3651 17697 3663 17731
rect 3605 17691 3663 17697
rect 3786 17688 3792 17740
rect 3844 17688 3850 17740
rect 4172 17737 4200 17768
rect 5810 17756 5816 17808
rect 5868 17756 5874 17808
rect 3881 17731 3939 17737
rect 3881 17697 3893 17731
rect 3927 17697 3939 17731
rect 3881 17691 3939 17697
rect 4157 17731 4215 17737
rect 4157 17697 4169 17731
rect 4203 17697 4215 17731
rect 4157 17691 4215 17697
rect 3896 17592 3924 17691
rect 4172 17660 4200 17691
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 5166 17728 5172 17740
rect 4304 17700 5172 17728
rect 4304 17688 4310 17700
rect 5166 17688 5172 17700
rect 5224 17728 5230 17740
rect 5997 17731 6055 17737
rect 5997 17728 6009 17731
rect 5224 17700 6009 17728
rect 5224 17688 5230 17700
rect 5997 17697 6009 17700
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 6086 17688 6092 17740
rect 6144 17688 6150 17740
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17697 6515 17731
rect 6457 17691 6515 17697
rect 4430 17660 4436 17672
rect 4172 17632 4436 17660
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 6472 17660 6500 17691
rect 6638 17688 6644 17740
rect 6696 17688 6702 17740
rect 6748 17737 6776 17836
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 9490 17824 9496 17876
rect 9548 17824 9554 17876
rect 10134 17824 10140 17876
rect 10192 17824 10198 17876
rect 10686 17824 10692 17876
rect 10744 17824 10750 17876
rect 11606 17824 11612 17876
rect 11664 17824 11670 17876
rect 13262 17824 13268 17876
rect 13320 17824 13326 17876
rect 14182 17824 14188 17876
rect 14240 17864 14246 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14240 17836 14657 17864
rect 14240 17824 14246 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 16117 17867 16175 17873
rect 16117 17864 16129 17867
rect 15804 17836 16129 17864
rect 15804 17824 15810 17836
rect 16117 17833 16129 17836
rect 16163 17833 16175 17867
rect 16117 17827 16175 17833
rect 16298 17824 16304 17876
rect 16356 17864 16362 17876
rect 17862 17864 17868 17876
rect 16356 17836 17868 17864
rect 16356 17824 16362 17836
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 25222 17824 25228 17876
rect 25280 17824 25286 17876
rect 28166 17824 28172 17876
rect 28224 17864 28230 17876
rect 28994 17864 29000 17876
rect 28224 17836 29000 17864
rect 28224 17824 28230 17836
rect 28994 17824 29000 17836
rect 29052 17824 29058 17876
rect 29270 17824 29276 17876
rect 29328 17824 29334 17876
rect 29362 17824 29368 17876
rect 29420 17824 29426 17876
rect 7374 17756 7380 17808
rect 7432 17796 7438 17808
rect 7432 17768 9674 17796
rect 7432 17756 7438 17768
rect 6733 17731 6791 17737
rect 6733 17697 6745 17731
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6822 17688 6828 17740
rect 6880 17688 6886 17740
rect 7282 17688 7288 17740
rect 7340 17688 7346 17740
rect 7558 17737 7564 17740
rect 7552 17728 7564 17737
rect 7519 17700 7564 17728
rect 7552 17691 7564 17700
rect 7558 17688 7564 17691
rect 7616 17688 7622 17740
rect 9646 17728 9674 17768
rect 10244 17768 10456 17796
rect 10244 17737 10272 17768
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9646 17700 9873 17728
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10229 17731 10287 17737
rect 10229 17697 10241 17731
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17697 10379 17731
rect 10321 17691 10379 17697
rect 6914 17660 6920 17672
rect 6472 17632 6920 17660
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 10336 17660 10364 17691
rect 9548 17632 10364 17660
rect 10428 17660 10456 17768
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 10928 17768 11284 17796
rect 10928 17756 10934 17768
rect 10502 17688 10508 17740
rect 10560 17688 10566 17740
rect 11256 17737 11284 17768
rect 11900 17768 12572 17796
rect 10965 17731 11023 17737
rect 10965 17697 10977 17731
rect 11011 17728 11023 17731
rect 11149 17731 11207 17737
rect 11011 17700 11100 17728
rect 11011 17697 11023 17700
rect 10965 17691 11023 17697
rect 11072 17672 11100 17700
rect 11149 17697 11161 17731
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17697 11299 17731
rect 11241 17691 11299 17697
rect 10428 17632 10548 17660
rect 9548 17620 9554 17632
rect 4706 17592 4712 17604
rect 3896 17564 4712 17592
rect 4706 17552 4712 17564
rect 4764 17552 4770 17604
rect 9953 17595 10011 17601
rect 8680 17564 9904 17592
rect 8680 17536 8708 17564
rect 3881 17527 3939 17533
rect 3881 17493 3893 17527
rect 3927 17524 3939 17527
rect 3970 17524 3976 17536
rect 3927 17496 3976 17524
rect 3927 17493 3939 17496
rect 3881 17487 3939 17493
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 4065 17527 4123 17533
rect 4065 17493 4077 17527
rect 4111 17524 4123 17527
rect 4154 17524 4160 17536
rect 4111 17496 4160 17524
rect 4111 17493 4123 17496
rect 4065 17487 4123 17493
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 6086 17484 6092 17536
rect 6144 17484 6150 17536
rect 7009 17527 7067 17533
rect 7009 17493 7021 17527
rect 7055 17524 7067 17527
rect 8386 17524 8392 17536
rect 7055 17496 8392 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 8662 17484 8668 17536
rect 8720 17484 8726 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 9769 17527 9827 17533
rect 9769 17524 9781 17527
rect 9732 17496 9781 17524
rect 9732 17484 9738 17496
rect 9769 17493 9781 17496
rect 9815 17493 9827 17527
rect 9876 17524 9904 17564
rect 9953 17561 9965 17595
rect 9999 17592 10011 17595
rect 9999 17564 10456 17592
rect 9999 17561 10011 17564
rect 9953 17555 10011 17561
rect 10428 17536 10456 17564
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 9876 17496 10333 17524
rect 9769 17487 9827 17493
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10321 17487 10379 17493
rect 10410 17484 10416 17536
rect 10468 17484 10474 17536
rect 10520 17524 10548 17632
rect 11054 17620 11060 17672
rect 11112 17620 11118 17672
rect 11173 17660 11201 17691
rect 11330 17688 11336 17740
rect 11388 17688 11394 17740
rect 11900 17672 11928 17768
rect 12544 17737 12572 17768
rect 12069 17731 12127 17737
rect 12069 17697 12081 17731
rect 12115 17728 12127 17731
rect 12345 17731 12403 17737
rect 12345 17728 12357 17731
rect 12115 17700 12357 17728
rect 12115 17697 12127 17700
rect 12069 17691 12127 17697
rect 12345 17697 12357 17700
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 12529 17731 12587 17737
rect 12529 17697 12541 17731
rect 12575 17697 12587 17731
rect 13280 17728 13308 17824
rect 13630 17756 13636 17808
rect 13688 17796 13694 17808
rect 16666 17796 16672 17808
rect 13688 17768 15792 17796
rect 13688 17756 13694 17768
rect 12529 17691 12587 17697
rect 12636 17700 13308 17728
rect 13541 17731 13599 17737
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11173 17632 11713 17660
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 11882 17620 11888 17672
rect 11940 17620 11946 17672
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17629 12219 17663
rect 12360 17660 12388 17691
rect 12636 17660 12664 17700
rect 13541 17697 13553 17731
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 12360 17632 12664 17660
rect 12161 17623 12219 17629
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 12176 17592 12204 17623
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 13556 17660 13584 17691
rect 13814 17688 13820 17740
rect 13872 17688 13878 17740
rect 14918 17688 14924 17740
rect 14976 17688 14982 17740
rect 15013 17731 15071 17737
rect 15013 17697 15025 17731
rect 15059 17697 15071 17731
rect 15013 17691 15071 17697
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15194 17728 15200 17740
rect 15151 17700 15200 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 13832 17660 13860 17688
rect 12860 17632 13584 17660
rect 13740 17632 13860 17660
rect 12860 17620 12866 17632
rect 11204 17564 12204 17592
rect 13173 17595 13231 17601
rect 11204 17552 11210 17564
rect 13173 17561 13185 17595
rect 13219 17592 13231 17595
rect 13740 17592 13768 17632
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 15028 17660 15056 17691
rect 15194 17688 15200 17700
rect 15252 17688 15258 17740
rect 15289 17731 15347 17737
rect 15289 17697 15301 17731
rect 15335 17728 15347 17731
rect 15378 17728 15384 17740
rect 15335 17700 15384 17728
rect 15335 17697 15347 17700
rect 15289 17691 15347 17697
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 15764 17737 15792 17768
rect 16500 17768 16672 17796
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 16390 17688 16396 17740
rect 16448 17688 16454 17740
rect 16500 17737 16528 17768
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 26326 17796 26332 17808
rect 24136 17768 26332 17796
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 16574 17688 16580 17740
rect 16632 17688 16638 17740
rect 16758 17688 16764 17740
rect 16816 17688 16822 17740
rect 17221 17731 17279 17737
rect 17221 17697 17233 17731
rect 17267 17728 17279 17731
rect 17310 17728 17316 17740
rect 17267 17700 17316 17728
rect 17267 17697 17279 17700
rect 17221 17691 17279 17697
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 20530 17688 20536 17740
rect 20588 17688 20594 17740
rect 20622 17688 20628 17740
rect 20680 17688 20686 17740
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17697 20775 17731
rect 20717 17691 20775 17697
rect 16206 17660 16212 17672
rect 14884 17632 16212 17660
rect 14884 17620 14890 17632
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 16408 17660 16436 17688
rect 16850 17660 16856 17672
rect 16408 17632 16856 17660
rect 16850 17620 16856 17632
rect 16908 17660 16914 17672
rect 17586 17660 17592 17672
rect 16908 17632 17592 17660
rect 16908 17620 16914 17632
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 20732 17660 20760 17691
rect 20898 17688 20904 17740
rect 20956 17688 20962 17740
rect 21910 17688 21916 17740
rect 21968 17688 21974 17740
rect 22186 17688 22192 17740
rect 22244 17688 22250 17740
rect 23201 17731 23259 17737
rect 23201 17697 23213 17731
rect 23247 17728 23259 17731
rect 23290 17728 23296 17740
rect 23247 17700 23296 17728
rect 23247 17697 23259 17700
rect 23201 17691 23259 17697
rect 23290 17688 23296 17700
rect 23348 17688 23354 17740
rect 23385 17731 23443 17737
rect 23385 17697 23397 17731
rect 23431 17728 23443 17731
rect 23474 17728 23480 17740
rect 23431 17700 23480 17728
rect 23431 17697 23443 17700
rect 23385 17691 23443 17697
rect 19306 17632 21496 17660
rect 13219 17564 13768 17592
rect 13817 17595 13875 17601
rect 13219 17561 13231 17564
rect 13173 17555 13231 17561
rect 13817 17561 13829 17595
rect 13863 17592 13875 17595
rect 15562 17592 15568 17604
rect 13863 17564 15568 17592
rect 13863 17561 13875 17564
rect 13817 17555 13875 17561
rect 12437 17527 12495 17533
rect 12437 17524 12449 17527
rect 10520 17496 12449 17524
rect 12437 17493 12449 17496
rect 12483 17493 12495 17527
rect 12437 17487 12495 17493
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 13832 17524 13860 17555
rect 15562 17552 15568 17564
rect 15620 17552 15626 17604
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 16758 17592 16764 17604
rect 16540 17564 16764 17592
rect 16540 17552 16546 17564
rect 16758 17552 16764 17564
rect 16816 17592 16822 17604
rect 17037 17595 17095 17601
rect 17037 17592 17049 17595
rect 16816 17564 17049 17592
rect 16816 17552 16822 17564
rect 17037 17561 17049 17564
rect 17083 17592 17095 17595
rect 19306 17592 19334 17632
rect 21468 17604 21496 17632
rect 21542 17620 21548 17672
rect 21600 17660 21606 17672
rect 22072 17663 22130 17669
rect 22072 17660 22084 17663
rect 21600 17632 22084 17660
rect 21600 17620 21606 17632
rect 22072 17629 22084 17632
rect 22118 17660 22130 17663
rect 22925 17663 22983 17669
rect 22118 17632 22600 17660
rect 22118 17629 22130 17632
rect 22072 17623 22130 17629
rect 17083 17564 19334 17592
rect 17083 17561 17095 17564
rect 17037 17555 17095 17561
rect 21266 17552 21272 17604
rect 21324 17552 21330 17604
rect 21450 17552 21456 17604
rect 21508 17552 21514 17604
rect 22462 17552 22468 17604
rect 22520 17552 22526 17604
rect 22572 17592 22600 17632
rect 22925 17629 22937 17663
rect 22971 17660 22983 17663
rect 23014 17660 23020 17672
rect 22971 17632 23020 17660
rect 22971 17629 22983 17632
rect 22925 17623 22983 17629
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 23106 17620 23112 17672
rect 23164 17620 23170 17672
rect 23400 17592 23428 17691
rect 23474 17688 23480 17700
rect 23532 17688 23538 17740
rect 24136 17660 24164 17768
rect 24210 17688 24216 17740
rect 24268 17728 24274 17740
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 24268 17700 24409 17728
rect 24268 17688 24274 17700
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 24489 17731 24547 17737
rect 24489 17697 24501 17731
rect 24535 17697 24547 17731
rect 24489 17691 24547 17697
rect 22572 17564 23428 17592
rect 23492 17632 24164 17660
rect 24504 17660 24532 17691
rect 24578 17688 24584 17740
rect 24636 17688 24642 17740
rect 24762 17688 24768 17740
rect 24820 17688 24826 17740
rect 24872 17737 24900 17768
rect 26326 17756 26332 17768
rect 26384 17796 26390 17808
rect 26602 17796 26608 17808
rect 26384 17768 26608 17796
rect 26384 17756 26390 17768
rect 26602 17756 26608 17768
rect 26660 17756 26666 17808
rect 28534 17796 28540 17808
rect 27816 17768 28540 17796
rect 27525 17753 27583 17759
rect 24857 17731 24915 17737
rect 24857 17697 24869 17731
rect 24903 17697 24915 17731
rect 24857 17691 24915 17697
rect 24946 17688 24952 17740
rect 25004 17688 25010 17740
rect 27525 17719 27537 17753
rect 27571 17719 27583 17753
rect 27816 17737 27844 17768
rect 28534 17756 28540 17768
rect 28592 17756 28598 17808
rect 29288 17796 29316 17824
rect 29288 17768 30512 17796
rect 27525 17713 27583 17719
rect 27617 17731 27675 17737
rect 27540 17672 27568 17713
rect 27617 17697 27629 17731
rect 27663 17697 27675 17731
rect 27617 17691 27675 17697
rect 27801 17731 27859 17737
rect 27801 17697 27813 17731
rect 27847 17697 27859 17731
rect 27801 17691 27859 17697
rect 27893 17731 27951 17737
rect 27893 17697 27905 17731
rect 27939 17728 27951 17731
rect 29273 17731 29331 17737
rect 27939 17700 28764 17728
rect 27939 17697 27951 17700
rect 27893 17691 27951 17697
rect 24504 17632 24900 17660
rect 12584 17496 13860 17524
rect 12584 17484 12590 17496
rect 15654 17484 15660 17536
rect 15712 17484 15718 17536
rect 20257 17527 20315 17533
rect 20257 17493 20269 17527
rect 20303 17524 20315 17527
rect 20438 17524 20444 17536
rect 20303 17496 20444 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 21468 17524 21496 17552
rect 22370 17524 22376 17536
rect 21468 17496 22376 17524
rect 22370 17484 22376 17496
rect 22428 17484 22434 17536
rect 23382 17484 23388 17536
rect 23440 17524 23446 17536
rect 23492 17524 23520 17632
rect 24872 17604 24900 17632
rect 27522 17620 27528 17672
rect 27580 17620 27586 17672
rect 27632 17660 27660 17691
rect 28626 17660 28632 17672
rect 27632 17632 28632 17660
rect 28626 17620 28632 17632
rect 28684 17620 28690 17672
rect 24854 17552 24860 17604
rect 24912 17552 24918 17604
rect 28077 17595 28135 17601
rect 28077 17561 28089 17595
rect 28123 17592 28135 17595
rect 28350 17592 28356 17604
rect 28123 17564 28356 17592
rect 28123 17561 28135 17564
rect 28077 17555 28135 17561
rect 28350 17552 28356 17564
rect 28408 17552 28414 17604
rect 28736 17592 28764 17700
rect 29273 17697 29285 17731
rect 29319 17697 29331 17731
rect 29273 17691 29331 17697
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17660 28871 17663
rect 29288 17660 29316 17691
rect 29546 17688 29552 17740
rect 29604 17728 29610 17740
rect 30484 17737 30512 17768
rect 30285 17731 30343 17737
rect 30285 17728 30297 17731
rect 29604 17700 30297 17728
rect 29604 17688 29610 17700
rect 30285 17697 30297 17700
rect 30331 17697 30343 17731
rect 30285 17691 30343 17697
rect 30469 17731 30527 17737
rect 30469 17697 30481 17731
rect 30515 17697 30527 17731
rect 30469 17691 30527 17697
rect 28859 17632 29316 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 28905 17595 28963 17601
rect 28905 17592 28917 17595
rect 28736 17564 28917 17592
rect 28905 17561 28917 17564
rect 28951 17561 28963 17595
rect 29288 17592 29316 17632
rect 29457 17663 29515 17669
rect 29457 17629 29469 17663
rect 29503 17660 29515 17663
rect 29638 17660 29644 17672
rect 29503 17632 29644 17660
rect 29503 17629 29515 17632
rect 29457 17623 29515 17629
rect 29638 17620 29644 17632
rect 29696 17620 29702 17672
rect 29546 17592 29552 17604
rect 29288 17564 29552 17592
rect 28905 17555 28963 17561
rect 29546 17552 29552 17564
rect 29604 17552 29610 17604
rect 23440 17496 23520 17524
rect 23440 17484 23446 17496
rect 23566 17484 23572 17536
rect 23624 17484 23630 17536
rect 23658 17484 23664 17536
rect 23716 17524 23722 17536
rect 24762 17524 24768 17536
rect 23716 17496 24768 17524
rect 23716 17484 23722 17496
rect 24762 17484 24768 17496
rect 24820 17524 24826 17536
rect 26234 17524 26240 17536
rect 24820 17496 26240 17524
rect 24820 17484 24826 17496
rect 26234 17484 26240 17496
rect 26292 17484 26298 17536
rect 27982 17484 27988 17536
rect 28040 17524 28046 17536
rect 28169 17527 28227 17533
rect 28169 17524 28181 17527
rect 28040 17496 28181 17524
rect 28040 17484 28046 17496
rect 28169 17493 28181 17496
rect 28215 17493 28227 17527
rect 28169 17487 28227 17493
rect 28994 17484 29000 17536
rect 29052 17524 29058 17536
rect 29733 17527 29791 17533
rect 29733 17524 29745 17527
rect 29052 17496 29745 17524
rect 29052 17484 29058 17496
rect 29733 17493 29745 17496
rect 29779 17493 29791 17527
rect 29733 17487 29791 17493
rect 30561 17527 30619 17533
rect 30561 17493 30573 17527
rect 30607 17524 30619 17527
rect 30650 17524 30656 17536
rect 30607 17496 30656 17524
rect 30607 17493 30619 17496
rect 30561 17487 30619 17493
rect 30650 17484 30656 17496
rect 30708 17484 30714 17536
rect 552 17434 31648 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 11436 17434
rect 11488 17382 11500 17434
rect 11552 17382 11564 17434
rect 11616 17382 11628 17434
rect 11680 17382 11692 17434
rect 11744 17382 19210 17434
rect 19262 17382 19274 17434
rect 19326 17382 19338 17434
rect 19390 17382 19402 17434
rect 19454 17382 19466 17434
rect 19518 17382 26984 17434
rect 27036 17382 27048 17434
rect 27100 17382 27112 17434
rect 27164 17382 27176 17434
rect 27228 17382 27240 17434
rect 27292 17382 31648 17434
rect 552 17360 31648 17382
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2409 17323 2467 17329
rect 2409 17320 2421 17323
rect 2280 17292 2421 17320
rect 2280 17280 2286 17292
rect 2409 17289 2421 17292
rect 2455 17289 2467 17323
rect 2409 17283 2467 17289
rect 2958 17280 2964 17332
rect 3016 17320 3022 17332
rect 3237 17323 3295 17329
rect 3237 17320 3249 17323
rect 3016 17292 3249 17320
rect 3016 17280 3022 17292
rect 3237 17289 3249 17292
rect 3283 17289 3295 17323
rect 3237 17283 3295 17289
rect 4341 17323 4399 17329
rect 4341 17289 4353 17323
rect 4387 17320 4399 17323
rect 6638 17320 6644 17332
rect 4387 17292 6644 17320
rect 4387 17289 4399 17292
rect 4341 17283 4399 17289
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7469 17323 7527 17329
rect 7469 17320 7481 17323
rect 6972 17292 7481 17320
rect 6972 17280 6978 17292
rect 7469 17289 7481 17292
rect 7515 17289 7527 17323
rect 7469 17283 7527 17289
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 7742 17320 7748 17332
rect 7699 17292 7748 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 7742 17280 7748 17292
rect 7800 17320 7806 17332
rect 8662 17320 8668 17332
rect 7800 17292 8668 17320
rect 7800 17280 7806 17292
rect 3050 17212 3056 17264
rect 3108 17212 3114 17264
rect 3697 17255 3755 17261
rect 3697 17221 3709 17255
rect 3743 17221 3755 17255
rect 3697 17215 3755 17221
rect 2682 17076 2688 17128
rect 2740 17076 2746 17128
rect 2774 17076 2780 17128
rect 2832 17076 2838 17128
rect 2866 17076 2872 17128
rect 2924 17076 2930 17128
rect 3068 17125 3096 17212
rect 3712 17184 3740 17215
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 7929 17255 7987 17261
rect 7929 17252 7941 17255
rect 6880 17224 7941 17252
rect 6880 17212 6886 17224
rect 7929 17221 7941 17224
rect 7975 17221 7987 17255
rect 7929 17215 7987 17221
rect 3712 17156 4384 17184
rect 3053 17119 3111 17125
rect 3053 17085 3065 17119
rect 3099 17085 3111 17119
rect 3053 17079 3111 17085
rect 3068 16980 3096 17079
rect 3142 17076 3148 17128
rect 3200 17116 3206 17128
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 3200 17088 3433 17116
rect 3200 17076 3206 17088
rect 3421 17085 3433 17088
rect 3467 17085 3479 17119
rect 3421 17079 3479 17085
rect 3513 17119 3571 17125
rect 3513 17085 3525 17119
rect 3559 17085 3571 17119
rect 3513 17079 3571 17085
rect 3234 17008 3240 17060
rect 3292 17008 3298 17060
rect 3326 17008 3332 17060
rect 3384 17048 3390 17060
rect 3528 17048 3556 17079
rect 4154 17076 4160 17128
rect 4212 17076 4218 17128
rect 4356 17125 4384 17156
rect 4430 17144 4436 17196
rect 4488 17184 4494 17196
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 4488 17156 6561 17184
rect 4488 17144 4494 17156
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17085 4399 17119
rect 4341 17079 4399 17085
rect 7926 17076 7932 17128
rect 7984 17076 7990 17128
rect 8128 17125 8156 17292
rect 8662 17280 8668 17292
rect 8720 17280 8726 17332
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 10502 17320 10508 17332
rect 10192 17292 10508 17320
rect 10192 17280 10198 17292
rect 10502 17280 10508 17292
rect 10560 17320 10566 17332
rect 11330 17320 11336 17332
rect 10560 17292 11336 17320
rect 10560 17280 10566 17292
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12618 17320 12624 17332
rect 12032 17292 12624 17320
rect 12032 17280 12038 17292
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 16666 17320 16672 17332
rect 15396 17292 16672 17320
rect 10962 17252 10968 17264
rect 10244 17224 10968 17252
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17116 8171 17119
rect 8202 17116 8208 17128
rect 8159 17088 8208 17116
rect 8159 17085 8171 17088
rect 8113 17079 8171 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 8570 17076 8576 17128
rect 8628 17116 8634 17128
rect 9582 17116 9588 17128
rect 8628 17088 9588 17116
rect 8628 17076 8634 17088
rect 9582 17076 9588 17088
rect 9640 17116 9646 17128
rect 10045 17119 10103 17125
rect 10045 17116 10057 17119
rect 9640 17088 10057 17116
rect 9640 17076 9646 17088
rect 10045 17085 10057 17088
rect 10091 17085 10103 17119
rect 10045 17079 10103 17085
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 10244 17116 10272 17224
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 15286 17252 15292 17264
rect 15120 17224 15292 17252
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10336 17156 10609 17184
rect 10336 17125 10364 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 12713 17187 12771 17193
rect 12713 17184 12725 17187
rect 11848 17156 12725 17184
rect 11848 17144 11854 17156
rect 12713 17153 12725 17156
rect 12759 17153 12771 17187
rect 13170 17184 13176 17196
rect 12713 17147 12771 17153
rect 13004 17156 13176 17184
rect 10183 17088 10272 17116
rect 10321 17119 10379 17125
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 10321 17085 10333 17119
rect 10367 17085 10379 17119
rect 10321 17079 10379 17085
rect 10410 17076 10416 17128
rect 10468 17076 10474 17128
rect 10686 17076 10692 17128
rect 10744 17076 10750 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 11112 17088 12449 17116
rect 11112 17076 11118 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12526 17076 12532 17128
rect 12584 17076 12590 17128
rect 12618 17076 12624 17128
rect 12676 17076 12682 17128
rect 13004 17125 13032 17156
rect 13170 17144 13176 17156
rect 13228 17184 13234 17196
rect 13630 17184 13636 17196
rect 13228 17156 13636 17184
rect 13228 17144 13234 17156
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 15120 17184 15148 17224
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 15396 17184 15424 17292
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 16853 17323 16911 17329
rect 16853 17289 16865 17323
rect 16899 17320 16911 17323
rect 16942 17320 16948 17332
rect 16899 17292 16948 17320
rect 16899 17289 16911 17292
rect 16853 17283 16911 17289
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 24118 17320 24124 17332
rect 21039 17292 24124 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 18046 17212 18052 17264
rect 18104 17252 18110 17264
rect 19242 17252 19248 17264
rect 18104 17224 19248 17252
rect 18104 17212 18110 17224
rect 19242 17212 19248 17224
rect 19300 17252 19306 17264
rect 19794 17252 19800 17264
rect 19300 17224 19800 17252
rect 19300 17212 19306 17224
rect 19794 17212 19800 17224
rect 19852 17212 19858 17264
rect 20438 17212 20444 17264
rect 20496 17212 20502 17264
rect 20530 17212 20536 17264
rect 20588 17252 20594 17264
rect 21269 17255 21327 17261
rect 21269 17252 21281 17255
rect 20588 17224 21281 17252
rect 20588 17212 20594 17224
rect 21269 17221 21281 17224
rect 21315 17252 21327 17255
rect 21542 17252 21548 17264
rect 21315 17224 21548 17252
rect 21315 17221 21327 17224
rect 21269 17215 21327 17221
rect 21542 17212 21548 17224
rect 21600 17212 21606 17264
rect 15654 17184 15660 17196
rect 15028 17156 15148 17184
rect 15304 17156 15424 17184
rect 15580 17156 15660 17184
rect 15028 17125 15056 17156
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17085 13047 17119
rect 12989 17079 13047 17085
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 15102 17076 15108 17128
rect 15160 17076 15166 17128
rect 15194 17076 15200 17128
rect 15252 17076 15258 17128
rect 15304 17113 15332 17156
rect 15381 17119 15439 17125
rect 15381 17113 15393 17119
rect 15304 17085 15393 17113
rect 15427 17085 15439 17119
rect 15381 17079 15439 17085
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 15580 17116 15608 17156
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 17402 17144 17408 17196
rect 17460 17184 17466 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17460 17156 17785 17184
rect 17460 17144 17466 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 20456 17184 20484 17212
rect 21634 17184 21640 17196
rect 20456 17156 20576 17184
rect 17773 17147 17831 17153
rect 15519 17088 15608 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 15746 17076 15752 17128
rect 15804 17076 15810 17128
rect 16942 17076 16948 17128
rect 17000 17116 17006 17128
rect 17681 17119 17739 17125
rect 17681 17116 17693 17119
rect 17000 17088 17693 17116
rect 17000 17076 17006 17088
rect 17681 17085 17693 17088
rect 17727 17085 17739 17119
rect 17681 17079 17739 17085
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 19852 17088 20177 17116
rect 19852 17076 19858 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 20349 17119 20407 17125
rect 20349 17085 20361 17119
rect 20395 17085 20407 17119
rect 20349 17079 20407 17085
rect 3384 17020 3556 17048
rect 3384 17008 3390 17020
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 7432 17020 7788 17048
rect 7432 17008 7438 17020
rect 3418 16980 3424 16992
rect 3068 16952 3424 16980
rect 3418 16940 3424 16952
rect 3476 16940 3482 16992
rect 7650 16989 7656 16992
rect 7637 16983 7656 16989
rect 7637 16949 7649 16983
rect 7637 16943 7656 16949
rect 7650 16940 7656 16943
rect 7708 16940 7714 16992
rect 7760 16980 7788 17020
rect 7834 17008 7840 17060
rect 7892 17008 7898 17060
rect 14461 17051 14519 17057
rect 14461 17048 14473 17051
rect 7944 17020 14473 17048
rect 7944 16980 7972 17020
rect 13004 16992 13032 17020
rect 14461 17017 14473 17020
rect 14507 17048 14519 17051
rect 20364 17048 20392 17079
rect 20438 17076 20444 17128
rect 20496 17076 20502 17128
rect 20548 17125 20576 17156
rect 20640 17156 21640 17184
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 20640 17048 20668 17156
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 22646 17144 22652 17196
rect 22704 17144 22710 17196
rect 22940 17184 22968 17292
rect 24118 17280 24124 17292
rect 24176 17280 24182 17332
rect 24394 17280 24400 17332
rect 24452 17320 24458 17332
rect 25130 17320 25136 17332
rect 24452 17292 25136 17320
rect 24452 17280 24458 17292
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 27430 17280 27436 17332
rect 27488 17320 27494 17332
rect 28166 17320 28172 17332
rect 27488 17292 28172 17320
rect 27488 17280 27494 17292
rect 28166 17280 28172 17292
rect 28224 17280 28230 17332
rect 28534 17280 28540 17332
rect 28592 17320 28598 17332
rect 29273 17323 29331 17329
rect 28592 17292 29224 17320
rect 28592 17280 28598 17292
rect 23106 17212 23112 17264
rect 23164 17252 23170 17264
rect 23164 17224 24992 17252
rect 23164 17212 23170 17224
rect 22940 17156 23060 17184
rect 20714 17076 20720 17128
rect 20772 17076 20778 17128
rect 21177 17119 21235 17125
rect 21177 17085 21189 17119
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 14507 17020 15608 17048
rect 20364 17020 20668 17048
rect 14507 17017 14519 17020
rect 14461 17011 14519 17017
rect 7760 16952 7972 16980
rect 9858 16940 9864 16992
rect 9916 16940 9922 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12897 16983 12955 16989
rect 12897 16980 12909 16983
rect 12584 16952 12909 16980
rect 12584 16940 12590 16952
rect 12897 16949 12909 16952
rect 12943 16949 12955 16983
rect 12897 16943 12955 16949
rect 12986 16940 12992 16992
rect 13044 16940 13050 16992
rect 14737 16983 14795 16989
rect 14737 16949 14749 16983
rect 14783 16980 14795 16983
rect 15470 16980 15476 16992
rect 14783 16952 15476 16980
rect 14783 16949 14795 16952
rect 14737 16943 14795 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15580 16980 15608 17020
rect 16574 16980 16580 16992
rect 15580 16952 16580 16980
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 17218 16940 17224 16992
rect 17276 16940 17282 16992
rect 17586 16940 17592 16992
rect 17644 16940 17650 16992
rect 19610 16940 19616 16992
rect 19668 16980 19674 16992
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 19668 16952 19993 16980
rect 19668 16940 19674 16952
rect 19981 16949 19993 16952
rect 20027 16949 20039 16983
rect 20732 16980 20760 17076
rect 21192 17048 21220 17079
rect 21818 17076 21824 17128
rect 21876 17116 21882 17128
rect 22741 17119 22799 17125
rect 22741 17116 22753 17119
rect 21876 17088 22753 17116
rect 21876 17076 21882 17088
rect 22741 17085 22753 17088
rect 22787 17085 22799 17119
rect 22741 17079 22799 17085
rect 22922 17076 22928 17128
rect 22980 17076 22986 17128
rect 23032 17125 23060 17156
rect 23198 17144 23204 17196
rect 23256 17184 23262 17196
rect 23569 17187 23627 17193
rect 23569 17184 23581 17187
rect 23256 17156 23581 17184
rect 23256 17144 23262 17156
rect 23569 17153 23581 17156
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 24394 17144 24400 17196
rect 24452 17144 24458 17196
rect 23017 17119 23075 17125
rect 23017 17085 23029 17119
rect 23063 17085 23075 17119
rect 23017 17079 23075 17085
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17116 23167 17119
rect 23474 17116 23480 17128
rect 23155 17088 23480 17116
rect 23155 17085 23167 17088
rect 23109 17079 23167 17085
rect 23474 17076 23480 17088
rect 23532 17076 23538 17128
rect 23661 17119 23719 17125
rect 23661 17085 23673 17119
rect 23707 17116 23719 17119
rect 24854 17116 24860 17128
rect 23707 17088 24860 17116
rect 23707 17085 23719 17088
rect 23661 17079 23719 17085
rect 24854 17076 24860 17088
rect 24912 17076 24918 17128
rect 24964 17125 24992 17224
rect 27614 17212 27620 17264
rect 27672 17252 27678 17264
rect 28258 17252 28264 17264
rect 27672 17224 28264 17252
rect 27672 17212 27678 17224
rect 28258 17212 28264 17224
rect 28316 17252 28322 17264
rect 28902 17252 28908 17264
rect 28316 17224 28908 17252
rect 28316 17212 28322 17224
rect 28902 17212 28908 17224
rect 28960 17212 28966 17264
rect 29196 17252 29224 17292
rect 29273 17289 29285 17323
rect 29319 17320 29331 17323
rect 29454 17320 29460 17332
rect 29319 17292 29460 17320
rect 29319 17289 29331 17292
rect 29273 17283 29331 17289
rect 29454 17280 29460 17292
rect 29512 17280 29518 17332
rect 30742 17320 30748 17332
rect 29748 17292 30748 17320
rect 29748 17252 29776 17292
rect 30742 17280 30748 17292
rect 30800 17280 30806 17332
rect 29196 17224 29776 17252
rect 25406 17144 25412 17196
rect 25464 17144 25470 17196
rect 25590 17144 25596 17196
rect 25648 17184 25654 17196
rect 29362 17184 29368 17196
rect 25648 17156 26464 17184
rect 25648 17144 25654 17156
rect 24949 17119 25007 17125
rect 24949 17085 24961 17119
rect 24995 17085 25007 17119
rect 24949 17079 25007 17085
rect 25133 17119 25191 17125
rect 25133 17085 25145 17119
rect 25179 17116 25191 17119
rect 26053 17119 26111 17125
rect 26053 17116 26065 17119
rect 25179 17088 26065 17116
rect 25179 17085 25191 17088
rect 25133 17079 25191 17085
rect 26053 17085 26065 17088
rect 26099 17085 26111 17119
rect 26053 17079 26111 17085
rect 22404 17051 22462 17057
rect 21192 17020 22094 17048
rect 21726 16980 21732 16992
rect 20732 16952 21732 16980
rect 19981 16943 20039 16949
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 22066 16980 22094 17020
rect 22404 17017 22416 17051
rect 22450 17048 22462 17051
rect 23385 17051 23443 17057
rect 23385 17048 23397 17051
rect 22450 17020 23397 17048
rect 22450 17017 22462 17020
rect 22404 17011 22462 17017
rect 23385 17017 23397 17020
rect 23431 17017 23443 17051
rect 23492 17048 23520 17076
rect 24305 17051 24363 17057
rect 24305 17048 24317 17051
rect 23492 17020 24317 17048
rect 23385 17011 23443 17017
rect 24305 17017 24317 17020
rect 24351 17017 24363 17051
rect 24305 17011 24363 17017
rect 24578 17008 24584 17060
rect 24636 17048 24642 17060
rect 24765 17051 24823 17057
rect 24765 17048 24777 17051
rect 24636 17020 24777 17048
rect 24636 17008 24642 17020
rect 24765 17017 24777 17020
rect 24811 17017 24823 17051
rect 24964 17048 24992 17079
rect 26234 17076 26240 17128
rect 26292 17076 26298 17128
rect 26326 17076 26332 17128
rect 26384 17076 26390 17128
rect 26436 17125 26464 17156
rect 27908 17156 29368 17184
rect 27908 17125 27936 17156
rect 29362 17144 29368 17156
rect 29420 17144 29426 17196
rect 30650 17144 30656 17196
rect 30708 17144 30714 17196
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 27893 17119 27951 17125
rect 27893 17085 27905 17119
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 28166 17076 28172 17128
rect 28224 17076 28230 17128
rect 28350 17076 28356 17128
rect 28408 17076 28414 17128
rect 28445 17119 28503 17125
rect 28445 17085 28457 17119
rect 28491 17085 28503 17119
rect 28445 17079 28503 17085
rect 28537 17119 28595 17125
rect 28537 17085 28549 17119
rect 28583 17116 28595 17119
rect 28994 17116 29000 17128
rect 28583 17088 29000 17116
rect 28583 17085 28595 17088
rect 28537 17079 28595 17085
rect 25498 17048 25504 17060
rect 24964 17020 25504 17048
rect 24765 17011 24823 17017
rect 25498 17008 25504 17020
rect 25556 17008 25562 17060
rect 25590 17008 25596 17060
rect 25648 17008 25654 17060
rect 25866 17008 25872 17060
rect 25924 17048 25930 17060
rect 26697 17051 26755 17057
rect 26697 17048 26709 17051
rect 25924 17020 26709 17048
rect 25924 17008 25930 17020
rect 26697 17017 26709 17020
rect 26743 17017 26755 17051
rect 26697 17011 26755 17017
rect 27614 17008 27620 17060
rect 27672 17048 27678 17060
rect 27709 17051 27767 17057
rect 27709 17048 27721 17051
rect 27672 17020 27721 17048
rect 27672 17008 27678 17020
rect 27709 17017 27721 17020
rect 27755 17017 27767 17051
rect 28460 17048 28488 17079
rect 28994 17076 29000 17088
rect 29052 17076 29058 17128
rect 29181 17119 29239 17125
rect 29181 17085 29193 17119
rect 29227 17116 29239 17119
rect 31018 17116 31024 17128
rect 29227 17088 31024 17116
rect 29227 17085 29239 17088
rect 29181 17079 29239 17085
rect 31018 17076 31024 17088
rect 31076 17076 31082 17128
rect 27709 17011 27767 17017
rect 28000 17020 28488 17048
rect 28813 17051 28871 17057
rect 22554 16980 22560 16992
rect 22066 16952 22560 16980
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 22646 16940 22652 16992
rect 22704 16980 22710 16992
rect 23198 16980 23204 16992
rect 22704 16952 23204 16980
rect 22704 16940 22710 16952
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 23474 16940 23480 16992
rect 23532 16980 23538 16992
rect 23845 16983 23903 16989
rect 23845 16980 23857 16983
rect 23532 16952 23857 16980
rect 23532 16940 23538 16952
rect 23845 16949 23857 16952
rect 23891 16949 23903 16983
rect 23845 16943 23903 16949
rect 23934 16940 23940 16992
rect 23992 16980 23998 16992
rect 24213 16983 24271 16989
rect 24213 16980 24225 16983
rect 23992 16952 24225 16980
rect 23992 16940 23998 16952
rect 24213 16949 24225 16952
rect 24259 16980 24271 16983
rect 25222 16980 25228 16992
rect 24259 16952 25228 16980
rect 24259 16949 24271 16952
rect 24213 16943 24271 16949
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 25961 16983 26019 16989
rect 25961 16949 25973 16983
rect 26007 16980 26019 16983
rect 26050 16980 26056 16992
rect 26007 16952 26056 16980
rect 26007 16949 26019 16952
rect 25961 16943 26019 16949
rect 26050 16940 26056 16952
rect 26108 16940 26114 16992
rect 26878 16940 26884 16992
rect 26936 16980 26942 16992
rect 28000 16980 28028 17020
rect 28813 17017 28825 17051
rect 28859 17048 28871 17051
rect 30386 17051 30444 17057
rect 30386 17048 30398 17051
rect 28859 17020 30398 17048
rect 28859 17017 28871 17020
rect 28813 17011 28871 17017
rect 30386 17017 30398 17020
rect 30432 17017 30444 17051
rect 30386 17011 30444 17017
rect 26936 16952 28028 16980
rect 28077 16983 28135 16989
rect 26936 16940 26942 16952
rect 28077 16949 28089 16983
rect 28123 16980 28135 16983
rect 28166 16980 28172 16992
rect 28123 16952 28172 16980
rect 28123 16949 28135 16952
rect 28077 16943 28135 16949
rect 28166 16940 28172 16952
rect 28224 16940 28230 16992
rect 29086 16940 29092 16992
rect 29144 16940 29150 16992
rect 552 16890 31648 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 12096 16890
rect 12148 16838 12160 16890
rect 12212 16838 12224 16890
rect 12276 16838 12288 16890
rect 12340 16838 12352 16890
rect 12404 16838 19870 16890
rect 19922 16838 19934 16890
rect 19986 16838 19998 16890
rect 20050 16838 20062 16890
rect 20114 16838 20126 16890
rect 20178 16838 27644 16890
rect 27696 16838 27708 16890
rect 27760 16838 27772 16890
rect 27824 16838 27836 16890
rect 27888 16838 27900 16890
rect 27952 16838 31648 16890
rect 552 16816 31648 16838
rect 2225 16779 2283 16785
rect 2225 16745 2237 16779
rect 2271 16776 2283 16779
rect 3142 16776 3148 16788
rect 2271 16748 3148 16776
rect 2271 16745 2283 16748
rect 2225 16739 2283 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 4893 16779 4951 16785
rect 4893 16745 4905 16779
rect 4939 16776 4951 16779
rect 6178 16776 6184 16788
rect 4939 16748 6184 16776
rect 4939 16745 4951 16748
rect 4893 16739 4951 16745
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 8570 16776 8576 16788
rect 7708 16748 8576 16776
rect 7708 16736 7714 16748
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 15194 16736 15200 16788
rect 15252 16776 15258 16788
rect 15565 16779 15623 16785
rect 15565 16776 15577 16779
rect 15252 16748 15577 16776
rect 15252 16736 15258 16748
rect 15565 16745 15577 16748
rect 15611 16745 15623 16779
rect 15565 16739 15623 16745
rect 16117 16779 16175 16785
rect 16117 16745 16129 16779
rect 16163 16745 16175 16779
rect 16117 16739 16175 16745
rect 1854 16668 1860 16720
rect 1912 16708 1918 16720
rect 2041 16711 2099 16717
rect 1912 16680 1992 16708
rect 1912 16668 1918 16680
rect 1578 16600 1584 16652
rect 1636 16600 1642 16652
rect 1964 16572 1992 16680
rect 2041 16677 2053 16711
rect 2087 16708 2099 16711
rect 2317 16711 2375 16717
rect 2317 16708 2329 16711
rect 2087 16680 2329 16708
rect 2087 16677 2099 16680
rect 2041 16671 2099 16677
rect 2317 16677 2329 16680
rect 2363 16677 2375 16711
rect 2317 16671 2375 16677
rect 6273 16711 6331 16717
rect 6273 16677 6285 16711
rect 6319 16708 6331 16711
rect 7374 16708 7380 16720
rect 6319 16680 7380 16708
rect 6319 16677 6331 16680
rect 6273 16671 6331 16677
rect 7374 16668 7380 16680
rect 7432 16668 7438 16720
rect 8389 16711 8447 16717
rect 8389 16677 8401 16711
rect 8435 16708 8447 16711
rect 9950 16708 9956 16720
rect 8435 16680 9956 16708
rect 8435 16677 8447 16680
rect 8389 16671 8447 16677
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 10042 16668 10048 16720
rect 10100 16708 10106 16720
rect 13633 16711 13691 16717
rect 13633 16708 13645 16711
rect 10100 16680 10548 16708
rect 10100 16668 10106 16680
rect 3050 16600 3056 16652
rect 3108 16600 3114 16652
rect 3234 16600 3240 16652
rect 3292 16600 3298 16652
rect 4246 16600 4252 16652
rect 4304 16600 4310 16652
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 6236 16612 7113 16640
rect 6236 16600 6242 16612
rect 7101 16609 7113 16612
rect 7147 16640 7159 16643
rect 7285 16643 7343 16649
rect 7285 16640 7297 16643
rect 7147 16612 7297 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 7285 16609 7297 16612
rect 7331 16609 7343 16643
rect 7285 16603 7343 16609
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 8202 16640 8208 16652
rect 7892 16612 8208 16640
rect 7892 16600 7898 16612
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8478 16600 8484 16652
rect 8536 16600 8542 16652
rect 8665 16643 8723 16649
rect 8665 16609 8677 16643
rect 8711 16640 8723 16643
rect 9030 16640 9036 16652
rect 8711 16612 9036 16640
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9490 16600 9496 16652
rect 9548 16600 9554 16652
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10318 16640 10324 16652
rect 9723 16612 10324 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10520 16649 10548 16680
rect 12820 16680 13645 16708
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 10686 16640 10692 16652
rect 10551 16612 10692 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 10686 16600 10692 16612
rect 10744 16600 10750 16652
rect 12820 16649 12848 16680
rect 13633 16677 13645 16680
rect 13679 16708 13691 16711
rect 14642 16708 14648 16720
rect 13679 16680 14648 16708
rect 13679 16677 13691 16680
rect 13633 16671 13691 16677
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 15102 16668 15108 16720
rect 15160 16708 15166 16720
rect 16132 16708 16160 16739
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16485 16779 16543 16785
rect 16485 16776 16497 16779
rect 16356 16748 16497 16776
rect 16356 16736 16362 16748
rect 16485 16745 16497 16748
rect 16531 16745 16543 16779
rect 16485 16739 16543 16745
rect 16577 16779 16635 16785
rect 16577 16745 16589 16779
rect 16623 16776 16635 16779
rect 17218 16776 17224 16788
rect 16623 16748 17224 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17402 16736 17408 16788
rect 17460 16736 17466 16788
rect 17586 16736 17592 16788
rect 17644 16776 17650 16788
rect 18509 16779 18567 16785
rect 18509 16776 18521 16779
rect 17644 16748 18521 16776
rect 17644 16736 17650 16748
rect 18509 16745 18521 16748
rect 18555 16745 18567 16779
rect 18509 16739 18567 16745
rect 18708 16748 22140 16776
rect 18708 16720 18736 16748
rect 16942 16708 16948 16720
rect 15160 16680 16160 16708
rect 16408 16680 16948 16708
rect 15160 16668 15166 16680
rect 12805 16643 12863 16649
rect 12805 16609 12817 16643
rect 12851 16609 12863 16643
rect 12805 16603 12863 16609
rect 12897 16643 12955 16649
rect 12897 16609 12909 16643
rect 12943 16640 12955 16643
rect 12986 16640 12992 16652
rect 12943 16612 12992 16640
rect 12943 16609 12955 16612
rect 12897 16603 12955 16609
rect 12986 16600 12992 16612
rect 13044 16600 13050 16652
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 15933 16643 15991 16649
rect 15795 16612 15884 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 2406 16572 2412 16584
rect 1964 16544 2412 16572
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 2958 16532 2964 16584
rect 3016 16532 3022 16584
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 3973 16575 4031 16581
rect 3973 16572 3985 16575
rect 3384 16544 3985 16572
rect 3384 16532 3390 16544
rect 3973 16541 3985 16544
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 4062 16532 4068 16584
rect 4120 16581 4126 16584
rect 4120 16575 4148 16581
rect 4136 16541 4148 16575
rect 4120 16535 4148 16541
rect 4120 16532 4126 16535
rect 8018 16532 8024 16584
rect 8076 16532 8082 16584
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 3697 16507 3755 16513
rect 3697 16473 3709 16507
rect 3743 16473 3755 16507
rect 3697 16467 3755 16473
rect 1670 16396 1676 16448
rect 1728 16396 1734 16448
rect 3712 16436 3740 16467
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 8128 16504 8156 16535
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 8444 16544 9873 16572
rect 8444 16532 8450 16544
rect 9861 16541 9873 16544
rect 9907 16572 9919 16575
rect 10042 16572 10048 16584
rect 9907 16544 10048 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16572 10287 16575
rect 11054 16572 11060 16584
rect 10275 16544 11060 16572
rect 10275 16541 10287 16544
rect 10229 16535 10287 16541
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 15654 16572 15660 16584
rect 12406 16544 15660 16572
rect 8202 16504 8208 16516
rect 7800 16476 8208 16504
rect 7800 16464 7806 16476
rect 8202 16464 8208 16476
rect 8260 16464 8266 16516
rect 10413 16507 10471 16513
rect 10413 16504 10425 16507
rect 9784 16476 10425 16504
rect 9784 16448 9812 16476
rect 10413 16473 10425 16476
rect 10459 16473 10471 16507
rect 10413 16467 10471 16473
rect 10502 16464 10508 16516
rect 10560 16504 10566 16516
rect 12406 16504 12434 16544
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 15856 16572 15884 16612
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16206 16640 16212 16652
rect 15979 16612 16212 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 16408 16640 16436 16680
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 18138 16708 18144 16720
rect 17144 16680 18144 16708
rect 17144 16649 17172 16680
rect 18138 16668 18144 16680
rect 18196 16708 18202 16720
rect 18690 16708 18696 16720
rect 18196 16680 18696 16708
rect 18196 16668 18202 16680
rect 18690 16668 18696 16680
rect 18748 16668 18754 16720
rect 19058 16668 19064 16720
rect 19116 16708 19122 16720
rect 22112 16717 22140 16748
rect 23014 16736 23020 16788
rect 23072 16776 23078 16788
rect 23198 16776 23204 16788
rect 23072 16748 23204 16776
rect 23072 16736 23078 16748
rect 23198 16736 23204 16748
rect 23256 16776 23262 16788
rect 23934 16776 23940 16788
rect 23256 16748 23940 16776
rect 23256 16736 23262 16748
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 25498 16736 25504 16788
rect 25556 16776 25562 16788
rect 25593 16779 25651 16785
rect 25593 16776 25605 16779
rect 25556 16748 25605 16776
rect 25556 16736 25562 16748
rect 25593 16745 25605 16748
rect 25639 16745 25651 16779
rect 30282 16776 30288 16788
rect 25593 16739 25651 16745
rect 27724 16748 30288 16776
rect 19153 16711 19211 16717
rect 19153 16708 19165 16711
rect 19116 16680 19165 16708
rect 19116 16668 19122 16680
rect 19153 16677 19165 16680
rect 19199 16677 19211 16711
rect 19153 16671 19211 16677
rect 22097 16711 22155 16717
rect 22097 16677 22109 16711
rect 22143 16708 22155 16711
rect 24854 16708 24860 16720
rect 22143 16680 24860 16708
rect 22143 16677 22155 16680
rect 22097 16671 22155 16677
rect 16316 16612 16436 16640
rect 17129 16643 17187 16649
rect 16316 16572 16344 16612
rect 17129 16609 17141 16643
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16609 17279 16643
rect 17221 16603 17279 16609
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 17494 16640 17500 16652
rect 17451 16612 17500 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 15856 16544 16344 16572
rect 16758 16532 16764 16584
rect 16816 16532 16822 16584
rect 17034 16532 17040 16584
rect 17092 16572 17098 16584
rect 17236 16572 17264 16603
rect 17092 16544 17264 16572
rect 17092 16532 17098 16544
rect 10560 16476 12434 16504
rect 10560 16464 10566 16476
rect 12894 16464 12900 16516
rect 12952 16504 12958 16516
rect 17420 16504 17448 16603
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 18782 16600 18788 16652
rect 18840 16600 18846 16652
rect 19242 16600 19248 16652
rect 19300 16600 19306 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16609 19487 16643
rect 19429 16603 19487 16609
rect 18673 16575 18731 16581
rect 18673 16541 18685 16575
rect 18719 16572 18731 16575
rect 18966 16572 18972 16584
rect 18719 16544 18972 16572
rect 18719 16541 18731 16544
rect 18673 16535 18731 16541
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 19061 16575 19119 16581
rect 19061 16541 19073 16575
rect 19107 16541 19119 16575
rect 19444 16572 19472 16603
rect 21266 16600 21272 16652
rect 21324 16600 21330 16652
rect 22756 16649 22784 16680
rect 24854 16668 24860 16680
rect 24912 16668 24918 16720
rect 25038 16668 25044 16720
rect 25096 16708 25102 16720
rect 26421 16711 26479 16717
rect 26421 16708 26433 16711
rect 25096 16680 26433 16708
rect 25096 16668 25102 16680
rect 26421 16677 26433 16680
rect 26467 16677 26479 16711
rect 27724 16708 27752 16748
rect 30282 16736 30288 16748
rect 30340 16736 30346 16788
rect 30377 16779 30435 16785
rect 30377 16745 30389 16779
rect 30423 16745 30435 16779
rect 30377 16739 30435 16745
rect 29086 16708 29092 16720
rect 26421 16671 26479 16677
rect 26804 16680 27016 16708
rect 26804 16652 26832 16680
rect 22741 16643 22799 16649
rect 22741 16609 22753 16643
rect 22787 16609 22799 16643
rect 22741 16603 22799 16609
rect 23198 16600 23204 16652
rect 23256 16640 23262 16652
rect 23293 16643 23351 16649
rect 23293 16640 23305 16643
rect 23256 16612 23305 16640
rect 23256 16600 23262 16612
rect 23293 16609 23305 16612
rect 23339 16609 23351 16643
rect 23293 16603 23351 16609
rect 23382 16600 23388 16652
rect 23440 16600 23446 16652
rect 23477 16643 23535 16649
rect 23477 16609 23489 16643
rect 23523 16609 23535 16643
rect 23477 16603 23535 16609
rect 19518 16572 19524 16584
rect 19444 16544 19524 16572
rect 19061 16535 19119 16541
rect 12952 16476 17448 16504
rect 19076 16504 19104 16535
rect 19518 16532 19524 16544
rect 19576 16572 19582 16584
rect 19794 16572 19800 16584
rect 19576 16544 19800 16572
rect 19576 16532 19582 16544
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 20346 16581 20352 16584
rect 20165 16575 20223 16581
rect 20165 16572 20177 16575
rect 19996 16544 20177 16572
rect 19886 16504 19892 16516
rect 19076 16476 19892 16504
rect 12952 16464 12958 16476
rect 19886 16464 19892 16476
rect 19944 16464 19950 16516
rect 5810 16436 5816 16448
rect 3712 16408 5816 16436
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 9766 16396 9772 16448
rect 9824 16396 9830 16448
rect 9950 16396 9956 16448
rect 10008 16396 10014 16448
rect 12802 16396 12808 16448
rect 12860 16436 12866 16448
rect 16298 16436 16304 16448
rect 12860 16408 16304 16436
rect 12860 16396 12866 16408
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 17037 16439 17095 16445
rect 17037 16436 17049 16439
rect 16908 16408 17049 16436
rect 16908 16396 16914 16408
rect 17037 16405 17049 16408
rect 17083 16405 17095 16439
rect 17037 16399 17095 16405
rect 17126 16396 17132 16448
rect 17184 16436 17190 16448
rect 19996 16436 20024 16544
rect 20165 16541 20177 16544
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 20303 16575 20352 16581
rect 20303 16541 20315 16575
rect 20349 16541 20352 16575
rect 20303 16535 20352 16541
rect 20346 16532 20352 16535
rect 20404 16532 20410 16584
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16572 20499 16575
rect 20622 16572 20628 16584
rect 20487 16544 20628 16572
rect 20487 16541 20499 16544
rect 20441 16535 20499 16541
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 23014 16532 23020 16584
rect 23072 16572 23078 16584
rect 23400 16572 23428 16600
rect 23072 16544 23428 16572
rect 23072 16532 23078 16544
rect 23492 16504 23520 16603
rect 23566 16600 23572 16652
rect 23624 16630 23630 16652
rect 23673 16643 23731 16649
rect 23673 16630 23685 16643
rect 23624 16609 23685 16630
rect 23719 16609 23731 16643
rect 23624 16603 23731 16609
rect 23624 16602 23704 16603
rect 23624 16600 23630 16602
rect 24210 16600 24216 16652
rect 24268 16600 24274 16652
rect 24486 16649 24492 16652
rect 24480 16603 24492 16649
rect 24486 16600 24492 16603
rect 24544 16600 24550 16652
rect 25682 16600 25688 16652
rect 25740 16600 25746 16652
rect 25777 16643 25835 16649
rect 25777 16609 25789 16643
rect 25823 16640 25835 16643
rect 25866 16640 25872 16652
rect 25823 16612 25872 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 25866 16600 25872 16612
rect 25924 16600 25930 16652
rect 25958 16600 25964 16652
rect 26016 16600 26022 16652
rect 26050 16600 26056 16652
rect 26108 16600 26114 16652
rect 26142 16600 26148 16652
rect 26200 16640 26206 16652
rect 26697 16643 26755 16649
rect 26697 16640 26709 16643
rect 26200 16612 26709 16640
rect 26200 16600 26206 16612
rect 26697 16609 26709 16612
rect 26743 16609 26755 16643
rect 26697 16603 26755 16609
rect 26786 16600 26792 16652
rect 26844 16600 26850 16652
rect 26881 16643 26939 16649
rect 26881 16609 26893 16643
rect 26927 16609 26939 16643
rect 26881 16603 26939 16609
rect 25222 16532 25228 16584
rect 25280 16572 25286 16584
rect 26160 16572 26188 16600
rect 25280 16544 26188 16572
rect 26237 16575 26295 16581
rect 25280 16532 25286 16544
rect 26237 16541 26249 16575
rect 26283 16572 26295 16575
rect 26896 16572 26924 16603
rect 26283 16544 26924 16572
rect 26988 16572 27016 16680
rect 27632 16680 27752 16708
rect 28184 16680 29092 16708
rect 27065 16643 27123 16649
rect 27065 16609 27077 16643
rect 27111 16640 27123 16643
rect 27430 16640 27436 16652
rect 27111 16612 27436 16640
rect 27111 16609 27123 16612
rect 27065 16603 27123 16609
rect 27430 16600 27436 16612
rect 27488 16600 27494 16652
rect 27632 16649 27660 16680
rect 27617 16643 27675 16649
rect 27617 16609 27629 16643
rect 27663 16609 27675 16643
rect 27617 16603 27675 16609
rect 27709 16643 27767 16649
rect 27709 16609 27721 16643
rect 27755 16609 27767 16643
rect 27709 16603 27767 16609
rect 27801 16643 27859 16649
rect 27801 16609 27813 16643
rect 27847 16640 27859 16643
rect 27982 16640 27988 16652
rect 27847 16612 27988 16640
rect 27847 16609 27859 16612
rect 27801 16603 27859 16609
rect 27724 16572 27752 16603
rect 27982 16600 27988 16612
rect 28040 16600 28046 16652
rect 28184 16649 28212 16680
rect 29086 16668 29092 16680
rect 29144 16668 29150 16720
rect 29454 16668 29460 16720
rect 29512 16708 29518 16720
rect 29914 16708 29920 16720
rect 29512 16680 29920 16708
rect 29512 16668 29518 16680
rect 29914 16668 29920 16680
rect 29972 16668 29978 16720
rect 30392 16708 30420 16739
rect 30392 16680 30880 16708
rect 28169 16643 28227 16649
rect 28169 16609 28181 16643
rect 28215 16609 28227 16643
rect 28425 16643 28483 16649
rect 28425 16640 28437 16643
rect 28169 16603 28227 16609
rect 28276 16612 28437 16640
rect 26988 16544 27752 16572
rect 28077 16575 28135 16581
rect 26283 16541 26295 16544
rect 26237 16535 26295 16541
rect 28077 16541 28089 16575
rect 28123 16572 28135 16575
rect 28276 16572 28304 16612
rect 28425 16609 28437 16612
rect 28471 16609 28483 16643
rect 28425 16603 28483 16609
rect 29362 16600 29368 16652
rect 29420 16640 29426 16652
rect 30009 16643 30067 16649
rect 30009 16640 30021 16643
rect 29420 16612 30021 16640
rect 29420 16600 29426 16612
rect 30009 16609 30021 16612
rect 30055 16609 30067 16643
rect 30469 16643 30527 16649
rect 30469 16640 30481 16643
rect 30009 16603 30067 16609
rect 30116 16612 30481 16640
rect 28123 16544 28304 16572
rect 28123 16541 28135 16544
rect 28077 16535 28135 16541
rect 29638 16532 29644 16584
rect 29696 16572 29702 16584
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29696 16544 29745 16572
rect 29696 16532 29702 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 23658 16504 23664 16516
rect 23492 16476 23664 16504
rect 23658 16464 23664 16476
rect 23716 16464 23722 16516
rect 30116 16504 30144 16612
rect 30469 16609 30481 16612
rect 30515 16609 30527 16643
rect 30469 16603 30527 16609
rect 30558 16600 30564 16652
rect 30616 16600 30622 16652
rect 30742 16600 30748 16652
rect 30800 16600 30806 16652
rect 30852 16649 30880 16680
rect 30837 16643 30895 16649
rect 30837 16609 30849 16643
rect 30883 16609 30895 16643
rect 30837 16603 30895 16609
rect 30282 16532 30288 16584
rect 30340 16572 30346 16584
rect 31021 16575 31079 16581
rect 31021 16572 31033 16575
rect 30340 16544 31033 16572
rect 30340 16532 30346 16544
rect 31021 16541 31033 16544
rect 31067 16541 31079 16575
rect 31021 16535 31079 16541
rect 29196 16476 30144 16504
rect 17184 16408 20024 16436
rect 17184 16396 17190 16408
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21085 16439 21143 16445
rect 21085 16436 21097 16439
rect 21048 16408 21097 16436
rect 21048 16396 21054 16408
rect 21085 16405 21097 16408
rect 21131 16405 21143 16439
rect 21085 16399 21143 16405
rect 23017 16439 23075 16445
rect 23017 16405 23029 16439
rect 23063 16436 23075 16439
rect 23198 16436 23204 16448
rect 23063 16408 23204 16436
rect 23063 16405 23075 16408
rect 23017 16399 23075 16405
rect 23198 16396 23204 16408
rect 23256 16396 23262 16448
rect 24946 16396 24952 16448
rect 25004 16436 25010 16448
rect 25682 16436 25688 16448
rect 25004 16408 25688 16436
rect 25004 16396 25010 16408
rect 25682 16396 25688 16408
rect 25740 16436 25746 16448
rect 27522 16436 27528 16448
rect 25740 16408 27528 16436
rect 25740 16396 25746 16408
rect 27522 16396 27528 16408
rect 27580 16436 27586 16448
rect 27982 16436 27988 16448
rect 27580 16408 27988 16436
rect 27580 16396 27586 16408
rect 27982 16396 27988 16408
rect 28040 16436 28046 16448
rect 29196 16436 29224 16476
rect 28040 16408 29224 16436
rect 28040 16396 28046 16408
rect 29546 16396 29552 16448
rect 29604 16396 29610 16448
rect 552 16346 31648 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 11436 16346
rect 11488 16294 11500 16346
rect 11552 16294 11564 16346
rect 11616 16294 11628 16346
rect 11680 16294 11692 16346
rect 11744 16294 19210 16346
rect 19262 16294 19274 16346
rect 19326 16294 19338 16346
rect 19390 16294 19402 16346
rect 19454 16294 19466 16346
rect 19518 16294 26984 16346
rect 27036 16294 27048 16346
rect 27100 16294 27112 16346
rect 27164 16294 27176 16346
rect 27228 16294 27240 16346
rect 27292 16294 31648 16346
rect 552 16272 31648 16294
rect 2958 16192 2964 16244
rect 3016 16232 3022 16244
rect 3053 16235 3111 16241
rect 3053 16232 3065 16235
rect 3016 16204 3065 16232
rect 3016 16192 3022 16204
rect 3053 16201 3065 16204
rect 3099 16232 3111 16235
rect 4062 16232 4068 16244
rect 3099 16204 4068 16232
rect 3099 16201 3111 16204
rect 3053 16195 3111 16201
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8168 16204 9444 16232
rect 8168 16192 8174 16204
rect 2682 16124 2688 16176
rect 2740 16164 2746 16176
rect 2740 16124 2774 16164
rect 2866 16124 2872 16176
rect 2924 16164 2930 16176
rect 3326 16164 3332 16176
rect 2924 16136 3332 16164
rect 2924 16124 2930 16136
rect 3326 16124 3332 16136
rect 3384 16124 3390 16176
rect 6733 16167 6791 16173
rect 6733 16133 6745 16167
rect 6779 16164 6791 16167
rect 7006 16164 7012 16176
rect 6779 16136 7012 16164
rect 6779 16133 6791 16136
rect 6733 16127 6791 16133
rect 7006 16124 7012 16136
rect 7064 16164 7070 16176
rect 7742 16164 7748 16176
rect 7064 16136 7748 16164
rect 7064 16124 7070 16136
rect 7742 16124 7748 16136
rect 7800 16124 7806 16176
rect 8478 16124 8484 16176
rect 8536 16164 8542 16176
rect 9309 16167 9367 16173
rect 9309 16164 9321 16167
rect 8536 16136 9321 16164
rect 8536 16124 8542 16136
rect 9309 16133 9321 16136
rect 9355 16133 9367 16167
rect 9416 16164 9444 16204
rect 9490 16192 9496 16244
rect 9548 16192 9554 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9824 16204 9873 16232
rect 9824 16192 9830 16204
rect 9861 16201 9873 16204
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 9674 16164 9680 16176
rect 9416 16136 9680 16164
rect 9309 16127 9367 16133
rect 1578 16096 1584 16108
rect 1412 16068 1584 16096
rect 1412 16037 1440 16068
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 2746 16096 2774 16124
rect 9324 16096 9352 16127
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 9490 16096 9496 16108
rect 2746 16068 9168 16096
rect 9324 16068 9496 16096
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1673 16031 1731 16037
rect 1673 16028 1685 16031
rect 1535 16000 1685 16028
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 1673 15997 1685 16000
rect 1719 15997 1731 16031
rect 1673 15991 1731 15997
rect 2406 15988 2412 16040
rect 2464 16028 2470 16040
rect 2464 16000 3188 16028
rect 2464 15988 2470 16000
rect 1940 15963 1998 15969
rect 1940 15929 1952 15963
rect 1986 15960 1998 15963
rect 3160 15960 3188 16000
rect 3326 15988 3332 16040
rect 3384 15988 3390 16040
rect 4246 15988 4252 16040
rect 4304 15988 4310 16040
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 15997 4399 16031
rect 4341 15991 4399 15997
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 5626 16028 5632 16040
rect 4663 16000 5632 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4154 15960 4160 15972
rect 1986 15932 2774 15960
rect 3160 15932 4160 15960
rect 1986 15929 1998 15932
rect 1940 15923 1998 15929
rect 2746 15892 2774 15932
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 2958 15892 2964 15904
rect 2746 15864 2964 15892
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 3878 15852 3884 15904
rect 3936 15852 3942 15904
rect 3970 15852 3976 15904
rect 4028 15852 4034 15904
rect 4062 15852 4068 15904
rect 4120 15892 4126 15904
rect 4356 15892 4384 15991
rect 4448 15960 4476 15991
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 16028 7527 16031
rect 7653 16031 7711 16037
rect 7653 16028 7665 16031
rect 7515 16000 7665 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 7653 15997 7665 16000
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 7742 15988 7748 16040
rect 7800 15988 7806 16040
rect 7834 15988 7840 16040
rect 7892 15988 7898 16040
rect 7929 16031 7987 16037
rect 7929 15997 7941 16031
rect 7975 16028 7987 16031
rect 8018 16028 8024 16040
rect 7975 16000 8024 16028
rect 7975 15997 7987 16000
rect 7929 15991 7987 15997
rect 4706 15960 4712 15972
rect 4448 15932 4712 15960
rect 4706 15920 4712 15932
rect 4764 15920 4770 15972
rect 6733 15963 6791 15969
rect 6733 15929 6745 15963
rect 6779 15960 6791 15963
rect 6914 15960 6920 15972
rect 6779 15932 6920 15960
rect 6779 15929 6791 15932
rect 6733 15923 6791 15929
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7558 15920 7564 15972
rect 7616 15960 7622 15972
rect 7944 15960 7972 15991
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 7616 15932 7972 15960
rect 7616 15920 7622 15932
rect 9030 15920 9036 15972
rect 9088 15920 9094 15972
rect 9140 15960 9168 16068
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 9692 16028 9720 16124
rect 9876 16096 9904 16195
rect 10042 16192 10048 16244
rect 10100 16192 10106 16244
rect 10410 16192 10416 16244
rect 10468 16192 10474 16244
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 11241 16235 11299 16241
rect 11241 16232 11253 16235
rect 10652 16204 11253 16232
rect 10652 16192 10658 16204
rect 11241 16201 11253 16204
rect 11287 16201 11299 16235
rect 11241 16195 11299 16201
rect 15562 16192 15568 16244
rect 15620 16232 15626 16244
rect 15620 16204 16160 16232
rect 15620 16192 15626 16204
rect 10321 16167 10379 16173
rect 10321 16133 10333 16167
rect 10367 16164 10379 16167
rect 10962 16164 10968 16176
rect 10367 16136 10968 16164
rect 10367 16133 10379 16136
rect 10321 16127 10379 16133
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 11057 16167 11115 16173
rect 11057 16133 11069 16167
rect 11103 16133 11115 16167
rect 11057 16127 11115 16133
rect 9876 16068 10916 16096
rect 9953 16031 10011 16037
rect 9953 16028 9965 16031
rect 9692 16000 9965 16028
rect 9953 15997 9965 16000
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 10597 16031 10655 16037
rect 10597 16028 10609 16031
rect 10376 16000 10609 16028
rect 10376 15988 10382 16000
rect 10597 15997 10609 16000
rect 10643 15997 10655 16031
rect 10597 15991 10655 15997
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 10778 16028 10784 16040
rect 10735 16000 10784 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 10888 16037 10916 16068
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11072 16028 11100 16127
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15749 16167 15807 16173
rect 15749 16164 15761 16167
rect 15344 16136 15761 16164
rect 15344 16124 15350 16136
rect 15749 16133 15761 16136
rect 15795 16133 15807 16167
rect 16132 16164 16160 16204
rect 16206 16192 16212 16244
rect 16264 16192 16270 16244
rect 19702 16192 19708 16244
rect 19760 16232 19766 16244
rect 22649 16235 22707 16241
rect 19760 16204 20484 16232
rect 19760 16192 19766 16204
rect 16132 16136 16712 16164
rect 15749 16127 15807 16133
rect 16684 16108 16712 16136
rect 16114 16096 16120 16108
rect 15764 16068 16120 16096
rect 11011 16000 11100 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 11146 15988 11152 16040
rect 11204 16028 11210 16040
rect 12345 16031 12403 16037
rect 12345 16028 12357 16031
rect 11204 16000 12357 16028
rect 11204 15988 11210 16000
rect 12345 15997 12357 16000
rect 12391 15997 12403 16031
rect 12345 15991 12403 15997
rect 12526 15988 12532 16040
rect 12584 15988 12590 16040
rect 12618 15988 12624 16040
rect 12676 15988 12682 16040
rect 12713 16031 12771 16037
rect 12713 15997 12725 16031
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 10502 15960 10508 15972
rect 9140 15932 10508 15960
rect 10502 15920 10508 15932
rect 10560 15920 10566 15972
rect 11425 15963 11483 15969
rect 11425 15960 11437 15963
rect 10980 15932 11437 15960
rect 4120 15864 4384 15892
rect 4120 15852 4126 15864
rect 7190 15852 7196 15904
rect 7248 15852 7254 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 9048 15892 9076 15920
rect 10980 15904 11008 15932
rect 11425 15929 11437 15932
rect 11471 15929 11483 15963
rect 11425 15923 11483 15929
rect 11974 15920 11980 15972
rect 12032 15960 12038 15972
rect 12728 15960 12756 15991
rect 13170 15988 13176 16040
rect 13228 15988 13234 16040
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 13311 16000 13553 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 13541 15997 13553 16000
rect 13587 15997 13599 16031
rect 13541 15991 13599 15997
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 15562 16028 15568 16040
rect 14148 16000 15568 16028
rect 14148 15988 14154 16000
rect 15562 15988 15568 16000
rect 15620 15988 15626 16040
rect 15764 16037 15792 16068
rect 16114 16056 16120 16068
rect 16172 16096 16178 16108
rect 16577 16099 16635 16105
rect 16577 16096 16589 16099
rect 16172 16068 16589 16096
rect 16172 16056 16178 16068
rect 16577 16065 16589 16068
rect 16623 16065 16635 16099
rect 16577 16059 16635 16065
rect 16666 16056 16672 16108
rect 16724 16056 16730 16108
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 16390 16028 16396 16040
rect 15749 15991 15807 15997
rect 16132 16000 16396 16028
rect 16132 15969 16160 16000
rect 16390 15988 16396 16000
rect 16448 16037 16454 16040
rect 16448 16031 16511 16037
rect 16448 15997 16465 16031
rect 16499 16028 16511 16031
rect 16499 16000 18368 16028
rect 16499 15997 16511 16000
rect 16448 15991 16511 15997
rect 16448 15988 16454 15991
rect 12032 15932 12756 15960
rect 12989 15963 13047 15969
rect 12032 15920 12038 15932
rect 12989 15929 13001 15963
rect 13035 15960 13047 15963
rect 13786 15963 13844 15969
rect 13786 15960 13798 15963
rect 13035 15932 13798 15960
rect 13035 15929 13047 15932
rect 12989 15923 13047 15929
rect 13786 15929 13798 15932
rect 13832 15929 13844 15963
rect 13786 15923 13844 15929
rect 16117 15963 16175 15969
rect 16117 15929 16129 15963
rect 16163 15929 16175 15963
rect 16117 15923 16175 15929
rect 17037 15963 17095 15969
rect 17037 15929 17049 15963
rect 17083 15960 17095 15963
rect 17497 15963 17555 15969
rect 17497 15960 17509 15963
rect 17083 15932 17509 15960
rect 17083 15929 17095 15932
rect 17037 15923 17095 15929
rect 17497 15929 17509 15932
rect 17543 15929 17555 15963
rect 17497 15923 17555 15929
rect 17865 15963 17923 15969
rect 17865 15929 17877 15963
rect 17911 15960 17923 15963
rect 18230 15960 18236 15972
rect 17911 15932 18236 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 7331 15864 9076 15892
rect 9677 15895 9735 15901
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 9677 15861 9689 15895
rect 9723 15892 9735 15895
rect 10962 15892 10968 15904
rect 9723 15864 10968 15892
rect 9723 15861 9735 15864
rect 9677 15855 9735 15861
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11225 15895 11283 15901
rect 11225 15892 11237 15895
rect 11112 15864 11237 15892
rect 11112 15852 11118 15864
rect 11225 15861 11237 15864
rect 11271 15861 11283 15895
rect 11225 15855 11283 15861
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 14921 15895 14979 15901
rect 14921 15892 14933 15895
rect 11572 15864 14933 15892
rect 11572 15852 11578 15864
rect 14921 15861 14933 15864
rect 14967 15861 14979 15895
rect 14921 15855 14979 15861
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 17052 15892 17080 15923
rect 18230 15920 18236 15932
rect 18288 15920 18294 15972
rect 18340 15960 18368 16000
rect 18690 15988 18696 16040
rect 18748 15988 18754 16040
rect 18785 16031 18843 16037
rect 18785 15997 18797 16031
rect 18831 16028 18843 16031
rect 18969 16031 19027 16037
rect 18969 16028 18981 16031
rect 18831 16000 18981 16028
rect 18831 15997 18843 16000
rect 18785 15991 18843 15997
rect 18969 15997 18981 16000
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 19236 16031 19294 16037
rect 19236 15997 19248 16031
rect 19282 16028 19294 16031
rect 19610 16028 19616 16040
rect 19282 16000 19616 16028
rect 19282 15997 19294 16000
rect 19236 15991 19294 15997
rect 19610 15988 19616 16000
rect 19668 15988 19674 16040
rect 20456 16028 20484 16204
rect 21652 16204 22600 16232
rect 21358 16056 21364 16108
rect 21416 16056 21422 16108
rect 21545 16099 21603 16105
rect 21545 16065 21557 16099
rect 21591 16096 21603 16099
rect 21652 16096 21680 16204
rect 22005 16167 22063 16173
rect 22005 16133 22017 16167
rect 22051 16133 22063 16167
rect 22572 16164 22600 16204
rect 22649 16201 22661 16235
rect 22695 16232 22707 16235
rect 22922 16232 22928 16244
rect 22695 16204 22928 16232
rect 22695 16201 22707 16204
rect 22649 16195 22707 16201
rect 22922 16192 22928 16204
rect 22980 16192 22986 16244
rect 23216 16204 24164 16232
rect 23106 16164 23112 16176
rect 22572 16136 23112 16164
rect 22005 16127 22063 16133
rect 21591 16068 21680 16096
rect 22020 16096 22048 16127
rect 23106 16124 23112 16136
rect 23164 16164 23170 16176
rect 23216 16164 23244 16204
rect 23164 16136 23244 16164
rect 23164 16124 23170 16136
rect 23658 16096 23664 16108
rect 22020 16068 22508 16096
rect 21591 16065 21603 16068
rect 21545 16059 21603 16065
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20456 16000 20545 16028
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20254 15960 20260 15972
rect 18340 15932 20260 15960
rect 20254 15920 20260 15932
rect 20312 15920 20318 15972
rect 20548 15960 20576 15991
rect 20622 15988 20628 16040
rect 20680 16028 20686 16040
rect 20717 16031 20775 16037
rect 20717 16028 20729 16031
rect 20680 16000 20729 16028
rect 20680 15988 20686 16000
rect 20717 15997 20729 16000
rect 20763 15997 20775 16031
rect 20717 15991 20775 15997
rect 20806 15988 20812 16040
rect 20864 15988 20870 16040
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 16028 20959 16031
rect 21560 16028 21588 16059
rect 20947 16000 21588 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 22094 15988 22100 16040
rect 22152 15988 22158 16040
rect 22189 16031 22247 16037
rect 22189 15997 22201 16031
rect 22235 16025 22247 16031
rect 22278 16025 22284 16040
rect 22235 15997 22284 16025
rect 22189 15991 22247 15997
rect 22278 15988 22284 15997
rect 22336 15988 22342 16040
rect 22370 15988 22376 16040
rect 22428 15988 22434 16040
rect 22480 16037 22508 16068
rect 23400 16068 23664 16096
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22646 15988 22652 16040
rect 22704 16028 22710 16040
rect 22741 16031 22799 16037
rect 22741 16028 22753 16031
rect 22704 16000 22753 16028
rect 22704 15988 22710 16000
rect 22741 15997 22753 16000
rect 22787 15997 22799 16031
rect 22741 15991 22799 15997
rect 23109 16031 23167 16037
rect 23109 15997 23121 16031
rect 23155 15997 23167 16031
rect 23109 15991 23167 15997
rect 21082 15960 21088 15972
rect 20548 15932 21088 15960
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 21177 15963 21235 15969
rect 21177 15929 21189 15963
rect 21223 15960 21235 15963
rect 21910 15960 21916 15972
rect 21223 15932 21916 15960
rect 21223 15929 21235 15932
rect 21177 15923 21235 15929
rect 21910 15920 21916 15932
rect 21968 15920 21974 15972
rect 23124 15904 23152 15991
rect 23198 15988 23204 16040
rect 23256 15988 23262 16040
rect 23400 16037 23428 16068
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 24136 16096 24164 16204
rect 24486 16192 24492 16244
rect 24544 16192 24550 16244
rect 26142 16192 26148 16244
rect 26200 16192 26206 16244
rect 28626 16192 28632 16244
rect 28684 16232 28690 16244
rect 28813 16235 28871 16241
rect 28813 16232 28825 16235
rect 28684 16204 28825 16232
rect 28684 16192 28690 16204
rect 28813 16201 28825 16204
rect 28859 16201 28871 16235
rect 28813 16195 28871 16201
rect 29641 16235 29699 16241
rect 29641 16201 29653 16235
rect 29687 16232 29699 16235
rect 30558 16232 30564 16244
rect 29687 16204 30564 16232
rect 29687 16201 29699 16204
rect 29641 16195 29699 16201
rect 30558 16192 30564 16204
rect 30616 16192 30622 16244
rect 26786 16124 26792 16176
rect 26844 16164 26850 16176
rect 26844 16136 28488 16164
rect 26844 16124 26850 16136
rect 24136 16068 24256 16096
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 23474 15988 23480 16040
rect 23532 15988 23538 16040
rect 23842 15988 23848 16040
rect 23900 15988 23906 16040
rect 24029 16031 24087 16037
rect 24029 15997 24041 16031
rect 24075 15997 24087 16031
rect 24029 15991 24087 15997
rect 23661 15963 23719 15969
rect 23661 15929 23673 15963
rect 23707 15960 23719 15963
rect 24044 15960 24072 15991
rect 24118 15988 24124 16040
rect 24176 15988 24182 16040
rect 24228 16037 24256 16068
rect 26050 16056 26056 16108
rect 26108 16096 26114 16108
rect 26602 16096 26608 16108
rect 26108 16068 26608 16096
rect 26108 16056 26114 16068
rect 26602 16056 26608 16068
rect 26660 16096 26666 16108
rect 26660 16068 28396 16096
rect 26660 16056 26666 16068
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 15997 24271 16031
rect 24213 15991 24271 15997
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 25038 16037 25044 16040
rect 25032 16028 25044 16037
rect 24999 16000 25044 16028
rect 25032 15991 25044 16000
rect 25038 15988 25044 15991
rect 25096 15988 25102 16040
rect 27617 16031 27675 16037
rect 27617 15997 27629 16031
rect 27663 15997 27675 16031
rect 27617 15991 27675 15997
rect 24946 15960 24952 15972
rect 23707 15932 24072 15960
rect 24105 15932 24952 15960
rect 23707 15929 23719 15932
rect 23661 15923 23719 15929
rect 15712 15864 17080 15892
rect 15712 15852 15718 15864
rect 17126 15852 17132 15904
rect 17184 15852 17190 15904
rect 19518 15852 19524 15904
rect 19576 15892 19582 15904
rect 19886 15892 19892 15904
rect 19576 15864 19892 15892
rect 19576 15852 19582 15864
rect 19886 15852 19892 15864
rect 19944 15892 19950 15904
rect 20349 15895 20407 15901
rect 20349 15892 20361 15895
rect 19944 15864 20361 15892
rect 19944 15852 19950 15864
rect 20349 15861 20361 15864
rect 20395 15892 20407 15895
rect 21450 15892 21456 15904
rect 20395 15864 21456 15892
rect 20395 15861 20407 15864
rect 20349 15855 20407 15861
rect 21450 15852 21456 15864
rect 21508 15892 21514 15904
rect 21637 15895 21695 15901
rect 21637 15892 21649 15895
rect 21508 15864 21649 15892
rect 21508 15852 21514 15864
rect 21637 15861 21649 15864
rect 21683 15892 21695 15895
rect 22094 15892 22100 15904
rect 21683 15864 22100 15892
rect 21683 15861 21695 15864
rect 21637 15855 21695 15861
rect 22094 15852 22100 15864
rect 22152 15852 22158 15904
rect 22922 15852 22928 15904
rect 22980 15852 22986 15904
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 24105 15892 24133 15932
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 26602 15920 26608 15972
rect 26660 15920 26666 15972
rect 27338 15920 27344 15972
rect 27396 15960 27402 15972
rect 27632 15960 27660 15991
rect 28166 15988 28172 16040
rect 28224 15988 28230 16040
rect 28368 16037 28396 16068
rect 28460 16037 28488 16136
rect 29546 16096 29552 16108
rect 28552 16068 29552 16096
rect 28552 16037 28580 16068
rect 29546 16056 29552 16068
rect 29604 16056 29610 16108
rect 28353 16031 28411 16037
rect 28353 15997 28365 16031
rect 28399 15997 28411 16031
rect 28353 15991 28411 15997
rect 28445 16031 28503 16037
rect 28445 15997 28457 16031
rect 28491 15997 28503 16031
rect 28445 15991 28503 15997
rect 28537 16031 28595 16037
rect 28537 15997 28549 16031
rect 28583 15997 28595 16031
rect 28537 15991 28595 15997
rect 28997 16031 29055 16037
rect 28997 15997 29009 16031
rect 29043 15997 29055 16031
rect 28997 15991 29055 15997
rect 27396 15932 27660 15960
rect 29012 15960 29040 15991
rect 29086 15988 29092 16040
rect 29144 16028 29150 16040
rect 29181 16031 29239 16037
rect 29181 16028 29193 16031
rect 29144 16000 29193 16028
rect 29144 15988 29150 16000
rect 29181 15997 29193 16000
rect 29227 15997 29239 16031
rect 29181 15991 29239 15997
rect 29270 15988 29276 16040
rect 29328 15988 29334 16040
rect 29362 15988 29368 16040
rect 29420 15988 29426 16040
rect 29914 15988 29920 16040
rect 29972 15988 29978 16040
rect 29733 15963 29791 15969
rect 29733 15960 29745 15963
rect 29012 15932 29745 15960
rect 27396 15920 27402 15932
rect 29733 15929 29745 15932
rect 29779 15929 29791 15963
rect 29733 15923 29791 15929
rect 30101 15963 30159 15969
rect 30101 15929 30113 15963
rect 30147 15929 30159 15963
rect 30101 15923 30159 15929
rect 23164 15864 24133 15892
rect 23164 15852 23170 15864
rect 24578 15852 24584 15904
rect 24636 15892 24642 15904
rect 29914 15892 29920 15904
rect 24636 15864 29920 15892
rect 24636 15852 24642 15864
rect 29914 15852 29920 15864
rect 29972 15892 29978 15904
rect 30116 15892 30144 15923
rect 29972 15864 30144 15892
rect 29972 15852 29978 15864
rect 552 15802 31648 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 12096 15802
rect 12148 15750 12160 15802
rect 12212 15750 12224 15802
rect 12276 15750 12288 15802
rect 12340 15750 12352 15802
rect 12404 15750 19870 15802
rect 19922 15750 19934 15802
rect 19986 15750 19998 15802
rect 20050 15750 20062 15802
rect 20114 15750 20126 15802
rect 20178 15750 27644 15802
rect 27696 15750 27708 15802
rect 27760 15750 27772 15802
rect 27824 15750 27836 15802
rect 27888 15750 27900 15802
rect 27952 15750 31648 15802
rect 552 15728 31648 15750
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3016 15660 3433 15688
rect 3016 15648 3022 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 3878 15648 3884 15700
rect 3936 15688 3942 15700
rect 4525 15691 4583 15697
rect 3936 15660 4384 15688
rect 3936 15648 3942 15660
rect 2216 15623 2274 15629
rect 2216 15589 2228 15623
rect 2262 15620 2274 15623
rect 3970 15620 3976 15632
rect 2262 15592 3976 15620
rect 2262 15589 2274 15592
rect 2216 15583 2274 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 4154 15580 4160 15632
rect 4212 15580 4218 15632
rect 4356 15629 4384 15660
rect 4525 15657 4537 15691
rect 4571 15688 4583 15691
rect 4706 15688 4712 15700
rect 4571 15660 4712 15688
rect 4571 15657 4583 15660
rect 4525 15651 4583 15657
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7834 15688 7840 15700
rect 6972 15660 7840 15688
rect 6972 15648 6978 15660
rect 7834 15648 7840 15660
rect 7892 15688 7898 15700
rect 13630 15688 13636 15700
rect 7892 15660 8248 15688
rect 7892 15648 7898 15660
rect 4341 15623 4399 15629
rect 4341 15589 4353 15623
rect 4387 15589 4399 15623
rect 4341 15583 4399 15589
rect 7101 15623 7159 15629
rect 7101 15589 7113 15623
rect 7147 15620 7159 15623
rect 7190 15620 7196 15632
rect 7147 15592 7196 15620
rect 7147 15589 7159 15592
rect 7101 15583 7159 15589
rect 7190 15580 7196 15592
rect 7248 15620 7254 15632
rect 8220 15620 8248 15660
rect 9692 15660 13636 15688
rect 9582 15620 9588 15632
rect 7248 15592 7880 15620
rect 8220 15592 9588 15620
rect 7248 15580 7254 15592
rect 1670 15512 1676 15564
rect 1728 15552 1734 15564
rect 1949 15555 2007 15561
rect 1949 15552 1961 15555
rect 1728 15524 1961 15552
rect 1728 15512 1734 15524
rect 1949 15521 1961 15524
rect 1995 15521 2007 15555
rect 1949 15515 2007 15521
rect 3694 15512 3700 15564
rect 3752 15512 3758 15564
rect 3786 15512 3792 15564
rect 3844 15512 3850 15564
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15521 3939 15555
rect 3881 15515 3939 15521
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 5626 15552 5632 15564
rect 4111 15524 5632 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 3142 15444 3148 15496
rect 3200 15484 3206 15496
rect 3896 15484 3924 15515
rect 3200 15456 3924 15484
rect 3200 15444 3206 15456
rect 2958 15376 2964 15428
rect 3016 15416 3022 15428
rect 3329 15419 3387 15425
rect 3329 15416 3341 15419
rect 3016 15388 3341 15416
rect 3016 15376 3022 15388
rect 3329 15385 3341 15388
rect 3375 15385 3387 15419
rect 3329 15379 3387 15385
rect 3418 15376 3424 15428
rect 3476 15416 3482 15428
rect 4080 15416 4108 15515
rect 5626 15512 5632 15524
rect 5684 15512 5690 15564
rect 7852 15561 7880 15592
rect 9582 15580 9588 15592
rect 9640 15580 9646 15632
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 7837 15555 7895 15561
rect 7837 15521 7849 15555
rect 7883 15552 7895 15555
rect 8478 15552 8484 15564
rect 7883 15524 8484 15552
rect 7883 15521 7895 15524
rect 7837 15515 7895 15521
rect 5534 15444 5540 15496
rect 5592 15444 5598 15496
rect 5994 15444 6000 15496
rect 6052 15484 6058 15496
rect 6181 15487 6239 15493
rect 6181 15484 6193 15487
rect 6052 15456 6193 15484
rect 6052 15444 6058 15456
rect 6181 15453 6193 15456
rect 6227 15453 6239 15487
rect 7668 15484 7696 15515
rect 8478 15512 8484 15524
rect 8536 15512 8542 15564
rect 9030 15484 9036 15496
rect 6181 15447 6239 15453
rect 7392 15456 9036 15484
rect 3476 15388 4108 15416
rect 3476 15376 3482 15388
rect 4246 15376 4252 15428
rect 4304 15416 4310 15428
rect 4798 15416 4804 15428
rect 4304 15388 4804 15416
rect 4304 15376 4310 15388
rect 4798 15376 4804 15388
rect 4856 15416 4862 15428
rect 7392 15425 7420 15456
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9692 15484 9720 15660
rect 13630 15648 13636 15660
rect 13688 15688 13694 15700
rect 14182 15688 14188 15700
rect 13688 15660 14188 15688
rect 13688 15648 13694 15660
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 17954 15688 17960 15700
rect 16500 15660 17960 15688
rect 10318 15580 10324 15632
rect 10376 15620 10382 15632
rect 10689 15623 10747 15629
rect 10689 15620 10701 15623
rect 10376 15592 10701 15620
rect 10376 15580 10382 15592
rect 10689 15589 10701 15592
rect 10735 15589 10747 15623
rect 10689 15583 10747 15589
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10226 15552 10232 15564
rect 10008 15524 10232 15552
rect 10008 15512 10014 15524
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 10413 15555 10471 15561
rect 10413 15521 10425 15555
rect 10459 15521 10471 15555
rect 10413 15515 10471 15521
rect 9140 15456 9720 15484
rect 10045 15487 10103 15493
rect 7377 15419 7435 15425
rect 4856 15388 6960 15416
rect 4856 15376 4862 15388
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 3510 15348 3516 15360
rect 2924 15320 3516 15348
rect 2924 15308 2930 15320
rect 3510 15308 3516 15320
rect 3568 15348 3574 15360
rect 3786 15348 3792 15360
rect 3568 15320 3792 15348
rect 3568 15308 3574 15320
rect 3786 15308 3792 15320
rect 3844 15348 3850 15360
rect 4062 15348 4068 15360
rect 3844 15320 4068 15348
rect 3844 15308 3850 15320
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4982 15308 4988 15360
rect 5040 15308 5046 15360
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6788 15320 6837 15348
rect 6788 15308 6794 15320
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6932 15348 6960 15388
rect 7377 15385 7389 15419
rect 7423 15385 7435 15419
rect 9140 15416 9168 15456
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10428 15484 10456 15515
rect 10594 15512 10600 15564
rect 10652 15512 10658 15564
rect 10778 15512 10784 15564
rect 10836 15552 10842 15564
rect 11514 15552 11520 15564
rect 10836 15524 11520 15552
rect 10836 15512 10842 15524
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 14369 15555 14427 15561
rect 14369 15521 14381 15555
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 10962 15484 10968 15496
rect 10091 15456 10968 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 14384 15484 14412 15515
rect 14642 15512 14648 15564
rect 14700 15512 14706 15564
rect 16022 15512 16028 15564
rect 16080 15552 16086 15564
rect 16301 15555 16359 15561
rect 16301 15552 16313 15555
rect 16080 15524 16313 15552
rect 16080 15512 16086 15524
rect 16301 15521 16313 15524
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 15378 15484 15384 15496
rect 14384 15456 15384 15484
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 7377 15379 7435 15385
rect 7475 15388 9168 15416
rect 7475 15348 7503 15388
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 9953 15419 10011 15425
rect 9953 15416 9965 15419
rect 9732 15388 9965 15416
rect 9732 15376 9738 15388
rect 9953 15385 9965 15388
rect 9999 15416 10011 15419
rect 10134 15416 10140 15428
rect 9999 15388 10140 15416
rect 9999 15385 10011 15388
rect 9953 15379 10011 15385
rect 10134 15376 10140 15388
rect 10192 15376 10198 15428
rect 10226 15376 10232 15428
rect 10284 15376 10290 15428
rect 10502 15376 10508 15428
rect 10560 15416 10566 15428
rect 10686 15416 10692 15428
rect 10560 15388 10692 15416
rect 10560 15376 10566 15388
rect 10686 15376 10692 15388
rect 10744 15416 10750 15428
rect 12618 15416 12624 15428
rect 10744 15388 12624 15416
rect 10744 15376 10750 15388
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 13998 15376 14004 15428
rect 14056 15416 14062 15428
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 14056 15388 14565 15416
rect 14056 15376 14062 15388
rect 14553 15385 14565 15388
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 6932 15320 7503 15348
rect 6825 15311 6883 15317
rect 7558 15308 7564 15360
rect 7616 15308 7622 15360
rect 7745 15351 7803 15357
rect 7745 15317 7757 15351
rect 7791 15348 7803 15351
rect 7926 15348 7932 15360
rect 7791 15320 7932 15348
rect 7791 15317 7803 15320
rect 7745 15311 7803 15317
rect 7926 15308 7932 15320
rect 7984 15348 7990 15360
rect 11054 15348 11060 15360
rect 7984 15320 11060 15348
rect 7984 15308 7990 15320
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11974 15348 11980 15360
rect 11204 15320 11980 15348
rect 11204 15308 11210 15320
rect 11974 15308 11980 15320
rect 12032 15348 12038 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 12032 15320 12081 15348
rect 12032 15308 12038 15320
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 15562 15308 15568 15360
rect 15620 15348 15626 15360
rect 16500 15357 16528 15660
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 18230 15648 18236 15700
rect 18288 15648 18294 15700
rect 19058 15648 19064 15700
rect 19116 15648 19122 15700
rect 19153 15691 19211 15697
rect 19153 15657 19165 15691
rect 19199 15657 19211 15691
rect 19153 15651 19211 15657
rect 20533 15691 20591 15697
rect 20533 15657 20545 15691
rect 20579 15688 20591 15691
rect 20714 15688 20720 15700
rect 20579 15660 20720 15688
rect 20579 15657 20591 15660
rect 20533 15651 20591 15657
rect 17494 15620 17500 15632
rect 16592 15592 17500 15620
rect 16592 15561 16620 15592
rect 17494 15580 17500 15592
rect 17552 15580 17558 15632
rect 18966 15580 18972 15632
rect 19024 15620 19030 15632
rect 19168 15620 19196 15651
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 20901 15691 20959 15697
rect 20901 15657 20913 15691
rect 20947 15688 20959 15691
rect 21082 15688 21088 15700
rect 20947 15660 21088 15688
rect 20947 15657 20959 15660
rect 20901 15651 20959 15657
rect 21082 15648 21088 15660
rect 21140 15688 21146 15700
rect 22281 15691 22339 15697
rect 22281 15688 22293 15691
rect 21140 15660 22293 15688
rect 21140 15648 21146 15660
rect 22281 15657 22293 15660
rect 22327 15688 22339 15691
rect 22462 15688 22468 15700
rect 22327 15660 22468 15688
rect 22327 15657 22339 15660
rect 22281 15651 22339 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 22649 15691 22707 15697
rect 22649 15657 22661 15691
rect 22695 15688 22707 15691
rect 22738 15688 22744 15700
rect 22695 15660 22744 15688
rect 22695 15657 22707 15660
rect 22649 15651 22707 15657
rect 22738 15648 22744 15660
rect 22796 15688 22802 15700
rect 23106 15688 23112 15700
rect 22796 15660 23112 15688
rect 22796 15648 22802 15660
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 23658 15648 23664 15700
rect 23716 15688 23722 15700
rect 24670 15688 24676 15700
rect 23716 15660 24676 15688
rect 23716 15648 23722 15660
rect 24670 15648 24676 15660
rect 24728 15648 24734 15700
rect 24762 15648 24768 15700
rect 24820 15688 24826 15700
rect 24949 15691 25007 15697
rect 24949 15688 24961 15691
rect 24820 15660 24961 15688
rect 24820 15648 24826 15660
rect 24949 15657 24961 15660
rect 24995 15657 25007 15691
rect 28258 15688 28264 15700
rect 24949 15651 25007 15657
rect 27632 15660 28264 15688
rect 19024 15592 19196 15620
rect 20257 15623 20315 15629
rect 19024 15580 19030 15592
rect 20257 15589 20269 15623
rect 20303 15620 20315 15623
rect 20806 15620 20812 15632
rect 20303 15592 20812 15620
rect 20303 15589 20315 15592
rect 20257 15583 20315 15589
rect 20548 15564 20576 15592
rect 20806 15580 20812 15592
rect 20864 15580 20870 15632
rect 21266 15580 21272 15632
rect 21324 15620 21330 15632
rect 26421 15623 26479 15629
rect 26421 15620 26433 15623
rect 21324 15592 26433 15620
rect 21324 15580 21330 15592
rect 26421 15589 26433 15592
rect 26467 15620 26479 15623
rect 26602 15620 26608 15632
rect 26467 15592 26608 15620
rect 26467 15589 26479 15592
rect 26421 15583 26479 15589
rect 26602 15580 26608 15592
rect 26660 15580 26666 15632
rect 27632 15629 27660 15660
rect 28258 15648 28264 15660
rect 28316 15648 28322 15700
rect 29086 15648 29092 15700
rect 29144 15688 29150 15700
rect 29270 15688 29276 15700
rect 29144 15660 29276 15688
rect 29144 15648 29150 15660
rect 29270 15648 29276 15660
rect 29328 15648 29334 15700
rect 27617 15623 27675 15629
rect 27617 15589 27629 15623
rect 27663 15589 27675 15623
rect 28813 15623 28871 15629
rect 28813 15620 28825 15623
rect 27617 15583 27675 15589
rect 28276 15592 28825 15620
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15521 16635 15555
rect 16577 15515 16635 15521
rect 16850 15512 16856 15564
rect 16908 15512 16914 15564
rect 16942 15512 16948 15564
rect 17000 15552 17006 15564
rect 17109 15555 17167 15561
rect 17109 15552 17121 15555
rect 17000 15524 17121 15552
rect 17000 15512 17006 15524
rect 17109 15521 17121 15524
rect 17155 15521 17167 15555
rect 17109 15515 17167 15521
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 18012 15524 18521 15552
rect 18012 15512 18018 15524
rect 18509 15521 18521 15524
rect 18555 15521 18567 15555
rect 18509 15515 18567 15521
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15552 18935 15555
rect 19337 15555 19395 15561
rect 19337 15552 19349 15555
rect 18923 15524 19349 15552
rect 18923 15521 18935 15524
rect 18877 15515 18935 15521
rect 19337 15521 19349 15524
rect 19383 15521 19395 15555
rect 19337 15515 19395 15521
rect 18414 15444 18420 15496
rect 18472 15444 18478 15496
rect 19352 15484 19380 15515
rect 19518 15512 19524 15564
rect 19576 15512 19582 15564
rect 19794 15512 19800 15564
rect 19852 15512 19858 15564
rect 20530 15512 20536 15564
rect 20588 15512 20594 15564
rect 20714 15512 20720 15564
rect 20772 15512 20778 15564
rect 20990 15512 20996 15564
rect 21048 15512 21054 15564
rect 21450 15512 21456 15564
rect 21508 15512 21514 15564
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15521 21695 15555
rect 21637 15515 21695 15521
rect 19610 15484 19616 15496
rect 19352 15456 19616 15484
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15484 20499 15487
rect 21652 15484 21680 15515
rect 21818 15512 21824 15564
rect 21876 15512 21882 15564
rect 22094 15512 22100 15564
rect 22152 15512 22158 15564
rect 22833 15555 22891 15561
rect 22833 15521 22845 15555
rect 22879 15552 22891 15555
rect 23382 15552 23388 15564
rect 22879 15524 23388 15552
rect 22879 15521 22891 15524
rect 22833 15515 22891 15521
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 24029 15555 24087 15561
rect 24029 15521 24041 15555
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 24213 15555 24271 15561
rect 24213 15521 24225 15555
rect 24259 15552 24271 15555
rect 24486 15552 24492 15564
rect 24259 15524 24492 15552
rect 24259 15521 24271 15524
rect 24213 15515 24271 15521
rect 23290 15484 23296 15496
rect 20487 15456 23296 15484
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 23290 15444 23296 15456
rect 23348 15484 23354 15496
rect 24044 15484 24072 15515
rect 24486 15512 24492 15524
rect 24544 15512 24550 15564
rect 24854 15512 24860 15564
rect 24912 15512 24918 15564
rect 25225 15555 25283 15561
rect 25225 15521 25237 15555
rect 25271 15521 25283 15555
rect 25225 15515 25283 15521
rect 23348 15456 24072 15484
rect 23348 15444 23354 15456
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 24670 15484 24676 15496
rect 24452 15456 24676 15484
rect 24452 15444 24458 15456
rect 24670 15444 24676 15456
rect 24728 15484 24734 15496
rect 25240 15484 25268 15515
rect 25774 15512 25780 15564
rect 25832 15552 25838 15564
rect 26145 15555 26203 15561
rect 26145 15552 26157 15555
rect 25832 15524 26157 15552
rect 25832 15512 25838 15524
rect 26145 15521 26157 15524
rect 26191 15552 26203 15555
rect 27157 15555 27215 15561
rect 27157 15552 27169 15555
rect 26191 15524 27169 15552
rect 26191 15521 26203 15524
rect 26145 15515 26203 15521
rect 27157 15521 27169 15524
rect 27203 15521 27215 15555
rect 27157 15515 27215 15521
rect 27801 15555 27859 15561
rect 27801 15521 27813 15555
rect 27847 15521 27859 15555
rect 27801 15515 27859 15521
rect 24728 15456 25268 15484
rect 27816 15484 27844 15515
rect 27982 15512 27988 15564
rect 28040 15552 28046 15564
rect 28276 15561 28304 15592
rect 28813 15589 28825 15592
rect 28859 15589 28871 15623
rect 28813 15583 28871 15589
rect 28169 15555 28227 15561
rect 28169 15552 28181 15555
rect 28040 15524 28181 15552
rect 28040 15512 28046 15524
rect 28169 15521 28181 15524
rect 28215 15521 28227 15555
rect 28169 15515 28227 15521
rect 28261 15555 28319 15561
rect 28261 15521 28273 15555
rect 28307 15521 28319 15555
rect 28261 15515 28319 15521
rect 28442 15512 28448 15564
rect 28500 15512 28506 15564
rect 28537 15555 28595 15561
rect 28537 15521 28549 15555
rect 28583 15552 28595 15555
rect 28994 15552 29000 15564
rect 28583 15524 29000 15552
rect 28583 15521 28595 15524
rect 28537 15515 28595 15521
rect 28994 15512 29000 15524
rect 29052 15512 29058 15564
rect 29086 15512 29092 15564
rect 29144 15512 29150 15564
rect 29178 15512 29184 15564
rect 29236 15512 29242 15564
rect 29270 15512 29276 15564
rect 29328 15561 29334 15564
rect 29328 15552 29336 15561
rect 29328 15524 29373 15552
rect 29328 15515 29336 15524
rect 29328 15512 29334 15515
rect 29454 15512 29460 15564
rect 29512 15512 29518 15564
rect 27816 15456 28994 15484
rect 24728 15444 24734 15456
rect 19058 15376 19064 15428
rect 19116 15416 19122 15428
rect 20622 15416 20628 15428
rect 19116 15388 20628 15416
rect 19116 15376 19122 15388
rect 20622 15376 20628 15388
rect 20680 15416 20686 15428
rect 21269 15419 21327 15425
rect 21269 15416 21281 15419
rect 20680 15388 21281 15416
rect 20680 15376 20686 15388
rect 21269 15385 21281 15388
rect 21315 15385 21327 15419
rect 21269 15379 21327 15385
rect 21634 15376 21640 15428
rect 21692 15416 21698 15428
rect 22738 15416 22744 15428
rect 21692 15388 22744 15416
rect 21692 15376 21698 15388
rect 22738 15376 22744 15388
rect 22796 15376 22802 15428
rect 28966 15416 28994 15456
rect 29086 15416 29092 15428
rect 28966 15388 29092 15416
rect 29086 15376 29092 15388
rect 29144 15376 29150 15428
rect 16485 15351 16543 15357
rect 16485 15348 16497 15351
rect 15620 15320 16497 15348
rect 15620 15308 15626 15320
rect 16485 15317 16497 15320
rect 16531 15317 16543 15351
rect 16485 15311 16543 15317
rect 16666 15308 16672 15360
rect 16724 15348 16730 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 16724 15320 18797 15348
rect 16724 15308 16730 15320
rect 18785 15317 18797 15320
rect 18831 15348 18843 15351
rect 19705 15351 19763 15357
rect 19705 15348 19717 15351
rect 18831 15320 19717 15348
rect 18831 15317 18843 15320
rect 18785 15311 18843 15317
rect 19705 15317 19717 15320
rect 19751 15348 19763 15351
rect 20806 15348 20812 15360
rect 19751 15320 20812 15348
rect 19751 15317 19763 15320
rect 19705 15311 19763 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 21450 15308 21456 15360
rect 21508 15348 21514 15360
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 21508 15320 21925 15348
rect 21508 15308 21514 15320
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 24397 15351 24455 15357
rect 24397 15317 24409 15351
rect 24443 15348 24455 15351
rect 24578 15348 24584 15360
rect 24443 15320 24584 15348
rect 24443 15317 24455 15320
rect 24397 15311 24455 15317
rect 24578 15308 24584 15320
rect 24636 15308 24642 15360
rect 25406 15308 25412 15360
rect 25464 15348 25470 15360
rect 25501 15351 25559 15357
rect 25501 15348 25513 15351
rect 25464 15320 25513 15348
rect 25464 15308 25470 15320
rect 25501 15317 25513 15320
rect 25547 15348 25559 15351
rect 25682 15348 25688 15360
rect 25547 15320 25688 15348
rect 25547 15317 25559 15320
rect 25501 15311 25559 15317
rect 25682 15308 25688 15320
rect 25740 15308 25746 15360
rect 27985 15351 28043 15357
rect 27985 15317 27997 15351
rect 28031 15348 28043 15351
rect 28534 15348 28540 15360
rect 28031 15320 28540 15348
rect 28031 15317 28043 15320
rect 27985 15311 28043 15317
rect 28534 15308 28540 15320
rect 28592 15308 28598 15360
rect 28721 15351 28779 15357
rect 28721 15317 28733 15351
rect 28767 15348 28779 15351
rect 30650 15348 30656 15360
rect 28767 15320 30656 15348
rect 28767 15317 28779 15320
rect 28721 15311 28779 15317
rect 30650 15308 30656 15320
rect 30708 15308 30714 15360
rect 552 15258 31648 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 11436 15258
rect 11488 15206 11500 15258
rect 11552 15206 11564 15258
rect 11616 15206 11628 15258
rect 11680 15206 11692 15258
rect 11744 15206 19210 15258
rect 19262 15206 19274 15258
rect 19326 15206 19338 15258
rect 19390 15206 19402 15258
rect 19454 15206 19466 15258
rect 19518 15206 26984 15258
rect 27036 15206 27048 15258
rect 27100 15206 27112 15258
rect 27164 15206 27176 15258
rect 27228 15206 27240 15258
rect 27292 15206 31648 15258
rect 552 15184 31648 15206
rect 4890 15144 4896 15156
rect 2746 15116 4896 15144
rect 2746 15008 2774 15116
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 5445 15147 5503 15153
rect 5445 15113 5457 15147
rect 5491 15144 5503 15147
rect 5534 15144 5540 15156
rect 5491 15116 5540 15144
rect 5491 15113 5503 15116
rect 5445 15107 5503 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 5684 15116 8064 15144
rect 5684 15104 5690 15116
rect 4706 15036 4712 15088
rect 4764 15076 4770 15088
rect 6273 15079 6331 15085
rect 6273 15076 6285 15079
rect 4764 15048 6285 15076
rect 4764 15036 4770 15048
rect 6273 15045 6285 15048
rect 6319 15045 6331 15079
rect 6273 15039 6331 15045
rect 2516 14980 2774 15008
rect 1578 14900 1584 14952
rect 1636 14940 1642 14952
rect 1946 14940 1952 14952
rect 1636 14912 1952 14940
rect 1636 14900 1642 14912
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 2516 14949 2544 14980
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4801 15011 4859 15017
rect 4212 14980 4384 15008
rect 4212 14968 4218 14980
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14909 2559 14943
rect 2501 14903 2559 14909
rect 2590 14900 2596 14952
rect 2648 14900 2654 14952
rect 2685 14943 2743 14949
rect 2685 14909 2697 14943
rect 2731 14940 2743 14943
rect 2774 14940 2780 14952
rect 2731 14912 2780 14940
rect 2731 14909 2743 14912
rect 2685 14903 2743 14909
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14909 2927 14943
rect 2869 14903 2927 14909
rect 2884 14872 2912 14903
rect 3050 14900 3056 14952
rect 3108 14940 3114 14952
rect 3234 14940 3240 14952
rect 3108 14912 3240 14940
rect 3108 14900 3114 14912
rect 3234 14900 3240 14912
rect 3292 14900 3298 14952
rect 4356 14949 4384 14980
rect 4801 14977 4813 15011
rect 4847 15008 4859 15011
rect 5534 15008 5540 15020
rect 4847 14980 5540 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 5534 14968 5540 14980
rect 5592 14968 5598 15020
rect 6089 15011 6147 15017
rect 6089 14977 6101 15011
rect 6135 14977 6147 15011
rect 6089 14971 6147 14977
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5905 14943 5963 14949
rect 5905 14940 5917 14943
rect 5399 14912 5917 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 5905 14909 5917 14912
rect 5951 14909 5963 14943
rect 6104 14940 6132 14971
rect 6730 14968 6736 15020
rect 6788 14968 6794 15020
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 6840 14940 6868 14971
rect 7190 14940 7196 14952
rect 6104 14912 7196 14940
rect 5905 14903 5963 14909
rect 3418 14872 3424 14884
rect 2884 14844 3424 14872
rect 3418 14832 3424 14844
rect 3476 14832 3482 14884
rect 3881 14875 3939 14881
rect 3881 14841 3893 14875
rect 3927 14872 3939 14875
rect 4157 14875 4215 14881
rect 4157 14872 4169 14875
rect 3927 14844 4169 14872
rect 3927 14841 3939 14844
rect 3881 14835 3939 14841
rect 4157 14841 4169 14844
rect 4203 14841 4215 14875
rect 4632 14872 4660 14903
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 8036 14949 8064 15116
rect 9582 15104 9588 15156
rect 9640 15144 9646 15156
rect 9953 15147 10011 15153
rect 9640 15116 9812 15144
rect 9640 15104 9646 15116
rect 9784 15085 9812 15116
rect 9953 15113 9965 15147
rect 9999 15144 10011 15147
rect 10318 15144 10324 15156
rect 9999 15116 10324 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 10468 15116 11652 15144
rect 10468 15104 10474 15116
rect 9769 15079 9827 15085
rect 9769 15045 9781 15079
rect 9815 15045 9827 15079
rect 9769 15039 9827 15045
rect 10042 15036 10048 15088
rect 10100 15036 10106 15088
rect 10336 15076 10364 15104
rect 11624 15076 11652 15116
rect 13722 15104 13728 15156
rect 13780 15144 13786 15156
rect 15286 15144 15292 15156
rect 13780 15116 15292 15144
rect 13780 15104 13786 15116
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 15378 15104 15384 15156
rect 15436 15104 15442 15156
rect 16390 15104 16396 15156
rect 16448 15104 16454 15156
rect 16574 15104 16580 15156
rect 16632 15144 16638 15156
rect 21266 15144 21272 15156
rect 16632 15116 21272 15144
rect 16632 15104 16638 15116
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 25958 15144 25964 15156
rect 24136 15116 25964 15144
rect 24136 15088 24164 15116
rect 25958 15104 25964 15116
rect 26016 15144 26022 15156
rect 26694 15144 26700 15156
rect 26016 15116 26700 15144
rect 26016 15104 26022 15116
rect 26694 15104 26700 15116
rect 26752 15104 26758 15156
rect 28994 15104 29000 15156
rect 29052 15144 29058 15156
rect 29089 15147 29147 15153
rect 29089 15144 29101 15147
rect 29052 15116 29101 15144
rect 29052 15104 29058 15116
rect 29089 15113 29101 15116
rect 29135 15113 29147 15147
rect 29089 15107 29147 15113
rect 29454 15104 29460 15156
rect 29512 15144 29518 15156
rect 30285 15147 30343 15153
rect 30285 15144 30297 15147
rect 29512 15116 30297 15144
rect 29512 15104 29518 15116
rect 30285 15113 30297 15116
rect 30331 15113 30343 15147
rect 30285 15107 30343 15113
rect 10336 15048 11560 15076
rect 11624 15048 11836 15076
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9088 14980 9628 15008
rect 9088 14968 9094 14980
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14909 8263 14943
rect 8205 14903 8263 14909
rect 6178 14872 6184 14884
rect 4632 14844 6184 14872
rect 4157 14835 4215 14841
rect 6178 14832 6184 14844
rect 6236 14832 6242 14884
rect 6914 14872 6920 14884
rect 6564 14844 6920 14872
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 1857 14807 1915 14813
rect 1857 14804 1869 14807
rect 1728 14776 1869 14804
rect 1728 14764 1734 14776
rect 1857 14773 1869 14776
rect 1903 14773 1915 14807
rect 1857 14767 1915 14773
rect 2222 14764 2228 14816
rect 2280 14764 2286 14816
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3660 14776 3985 14804
rect 3660 14764 3666 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 3973 14767 4031 14773
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 4525 14807 4583 14813
rect 4525 14804 4537 14807
rect 4304 14776 4537 14804
rect 4304 14764 4310 14776
rect 4525 14773 4537 14776
rect 4571 14773 4583 14807
rect 4525 14767 4583 14773
rect 5813 14807 5871 14813
rect 5813 14773 5825 14807
rect 5859 14804 5871 14807
rect 6564 14804 6592 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7208 14872 7236 14900
rect 8113 14875 8171 14881
rect 8113 14872 8125 14875
rect 7208 14844 8125 14872
rect 8113 14841 8125 14844
rect 8159 14841 8171 14875
rect 8220 14872 8248 14903
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 9490 14940 9496 14952
rect 8352 14912 9496 14940
rect 8352 14900 8358 14912
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9600 14940 9628 14980
rect 9858 14968 9864 15020
rect 9916 15008 9922 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 9916 14980 10517 15008
rect 9916 14968 9922 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 11532 15017 11560 15048
rect 11517 15011 11575 15017
rect 10744 14980 11100 15008
rect 10744 14968 10750 14980
rect 10134 14940 10140 14952
rect 9600 14912 10140 14940
rect 10134 14900 10140 14912
rect 10192 14940 10198 14952
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 10192 14912 10241 14940
rect 10192 14900 10198 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 10428 14872 10456 14903
rect 10594 14900 10600 14952
rect 10652 14900 10658 14952
rect 10781 14943 10839 14949
rect 10781 14909 10793 14943
rect 10827 14940 10839 14943
rect 10870 14940 10876 14952
rect 10827 14912 10876 14940
rect 10827 14909 10839 14912
rect 10781 14903 10839 14909
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 10962 14900 10968 14952
rect 11020 14900 11026 14952
rect 11072 14940 11100 14980
rect 11517 14977 11529 15011
rect 11563 15008 11575 15011
rect 11609 15011 11667 15017
rect 11609 15008 11621 15011
rect 11563 14980 11621 15008
rect 11563 14977 11575 14980
rect 11517 14971 11575 14977
rect 11609 14977 11621 14980
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 11808 14949 11836 15048
rect 15838 15036 15844 15088
rect 15896 15076 15902 15088
rect 16025 15079 16083 15085
rect 16025 15076 16037 15079
rect 15896 15048 16037 15076
rect 15896 15036 15902 15048
rect 16025 15045 16037 15048
rect 16071 15045 16083 15079
rect 16025 15039 16083 15045
rect 16669 15079 16727 15085
rect 16669 15045 16681 15079
rect 16715 15076 16727 15079
rect 16942 15076 16948 15088
rect 16715 15048 16948 15076
rect 16715 15045 16727 15048
rect 16669 15039 16727 15045
rect 16942 15036 16948 15048
rect 17000 15036 17006 15088
rect 18417 15079 18475 15085
rect 18417 15045 18429 15079
rect 18463 15076 18475 15079
rect 19610 15076 19616 15088
rect 18463 15048 19616 15076
rect 18463 15045 18475 15048
rect 18417 15039 18475 15045
rect 19610 15036 19616 15048
rect 19668 15036 19674 15088
rect 20714 15036 20720 15088
rect 20772 15076 20778 15088
rect 21177 15079 21235 15085
rect 21177 15076 21189 15079
rect 20772 15048 21189 15076
rect 20772 15036 20778 15048
rect 21177 15045 21189 15048
rect 21223 15076 21235 15079
rect 21910 15076 21916 15088
rect 21223 15048 21916 15076
rect 21223 15045 21235 15048
rect 21177 15039 21235 15045
rect 21910 15036 21916 15048
rect 21968 15076 21974 15088
rect 22373 15079 22431 15085
rect 21968 15048 22094 15076
rect 21968 15036 21974 15048
rect 13998 14968 14004 15020
rect 14056 14968 14062 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15436 14980 16436 15008
rect 15436 14968 15442 14980
rect 11333 14943 11391 14949
rect 11333 14940 11345 14943
rect 11072 14912 11345 14940
rect 11333 14909 11345 14912
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13630 14940 13636 14952
rect 13228 14912 13636 14940
rect 13228 14900 13234 14912
rect 13630 14900 13636 14912
rect 13688 14900 13694 14952
rect 15746 14900 15752 14952
rect 15804 14900 15810 14952
rect 16408 14949 16436 14980
rect 16482 14968 16488 15020
rect 16540 15008 16546 15020
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 16540 14980 17080 15008
rect 16540 14968 16546 14980
rect 16025 14943 16083 14949
rect 16025 14909 16037 14943
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 16393 14943 16451 14949
rect 16393 14909 16405 14943
rect 16439 14909 16451 14943
rect 16393 14903 16451 14909
rect 16577 14943 16635 14949
rect 16577 14909 16589 14943
rect 16623 14940 16635 14943
rect 16850 14940 16856 14952
rect 16623 14912 16856 14940
rect 16623 14909 16635 14912
rect 16577 14903 16635 14909
rect 10502 14872 10508 14884
rect 8220 14844 10508 14872
rect 8113 14835 8171 14841
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 13538 14872 13544 14884
rect 11348 14844 13544 14872
rect 5859 14776 6592 14804
rect 6641 14807 6699 14813
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 7006 14804 7012 14816
rect 6687 14776 7012 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 7156 14776 7297 14804
rect 7156 14764 7162 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 11238 14804 11244 14816
rect 7432 14776 11244 14804
rect 7432 14764 7438 14776
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11348 14813 11376 14844
rect 13538 14832 13544 14844
rect 13596 14832 13602 14884
rect 14268 14875 14326 14881
rect 14268 14841 14280 14875
rect 14314 14872 14326 14875
rect 14366 14872 14372 14884
rect 14314 14844 14372 14872
rect 14314 14841 14326 14844
rect 14268 14835 14326 14841
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14773 11391 14807
rect 11333 14767 11391 14773
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 11977 14807 12035 14813
rect 11977 14804 11989 14807
rect 11940 14776 11989 14804
rect 11940 14764 11946 14776
rect 11977 14773 11989 14776
rect 12023 14773 12035 14807
rect 11977 14767 12035 14773
rect 13817 14807 13875 14813
rect 13817 14773 13829 14807
rect 13863 14804 13875 14807
rect 14090 14804 14096 14816
rect 13863 14776 14096 14804
rect 13863 14773 13875 14776
rect 13817 14767 13875 14773
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 16040 14804 16068 14903
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 16942 14900 16948 14952
rect 17000 14900 17006 14952
rect 17052 14949 17080 14980
rect 17144 14980 17785 15008
rect 17144 14949 17172 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 19334 15008 19340 15020
rect 17773 14971 17831 14977
rect 17880 14980 19340 15008
rect 17037 14943 17095 14949
rect 17037 14909 17049 14943
rect 17083 14909 17095 14943
rect 17037 14903 17095 14909
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17218 14900 17224 14952
rect 17276 14940 17282 14952
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 17276 14912 17325 14940
rect 17276 14900 17282 14912
rect 17313 14909 17325 14912
rect 17359 14940 17371 14943
rect 17359 14912 17540 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 16114 14832 16120 14884
rect 16172 14872 16178 14884
rect 17405 14875 17463 14881
rect 17405 14872 17417 14875
rect 16172 14844 17417 14872
rect 16172 14832 16178 14844
rect 17405 14841 17417 14844
rect 17451 14841 17463 14875
rect 17512 14872 17540 14912
rect 17586 14900 17592 14952
rect 17644 14900 17650 14952
rect 17880 14940 17908 14980
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 22066 15008 22094 15048
rect 22373 15045 22385 15079
rect 22419 15076 22431 15079
rect 22554 15076 22560 15088
rect 22419 15048 22560 15076
rect 22419 15045 22431 15048
rect 22373 15039 22431 15045
rect 22554 15036 22560 15048
rect 22612 15036 22618 15088
rect 22922 15036 22928 15088
rect 22980 15076 22986 15088
rect 22980 15048 23612 15076
rect 22980 15036 22986 15048
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 22066 14980 22293 15008
rect 22281 14977 22293 14980
rect 22327 15008 22339 15011
rect 23584 15008 23612 15048
rect 23658 15036 23664 15088
rect 23716 15076 23722 15088
rect 24118 15076 24124 15088
rect 23716 15048 24124 15076
rect 23716 15036 23722 15048
rect 24118 15036 24124 15048
rect 24176 15036 24182 15088
rect 26786 15076 26792 15088
rect 24320 15048 26792 15076
rect 24320 15008 24348 15048
rect 26786 15036 26792 15048
rect 26844 15036 26850 15088
rect 27154 15036 27160 15088
rect 27212 15076 27218 15088
rect 27430 15076 27436 15088
rect 27212 15048 27436 15076
rect 27212 15036 27218 15048
rect 27430 15036 27436 15048
rect 27488 15036 27494 15088
rect 28350 15036 28356 15088
rect 28408 15076 28414 15088
rect 29270 15076 29276 15088
rect 28408 15048 29276 15076
rect 28408 15036 28414 15048
rect 29270 15036 29276 15048
rect 29328 15076 29334 15088
rect 30558 15076 30564 15088
rect 29328 15048 30564 15076
rect 29328 15036 29334 15048
rect 30558 15036 30564 15048
rect 30616 15036 30622 15088
rect 22327 14980 23244 15008
rect 23584 14980 24348 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 18233 14943 18291 14949
rect 18233 14940 18245 14943
rect 17696 14912 17908 14940
rect 18064 14912 18245 14940
rect 17696 14872 17724 14912
rect 17512 14844 17724 14872
rect 17405 14835 17463 14841
rect 17770 14832 17776 14884
rect 17828 14872 17834 14884
rect 17957 14875 18015 14881
rect 17957 14872 17969 14875
rect 17828 14844 17969 14872
rect 17828 14832 17834 14844
rect 17957 14841 17969 14844
rect 18003 14841 18015 14875
rect 17957 14835 18015 14841
rect 16942 14804 16948 14816
rect 16040 14776 16948 14804
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17862 14764 17868 14816
rect 17920 14804 17926 14816
rect 18064 14813 18092 14912
rect 18233 14909 18245 14912
rect 18279 14909 18291 14943
rect 18233 14903 18291 14909
rect 19610 14900 19616 14952
rect 19668 14940 19674 14952
rect 20993 14943 21051 14949
rect 20993 14940 21005 14943
rect 19668 14912 21005 14940
rect 19668 14900 19674 14912
rect 20993 14909 21005 14912
rect 21039 14940 21051 14943
rect 21542 14940 21548 14952
rect 21039 14912 21548 14940
rect 21039 14909 21051 14912
rect 20993 14903 21051 14909
rect 21542 14900 21548 14912
rect 21600 14900 21606 14952
rect 22002 14900 22008 14952
rect 22060 14900 22066 14952
rect 22649 14943 22707 14949
rect 22649 14909 22661 14943
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 22833 14943 22891 14949
rect 22833 14909 22845 14943
rect 22879 14940 22891 14943
rect 22922 14940 22928 14952
rect 22879 14912 22928 14940
rect 22879 14909 22891 14912
rect 22833 14903 22891 14909
rect 18874 14832 18880 14884
rect 18932 14872 18938 14884
rect 20622 14872 20628 14884
rect 18932 14844 20628 14872
rect 18932 14832 18938 14844
rect 20622 14832 20628 14844
rect 20680 14872 20686 14884
rect 20809 14875 20867 14881
rect 20809 14872 20821 14875
rect 20680 14844 20821 14872
rect 20680 14832 20686 14844
rect 20809 14841 20821 14844
rect 20855 14841 20867 14875
rect 20809 14835 20867 14841
rect 21450 14832 21456 14884
rect 21508 14872 21514 14884
rect 22664 14872 22692 14903
rect 22922 14900 22928 14912
rect 22980 14900 22986 14952
rect 23216 14949 23244 14980
rect 23201 14943 23259 14949
rect 23201 14909 23213 14943
rect 23247 14909 23259 14943
rect 23201 14903 23259 14909
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 24320 14949 24348 14980
rect 24486 14968 24492 15020
rect 24544 15008 24550 15020
rect 26605 15011 26663 15017
rect 26605 15008 26617 15011
rect 24544 14980 26617 15008
rect 24544 14968 24550 14980
rect 26605 14977 26617 14980
rect 26651 15008 26663 15011
rect 26694 15008 26700 15020
rect 26651 14980 26700 15008
rect 26651 14977 26663 14980
rect 26605 14971 26663 14977
rect 26694 14968 26700 14980
rect 26752 14968 26758 15020
rect 28994 14968 29000 15020
rect 29052 15008 29058 15020
rect 29638 15008 29644 15020
rect 29052 14980 29644 15008
rect 29052 14968 29058 14980
rect 29638 14968 29644 14980
rect 29696 14968 29702 15020
rect 29730 14968 29736 15020
rect 29788 15008 29794 15020
rect 29788 14980 30236 15008
rect 29788 14968 29794 14980
rect 24213 14943 24271 14949
rect 24213 14940 24225 14943
rect 24176 14912 24225 14940
rect 24176 14900 24182 14912
rect 24213 14909 24225 14912
rect 24259 14909 24271 14943
rect 24213 14903 24271 14909
rect 24305 14943 24363 14949
rect 24305 14909 24317 14943
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24394 14900 24400 14952
rect 24452 14900 24458 14952
rect 24578 14900 24584 14952
rect 24636 14900 24642 14952
rect 24946 14900 24952 14952
rect 25004 14900 25010 14952
rect 25038 14900 25044 14952
rect 25096 14900 25102 14952
rect 25222 14900 25228 14952
rect 25280 14900 25286 14952
rect 25317 14943 25375 14949
rect 25317 14909 25329 14943
rect 25363 14909 25375 14943
rect 25317 14903 25375 14909
rect 23017 14875 23075 14881
rect 23017 14872 23029 14875
rect 21508 14844 23029 14872
rect 21508 14832 21514 14844
rect 23017 14841 23029 14844
rect 23063 14841 23075 14875
rect 23017 14835 23075 14841
rect 25130 14832 25136 14884
rect 25188 14872 25194 14884
rect 25332 14872 25360 14903
rect 26878 14900 26884 14952
rect 26936 14940 26942 14952
rect 27157 14943 27215 14949
rect 27157 14940 27169 14943
rect 26936 14912 27169 14940
rect 26936 14900 26942 14912
rect 27157 14909 27169 14912
rect 27203 14909 27215 14943
rect 27157 14903 27215 14909
rect 27249 14943 27307 14949
rect 27249 14909 27261 14943
rect 27295 14909 27307 14943
rect 27249 14903 27307 14909
rect 25188 14844 25360 14872
rect 25188 14832 25194 14844
rect 25590 14832 25596 14884
rect 25648 14872 25654 14884
rect 27264 14872 27292 14903
rect 27430 14900 27436 14952
rect 27488 14900 27494 14952
rect 27525 14943 27583 14949
rect 27525 14909 27537 14943
rect 27571 14940 27583 14943
rect 27982 14940 27988 14952
rect 27571 14912 27988 14940
rect 27571 14909 27583 14912
rect 27525 14903 27583 14909
rect 27982 14900 27988 14912
rect 28040 14900 28046 14952
rect 28626 14900 28632 14952
rect 28684 14900 28690 14952
rect 29546 14900 29552 14952
rect 29604 14940 29610 14952
rect 30101 14943 30159 14949
rect 30101 14940 30113 14943
rect 29604 14912 30113 14940
rect 29604 14900 29610 14912
rect 30101 14909 30113 14912
rect 30147 14909 30159 14943
rect 30101 14903 30159 14909
rect 30208 14884 30236 14980
rect 30466 14900 30472 14952
rect 30524 14900 30530 14952
rect 30650 14900 30656 14952
rect 30708 14900 30714 14952
rect 30745 14943 30803 14949
rect 30745 14909 30757 14943
rect 30791 14909 30803 14943
rect 30745 14903 30803 14909
rect 28442 14872 28448 14884
rect 25648 14844 28448 14872
rect 25648 14832 25654 14844
rect 28442 14832 28448 14844
rect 28500 14832 28506 14884
rect 29914 14832 29920 14884
rect 29972 14832 29978 14884
rect 30190 14832 30196 14884
rect 30248 14872 30254 14884
rect 30760 14872 30788 14903
rect 30834 14900 30840 14952
rect 30892 14900 30898 14952
rect 30248 14844 30788 14872
rect 30248 14832 30254 14844
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 17920 14776 18061 14804
rect 17920 14764 17926 14776
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 18049 14767 18107 14773
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 22646 14804 22652 14816
rect 21048 14776 22652 14804
rect 21048 14764 21054 14776
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 23382 14764 23388 14816
rect 23440 14764 23446 14816
rect 23937 14807 23995 14813
rect 23937 14773 23949 14807
rect 23983 14804 23995 14807
rect 24210 14804 24216 14816
rect 23983 14776 24216 14804
rect 23983 14773 23995 14776
rect 23937 14767 23995 14773
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 25498 14764 25504 14816
rect 25556 14764 25562 14816
rect 25866 14764 25872 14816
rect 25924 14804 25930 14816
rect 26053 14807 26111 14813
rect 26053 14804 26065 14807
rect 25924 14776 26065 14804
rect 25924 14764 25930 14776
rect 26053 14773 26065 14776
rect 26099 14773 26111 14807
rect 26053 14767 26111 14773
rect 26973 14807 27031 14813
rect 26973 14773 26985 14807
rect 27019 14804 27031 14807
rect 27246 14804 27252 14816
rect 27019 14776 27252 14804
rect 27019 14773 27031 14776
rect 26973 14767 27031 14773
rect 27246 14764 27252 14776
rect 27304 14764 27310 14816
rect 27522 14764 27528 14816
rect 27580 14804 27586 14816
rect 27985 14807 28043 14813
rect 27985 14804 27997 14807
rect 27580 14776 27997 14804
rect 27580 14764 27586 14776
rect 27985 14773 27997 14776
rect 28031 14773 28043 14807
rect 27985 14767 28043 14773
rect 29086 14764 29092 14816
rect 29144 14804 29150 14816
rect 29270 14804 29276 14816
rect 29144 14776 29276 14804
rect 29144 14764 29150 14776
rect 29270 14764 29276 14776
rect 29328 14804 29334 14816
rect 29457 14807 29515 14813
rect 29457 14804 29469 14807
rect 29328 14776 29469 14804
rect 29328 14764 29334 14776
rect 29457 14773 29469 14776
rect 29503 14773 29515 14807
rect 29457 14767 29515 14773
rect 29822 14764 29828 14816
rect 29880 14804 29886 14816
rect 31113 14807 31171 14813
rect 31113 14804 31125 14807
rect 29880 14776 31125 14804
rect 29880 14764 29886 14776
rect 31113 14773 31125 14776
rect 31159 14773 31171 14807
rect 31113 14767 31171 14773
rect 552 14714 31648 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 12096 14714
rect 12148 14662 12160 14714
rect 12212 14662 12224 14714
rect 12276 14662 12288 14714
rect 12340 14662 12352 14714
rect 12404 14662 19870 14714
rect 19922 14662 19934 14714
rect 19986 14662 19998 14714
rect 20050 14662 20062 14714
rect 20114 14662 20126 14714
rect 20178 14662 27644 14714
rect 27696 14662 27708 14714
rect 27760 14662 27772 14714
rect 27824 14662 27836 14714
rect 27888 14662 27900 14714
rect 27952 14662 31648 14714
rect 552 14640 31648 14662
rect 3418 14560 3424 14612
rect 3476 14560 3482 14612
rect 5534 14560 5540 14612
rect 5592 14560 5598 14612
rect 7098 14560 7104 14612
rect 7156 14560 7162 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 10410 14600 10416 14612
rect 7616 14572 10416 14600
rect 7616 14560 7622 14572
rect 10410 14560 10416 14572
rect 10468 14560 10474 14612
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 10652 14572 11437 14600
rect 10652 14560 10658 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11425 14563 11483 14569
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12710 14600 12716 14612
rect 12299 14572 12716 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 13262 14560 13268 14612
rect 13320 14560 13326 14612
rect 14366 14560 14372 14612
rect 14424 14560 14430 14612
rect 16761 14603 16819 14609
rect 16761 14600 16773 14603
rect 16224 14572 16773 14600
rect 1940 14535 1998 14541
rect 1940 14501 1952 14535
rect 1986 14532 1998 14535
rect 2222 14532 2228 14544
rect 1986 14504 2228 14532
rect 1986 14501 1998 14504
rect 1940 14495 1998 14501
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 3436 14532 3464 14560
rect 4424 14535 4482 14541
rect 3436 14504 3832 14532
rect 1670 14424 1676 14476
rect 1728 14424 1734 14476
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 3053 14331 3111 14337
rect 3053 14297 3065 14331
rect 3099 14328 3111 14331
rect 3234 14328 3240 14340
rect 3099 14300 3240 14328
rect 3099 14297 3111 14300
rect 3053 14291 3111 14297
rect 3234 14288 3240 14300
rect 3292 14288 3298 14340
rect 3142 14220 3148 14272
rect 3200 14220 3206 14272
rect 3436 14260 3464 14427
rect 3510 14424 3516 14476
rect 3568 14424 3574 14476
rect 3602 14424 3608 14476
rect 3660 14424 3666 14476
rect 3804 14473 3832 14504
rect 4424 14501 4436 14535
rect 4470 14532 4482 14535
rect 4982 14532 4988 14544
rect 4470 14504 4988 14532
rect 4470 14501 4482 14504
rect 4424 14495 4482 14501
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 5552 14532 5580 14560
rect 5902 14532 5908 14544
rect 5552 14504 5908 14532
rect 5902 14492 5908 14504
rect 5960 14532 5966 14544
rect 7009 14535 7067 14541
rect 5960 14504 6592 14532
rect 5960 14492 5966 14504
rect 3789 14467 3847 14473
rect 3789 14433 3801 14467
rect 3835 14433 3847 14467
rect 3789 14427 3847 14433
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14464 4215 14467
rect 4246 14464 4252 14476
rect 4203 14436 4252 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 5994 14424 6000 14476
rect 6052 14424 6058 14476
rect 6564 14473 6592 14504
rect 7009 14501 7021 14535
rect 7055 14532 7067 14535
rect 9030 14532 9036 14544
rect 7055 14504 9036 14532
rect 7055 14501 7067 14504
rect 7009 14495 7067 14501
rect 9030 14492 9036 14504
rect 9088 14492 9094 14544
rect 10134 14492 10140 14544
rect 10192 14532 10198 14544
rect 10192 14504 10456 14532
rect 10192 14492 10198 14504
rect 10428 14473 10456 14504
rect 10686 14492 10692 14544
rect 10744 14532 10750 14544
rect 10781 14535 10839 14541
rect 10781 14532 10793 14535
rect 10744 14504 10793 14532
rect 10744 14492 10750 14504
rect 10781 14501 10793 14504
rect 10827 14501 10839 14535
rect 10781 14495 10839 14501
rect 11882 14492 11888 14544
rect 11940 14492 11946 14544
rect 11974 14492 11980 14544
rect 12032 14532 12038 14544
rect 12085 14535 12143 14541
rect 12085 14532 12097 14535
rect 12032 14504 12097 14532
rect 12032 14492 12038 14504
rect 12085 14501 12097 14504
rect 12131 14501 12143 14535
rect 12085 14495 12143 14501
rect 13538 14492 13544 14544
rect 13596 14532 13602 14544
rect 14829 14535 14887 14541
rect 14829 14532 14841 14535
rect 13596 14504 14841 14532
rect 13596 14492 13602 14504
rect 14829 14501 14841 14504
rect 14875 14532 14887 14535
rect 15194 14532 15200 14544
rect 14875 14504 15200 14532
rect 14875 14501 14887 14504
rect 14829 14495 14887 14501
rect 15194 14492 15200 14504
rect 15252 14492 15258 14544
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 10413 14467 10471 14473
rect 7883 14436 10364 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 6914 14396 6920 14408
rect 6411 14368 6920 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 6914 14356 6920 14368
rect 6972 14356 6978 14408
rect 7190 14356 7196 14408
rect 7248 14356 7254 14408
rect 7926 14356 7932 14408
rect 7984 14356 7990 14408
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 10336 14396 10364 14436
rect 10413 14433 10425 14467
rect 10459 14464 10471 14467
rect 10502 14464 10508 14476
rect 10459 14436 10508 14464
rect 10459 14433 10471 14436
rect 10413 14427 10471 14433
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 10870 14464 10876 14476
rect 10643 14436 10876 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11238 14424 11244 14476
rect 11296 14424 11302 14476
rect 11333 14467 11391 14473
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 11606 14464 11612 14476
rect 11379 14436 11612 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 11146 14396 11152 14408
rect 10336 14368 11152 14396
rect 8021 14359 8079 14365
rect 7208 14328 7236 14356
rect 8036 14328 8064 14359
rect 11146 14356 11152 14368
rect 11204 14356 11210 14408
rect 6564 14300 7144 14328
rect 7208 14300 8064 14328
rect 6564 14260 6592 14300
rect 3436 14232 6592 14260
rect 6638 14220 6644 14272
rect 6696 14220 6702 14272
rect 7116 14260 7144 14300
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 11348 14328 11376 14427
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 11701 14467 11759 14473
rect 11701 14433 11713 14467
rect 11747 14464 11759 14467
rect 11900 14464 11928 14492
rect 16224 14476 16252 14572
rect 16761 14569 16773 14572
rect 16807 14569 16819 14603
rect 16761 14563 16819 14569
rect 16776 14532 16804 14563
rect 17310 14560 17316 14612
rect 17368 14600 17374 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 17368 14572 18521 14600
rect 17368 14560 17374 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 19058 14560 19064 14612
rect 19116 14560 19122 14612
rect 19153 14603 19211 14609
rect 19153 14569 19165 14603
rect 19199 14600 19211 14603
rect 20717 14603 20775 14609
rect 20717 14600 20729 14603
rect 19199 14572 20729 14600
rect 19199 14569 19211 14572
rect 19153 14563 19211 14569
rect 20717 14569 20729 14572
rect 20763 14600 20775 14603
rect 21358 14600 21364 14612
rect 20763 14572 21364 14600
rect 20763 14569 20775 14572
rect 20717 14563 20775 14569
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 22370 14560 22376 14612
rect 22428 14600 22434 14612
rect 23566 14600 23572 14612
rect 22428 14572 23572 14600
rect 22428 14560 22434 14572
rect 23566 14560 23572 14572
rect 23624 14560 23630 14612
rect 24486 14560 24492 14612
rect 24544 14560 24550 14612
rect 25038 14560 25044 14612
rect 25096 14600 25102 14612
rect 26326 14600 26332 14612
rect 25096 14572 26332 14600
rect 25096 14560 25102 14572
rect 26326 14560 26332 14572
rect 26384 14560 26390 14612
rect 27154 14600 27160 14612
rect 26528 14572 27160 14600
rect 18414 14532 18420 14544
rect 16776 14504 18420 14532
rect 18414 14492 18420 14504
rect 18472 14492 18478 14544
rect 18524 14504 20852 14532
rect 11747 14436 11928 14464
rect 11747 14433 11759 14436
rect 11701 14427 11759 14433
rect 12802 14424 12808 14476
rect 12860 14464 12866 14476
rect 13081 14467 13139 14473
rect 13081 14464 13093 14467
rect 12860 14436 13093 14464
rect 12860 14424 12866 14436
rect 13081 14433 13093 14436
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 13722 14424 13728 14476
rect 13780 14424 13786 14476
rect 13909 14467 13967 14473
rect 13909 14433 13921 14467
rect 13955 14433 13967 14467
rect 13909 14427 13967 14433
rect 13814 14396 13820 14408
rect 9640 14300 11376 14328
rect 11440 14368 13820 14396
rect 9640 14288 9646 14300
rect 7190 14260 7196 14272
rect 7116 14232 7196 14260
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7466 14220 7472 14272
rect 7524 14220 7530 14272
rect 9950 14220 9956 14272
rect 10008 14260 10014 14272
rect 11440 14260 11468 14368
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 13924 14396 13952 14427
rect 13998 14424 14004 14476
rect 14056 14424 14062 14476
rect 14090 14424 14096 14476
rect 14148 14424 14154 14476
rect 14550 14424 14556 14476
rect 14608 14464 14614 14476
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 14608 14436 14657 14464
rect 14608 14424 14614 14436
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 13924 14368 14473 14396
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14660 14396 14688 14427
rect 16206 14424 16212 14476
rect 16264 14424 16270 14476
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 16356 14436 16589 14464
rect 16356 14424 16362 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 17862 14464 17868 14476
rect 16577 14427 16635 14433
rect 16776 14436 17868 14464
rect 16776 14408 16804 14436
rect 17862 14424 17868 14436
rect 17920 14464 17926 14476
rect 18322 14473 18328 14476
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 17920 14436 18153 14464
rect 17920 14424 17926 14436
rect 18141 14433 18153 14436
rect 18187 14433 18199 14467
rect 18141 14427 18199 14433
rect 18295 14467 18328 14473
rect 18295 14433 18307 14467
rect 18380 14464 18386 14476
rect 18524 14464 18552 14504
rect 20824 14476 20852 14504
rect 21266 14492 21272 14544
rect 21324 14532 21330 14544
rect 21453 14535 21511 14541
rect 21453 14532 21465 14535
rect 21324 14504 21465 14532
rect 21324 14492 21330 14504
rect 21453 14501 21465 14504
rect 21499 14501 21511 14535
rect 24857 14535 24915 14541
rect 24857 14532 24869 14535
rect 21453 14495 21511 14501
rect 23584 14504 24869 14532
rect 18380 14436 18552 14464
rect 18295 14427 18328 14433
rect 18322 14424 18328 14427
rect 18380 14424 18386 14436
rect 18966 14424 18972 14476
rect 19024 14424 19030 14476
rect 19610 14464 19616 14476
rect 19260 14436 19616 14464
rect 16758 14396 16764 14408
rect 14660 14368 16764 14396
rect 14461 14359 14519 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 16908 14368 17601 14396
rect 16908 14356 16914 14368
rect 17589 14365 17601 14368
rect 17635 14396 17647 14399
rect 19260 14396 19288 14436
rect 19610 14424 19616 14436
rect 19668 14424 19674 14476
rect 20533 14467 20591 14473
rect 20533 14433 20545 14467
rect 20579 14433 20591 14467
rect 20533 14427 20591 14433
rect 17635 14368 19288 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19886 14396 19892 14408
rect 19392 14368 19892 14396
rect 19392 14356 19398 14368
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 20548 14396 20576 14427
rect 20806 14424 20812 14476
rect 20864 14424 20870 14476
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21634 14464 21640 14476
rect 20947 14436 21640 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21634 14424 21640 14436
rect 21692 14424 21698 14476
rect 21910 14424 21916 14476
rect 21968 14464 21974 14476
rect 22649 14467 22707 14473
rect 22649 14464 22661 14467
rect 21968 14436 22661 14464
rect 21968 14424 21974 14436
rect 22649 14433 22661 14436
rect 22695 14433 22707 14467
rect 22649 14427 22707 14433
rect 22830 14424 22836 14476
rect 22888 14464 22894 14476
rect 23584 14473 23612 14504
rect 24857 14501 24869 14504
rect 24903 14501 24915 14535
rect 24857 14495 24915 14501
rect 25498 14492 25504 14544
rect 25556 14532 25562 14544
rect 25556 14504 26096 14532
rect 25556 14492 25562 14504
rect 23017 14467 23075 14473
rect 23017 14464 23029 14467
rect 22888 14436 23029 14464
rect 22888 14424 22894 14436
rect 23017 14433 23029 14436
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 23569 14467 23627 14473
rect 23569 14433 23581 14467
rect 23615 14433 23627 14467
rect 23569 14427 23627 14433
rect 23658 14424 23664 14476
rect 23716 14424 23722 14476
rect 23750 14424 23756 14476
rect 23808 14424 23814 14476
rect 23842 14424 23848 14476
rect 23900 14464 23906 14476
rect 23937 14467 23995 14473
rect 23937 14464 23949 14467
rect 23900 14436 23949 14464
rect 23900 14424 23906 14436
rect 23937 14433 23949 14436
rect 23983 14464 23995 14467
rect 24302 14464 24308 14476
rect 23983 14436 24308 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24302 14424 24308 14436
rect 24360 14424 24366 14476
rect 24397 14467 24455 14473
rect 24397 14433 24409 14467
rect 24443 14433 24455 14467
rect 24397 14427 24455 14433
rect 21542 14396 21548 14408
rect 20548 14368 21548 14396
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 22002 14356 22008 14408
rect 22060 14396 22066 14408
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 22060 14368 22201 14396
rect 22060 14356 22066 14368
rect 22189 14365 22201 14368
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 24118 14396 24124 14408
rect 23256 14368 24124 14396
rect 23256 14356 23262 14368
rect 24118 14356 24124 14368
rect 24176 14396 24182 14408
rect 24412 14396 24440 14427
rect 24578 14424 24584 14476
rect 24636 14464 24642 14476
rect 24762 14464 24768 14476
rect 24636 14436 24768 14464
rect 24636 14424 24642 14436
rect 24762 14424 24768 14436
rect 24820 14464 24826 14476
rect 25222 14464 25228 14476
rect 24820 14436 25228 14464
rect 24820 14424 24826 14436
rect 25222 14424 25228 14436
rect 25280 14424 25286 14476
rect 25866 14424 25872 14476
rect 25924 14424 25930 14476
rect 25958 14424 25964 14476
rect 26016 14424 26022 14476
rect 26068 14473 26096 14504
rect 26053 14467 26111 14473
rect 26053 14433 26065 14467
rect 26099 14433 26111 14467
rect 26053 14427 26111 14433
rect 26142 14424 26148 14476
rect 26200 14464 26206 14476
rect 26237 14467 26295 14473
rect 26237 14464 26249 14467
rect 26200 14436 26249 14464
rect 26200 14424 26206 14436
rect 26237 14433 26249 14436
rect 26283 14464 26295 14467
rect 26528 14464 26556 14572
rect 27154 14560 27160 14572
rect 27212 14560 27218 14612
rect 27430 14560 27436 14612
rect 27488 14600 27494 14612
rect 27893 14603 27951 14609
rect 27893 14600 27905 14603
rect 27488 14572 27905 14600
rect 27488 14560 27494 14572
rect 27893 14569 27905 14572
rect 27939 14569 27951 14603
rect 27893 14563 27951 14569
rect 29362 14560 29368 14612
rect 29420 14600 29426 14612
rect 30926 14600 30932 14612
rect 29420 14572 30932 14600
rect 29420 14560 29426 14572
rect 30926 14560 30932 14572
rect 30984 14560 30990 14612
rect 26602 14492 26608 14544
rect 26660 14532 26666 14544
rect 29178 14532 29184 14544
rect 26660 14504 27476 14532
rect 26660 14492 26666 14504
rect 26283 14436 26556 14464
rect 26697 14467 26755 14473
rect 26283 14433 26295 14436
rect 26237 14427 26295 14433
rect 26697 14433 26709 14467
rect 26743 14433 26755 14467
rect 26697 14427 26755 14433
rect 24176 14368 24440 14396
rect 24176 14356 24182 14368
rect 24670 14356 24676 14408
rect 24728 14356 24734 14408
rect 25409 14399 25467 14405
rect 25409 14365 25421 14399
rect 25455 14396 25467 14399
rect 26712 14396 26740 14427
rect 26786 14424 26792 14476
rect 26844 14424 26850 14476
rect 26881 14467 26939 14473
rect 26881 14433 26893 14467
rect 26927 14464 26939 14467
rect 26970 14464 26976 14476
rect 26927 14436 26976 14464
rect 26927 14433 26939 14436
rect 26881 14427 26939 14433
rect 26970 14424 26976 14436
rect 27028 14424 27034 14476
rect 27065 14467 27123 14473
rect 27065 14433 27077 14467
rect 27111 14433 27123 14467
rect 27065 14427 27123 14433
rect 25455 14368 26740 14396
rect 25455 14365 25467 14368
rect 25409 14359 25467 14365
rect 11606 14288 11612 14340
rect 11664 14328 11670 14340
rect 15746 14328 15752 14340
rect 11664 14300 15752 14328
rect 11664 14288 11670 14300
rect 15746 14288 15752 14300
rect 15804 14288 15810 14340
rect 16942 14288 16948 14340
rect 17000 14328 17006 14340
rect 17402 14328 17408 14340
rect 17000 14300 17408 14328
rect 17000 14288 17006 14300
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 17957 14331 18015 14337
rect 17957 14297 17969 14331
rect 18003 14297 18015 14331
rect 17957 14291 18015 14297
rect 18049 14331 18107 14337
rect 18049 14297 18061 14331
rect 18095 14328 18107 14331
rect 22094 14328 22100 14340
rect 18095 14300 22100 14328
rect 18095 14297 18107 14300
rect 18049 14291 18107 14297
rect 10008 14232 11468 14260
rect 12069 14263 12127 14269
rect 10008 14220 10014 14232
rect 12069 14229 12081 14263
rect 12115 14260 12127 14263
rect 12710 14260 12716 14272
rect 12115 14232 12716 14260
rect 12115 14229 12127 14232
rect 12069 14223 12127 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 16206 14260 16212 14272
rect 14240 14232 16212 14260
rect 14240 14220 14246 14232
rect 16206 14220 16212 14232
rect 16264 14260 16270 14272
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 16264 14232 16405 14260
rect 16264 14220 16270 14232
rect 16393 14229 16405 14232
rect 16439 14260 16451 14263
rect 17494 14260 17500 14272
rect 16439 14232 17500 14260
rect 16439 14229 16451 14232
rect 16393 14223 16451 14229
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 17972 14260 18000 14291
rect 22094 14288 22100 14300
rect 22152 14288 22158 14340
rect 25222 14328 25228 14340
rect 22940 14300 25228 14328
rect 18322 14260 18328 14272
rect 17972 14232 18328 14260
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 19058 14220 19064 14272
rect 19116 14220 19122 14272
rect 22462 14220 22468 14272
rect 22520 14220 22526 14272
rect 22940 14269 22968 14300
rect 25222 14288 25228 14300
rect 25280 14328 25286 14340
rect 25424 14328 25452 14359
rect 26142 14328 26148 14340
rect 25280 14300 25452 14328
rect 25486 14300 26148 14328
rect 25280 14288 25286 14300
rect 22925 14263 22983 14269
rect 22925 14229 22937 14263
rect 22971 14229 22983 14263
rect 22925 14223 22983 14229
rect 23290 14220 23296 14272
rect 23348 14220 23354 14272
rect 23934 14220 23940 14272
rect 23992 14260 23998 14272
rect 24029 14263 24087 14269
rect 24029 14260 24041 14263
rect 23992 14232 24041 14260
rect 23992 14220 23998 14232
rect 24029 14229 24041 14232
rect 24075 14229 24087 14263
rect 24029 14223 24087 14229
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 25486 14260 25514 14300
rect 26142 14288 26148 14300
rect 26200 14288 26206 14340
rect 26326 14288 26332 14340
rect 26384 14328 26390 14340
rect 26421 14331 26479 14337
rect 26421 14328 26433 14331
rect 26384 14300 26433 14328
rect 26384 14288 26390 14300
rect 26421 14297 26433 14300
rect 26467 14297 26479 14331
rect 26421 14291 26479 14297
rect 26786 14288 26792 14340
rect 26844 14328 26850 14340
rect 27080 14328 27108 14427
rect 27154 14424 27160 14476
rect 27212 14424 27218 14476
rect 27246 14424 27252 14476
rect 27304 14464 27310 14476
rect 27448 14473 27476 14504
rect 28276 14504 29184 14532
rect 28276 14476 28304 14504
rect 29178 14492 29184 14504
rect 29236 14492 29242 14544
rect 29288 14504 30880 14532
rect 27341 14467 27399 14473
rect 27341 14464 27353 14467
rect 27304 14436 27353 14464
rect 27304 14424 27310 14436
rect 27341 14433 27353 14436
rect 27387 14433 27399 14467
rect 27341 14427 27399 14433
rect 27433 14467 27491 14473
rect 27433 14433 27445 14467
rect 27479 14433 27491 14467
rect 27433 14427 27491 14433
rect 27522 14424 27528 14476
rect 27580 14424 27586 14476
rect 27798 14424 27804 14476
rect 27856 14464 27862 14476
rect 28169 14467 28227 14473
rect 28169 14464 28181 14467
rect 27856 14436 28181 14464
rect 27856 14424 27862 14436
rect 28169 14433 28181 14436
rect 28215 14433 28227 14467
rect 28169 14427 28227 14433
rect 28258 14424 28264 14476
rect 28316 14424 28322 14476
rect 28350 14424 28356 14476
rect 28408 14424 28414 14476
rect 28534 14424 28540 14476
rect 28592 14424 28598 14476
rect 28626 14424 28632 14476
rect 28684 14464 28690 14476
rect 29288 14473 29316 14504
rect 29273 14467 29331 14473
rect 29273 14464 29285 14467
rect 28684 14436 29285 14464
rect 28684 14424 28690 14436
rect 29273 14433 29285 14436
rect 29319 14433 29331 14467
rect 29273 14427 29331 14433
rect 29380 14436 30420 14464
rect 27172 14396 27200 14424
rect 27890 14396 27896 14408
rect 27172 14368 27896 14396
rect 27890 14356 27896 14368
rect 27948 14356 27954 14408
rect 28994 14396 29000 14408
rect 28276 14368 29000 14396
rect 26844 14300 27108 14328
rect 27801 14331 27859 14337
rect 26844 14288 26850 14300
rect 27801 14297 27813 14331
rect 27847 14328 27859 14331
rect 27982 14328 27988 14340
rect 27847 14300 27988 14328
rect 27847 14297 27859 14300
rect 27801 14291 27859 14297
rect 27982 14288 27988 14300
rect 28040 14288 28046 14340
rect 24360 14232 25514 14260
rect 24360 14220 24366 14232
rect 25590 14220 25596 14272
rect 25648 14220 25654 14272
rect 25682 14220 25688 14272
rect 25740 14260 25746 14272
rect 27706 14260 27712 14272
rect 25740 14232 27712 14260
rect 25740 14220 25746 14232
rect 27706 14220 27712 14232
rect 27764 14260 27770 14272
rect 28276 14260 28304 14368
rect 28994 14356 29000 14368
rect 29052 14356 29058 14408
rect 29178 14356 29184 14408
rect 29236 14396 29242 14408
rect 29380 14396 29408 14436
rect 29236 14368 29408 14396
rect 29549 14399 29607 14405
rect 29236 14356 29242 14368
rect 29549 14365 29561 14399
rect 29595 14396 29607 14399
rect 29638 14396 29644 14408
rect 29595 14368 29644 14396
rect 29595 14365 29607 14368
rect 29549 14359 29607 14365
rect 29638 14356 29644 14368
rect 29696 14356 29702 14408
rect 30285 14399 30343 14405
rect 30285 14365 30297 14399
rect 30331 14365 30343 14399
rect 30392 14396 30420 14436
rect 30466 14424 30472 14476
rect 30524 14424 30530 14476
rect 30558 14424 30564 14476
rect 30616 14464 30622 14476
rect 30852 14473 30880 14504
rect 30653 14467 30711 14473
rect 30653 14464 30665 14467
rect 30616 14436 30665 14464
rect 30616 14424 30622 14436
rect 30653 14433 30665 14436
rect 30699 14433 30711 14467
rect 30653 14427 30711 14433
rect 30745 14467 30803 14473
rect 30745 14433 30757 14467
rect 30791 14433 30803 14467
rect 30745 14427 30803 14433
rect 30837 14467 30895 14473
rect 30837 14433 30849 14467
rect 30883 14433 30895 14467
rect 30837 14427 30895 14433
rect 30760 14396 30788 14427
rect 30392 14368 30788 14396
rect 30285 14359 30343 14365
rect 29270 14288 29276 14340
rect 29328 14328 29334 14340
rect 30300 14328 30328 14359
rect 29328 14300 30328 14328
rect 29328 14288 29334 14300
rect 27764 14232 28304 14260
rect 28905 14263 28963 14269
rect 27764 14220 27770 14232
rect 28905 14229 28917 14263
rect 28951 14260 28963 14263
rect 28994 14260 29000 14272
rect 28951 14232 29000 14260
rect 28951 14229 28963 14232
rect 28905 14223 28963 14229
rect 28994 14220 29000 14232
rect 29052 14220 29058 14272
rect 29086 14220 29092 14272
rect 29144 14260 29150 14272
rect 29733 14263 29791 14269
rect 29733 14260 29745 14263
rect 29144 14232 29745 14260
rect 29144 14220 29150 14232
rect 29733 14229 29745 14232
rect 29779 14229 29791 14263
rect 29733 14223 29791 14229
rect 30098 14220 30104 14272
rect 30156 14260 30162 14272
rect 31113 14263 31171 14269
rect 31113 14260 31125 14263
rect 30156 14232 31125 14260
rect 30156 14220 30162 14232
rect 31113 14229 31125 14232
rect 31159 14229 31171 14263
rect 31113 14223 31171 14229
rect 552 14170 31648 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 11436 14170
rect 11488 14118 11500 14170
rect 11552 14118 11564 14170
rect 11616 14118 11628 14170
rect 11680 14118 11692 14170
rect 11744 14118 19210 14170
rect 19262 14118 19274 14170
rect 19326 14118 19338 14170
rect 19390 14118 19402 14170
rect 19454 14118 19466 14170
rect 19518 14118 26984 14170
rect 27036 14118 27048 14170
rect 27100 14118 27112 14170
rect 27164 14118 27176 14170
rect 27228 14118 27240 14170
rect 27292 14118 31648 14170
rect 552 14096 31648 14118
rect 1946 14056 1952 14068
rect 1412 14028 1952 14056
rect 1412 13861 1440 14028
rect 1946 14016 1952 14028
rect 2004 14056 2010 14068
rect 2004 14028 2636 14056
rect 2004 14016 2010 14028
rect 2608 13988 2636 14028
rect 3050 14016 3056 14068
rect 3108 14016 3114 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5592 14028 5641 14056
rect 5592 14016 5598 14028
rect 5629 14025 5641 14028
rect 5675 14056 5687 14059
rect 5994 14056 6000 14068
rect 5675 14028 6000 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 10652 14028 10916 14056
rect 10652 14016 10658 14028
rect 10888 13988 10916 14028
rect 11238 14016 11244 14068
rect 11296 14056 11302 14068
rect 12069 14059 12127 14065
rect 12069 14056 12081 14059
rect 11296 14028 12081 14056
rect 11296 14016 11302 14028
rect 12069 14025 12081 14028
rect 12115 14025 12127 14059
rect 12069 14019 12127 14025
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14025 12311 14059
rect 15933 14059 15991 14065
rect 12253 14019 12311 14025
rect 13096 14028 15884 14056
rect 11333 13991 11391 13997
rect 11333 13988 11345 13991
rect 2608 13960 4016 13988
rect 10888 13960 11345 13988
rect 3234 13880 3240 13932
rect 3292 13920 3298 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3292 13892 3801 13920
rect 3292 13880 3298 13892
rect 3789 13889 3801 13892
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3988 13920 4016 13960
rect 11333 13957 11345 13960
rect 11379 13957 11391 13991
rect 11333 13951 11391 13957
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 12268 13988 12296 14019
rect 12032 13960 12296 13988
rect 12032 13948 12038 13960
rect 5813 13923 5871 13929
rect 3988 13892 4384 13920
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 1397 13815 1455 13821
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13852 1547 13855
rect 1673 13855 1731 13861
rect 1673 13852 1685 13855
rect 1535 13824 1685 13852
rect 1535 13821 1547 13824
rect 1489 13815 1547 13821
rect 1673 13821 1685 13824
rect 1719 13821 1731 13855
rect 1673 13815 1731 13821
rect 1940 13855 1998 13861
rect 1940 13821 1952 13855
rect 1986 13852 1998 13855
rect 3142 13852 3148 13864
rect 1986 13824 3148 13852
rect 1986 13821 1998 13824
rect 1940 13815 1998 13821
rect 3142 13812 3148 13824
rect 3200 13812 3206 13864
rect 3988 13861 4016 13892
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 4111 13824 4261 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4249 13821 4261 13824
rect 4295 13821 4307 13855
rect 4356 13852 4384 13892
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6273 13923 6331 13929
rect 6273 13920 6285 13923
rect 5859 13892 6285 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6273 13889 6285 13892
rect 6319 13889 6331 13923
rect 6273 13883 6331 13889
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 9953 13923 10011 13929
rect 9953 13920 9965 13923
rect 9815 13892 9965 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 9953 13889 9965 13892
rect 9999 13889 10011 13923
rect 9953 13883 10011 13889
rect 5721 13855 5779 13861
rect 5721 13852 5733 13855
rect 4356 13824 5733 13852
rect 4249 13815 4307 13821
rect 5721 13821 5733 13824
rect 5767 13852 5779 13855
rect 6178 13852 6184 13864
rect 5767 13824 6184 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6540 13855 6598 13861
rect 6540 13821 6552 13855
rect 6586 13852 6598 13855
rect 7466 13852 7472 13864
rect 6586 13824 7472 13852
rect 6586 13821 6598 13824
rect 6540 13815 6598 13821
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 11882 13852 11888 13864
rect 9907 13824 11888 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 12894 13852 12900 13864
rect 12851 13824 12900 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13096 13861 13124 14028
rect 13998 13948 14004 14000
rect 14056 13988 14062 14000
rect 15856 13988 15884 14028
rect 15933 14025 15945 14059
rect 15979 14056 15991 14059
rect 16298 14056 16304 14068
rect 15979 14028 16304 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 16500 14028 18061 14056
rect 16500 13988 16528 14028
rect 18049 14025 18061 14028
rect 18095 14056 18107 14059
rect 18966 14056 18972 14068
rect 18095 14028 18972 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19300 14028 20760 14056
rect 19300 14016 19306 14028
rect 14056 13960 14136 13988
rect 15856 13960 16528 13988
rect 14056 13948 14062 13960
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13852 13323 13855
rect 13446 13852 13452 13864
rect 13311 13824 13452 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13780 13824 13829 13852
rect 13780 13812 13786 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 13998 13812 14004 13864
rect 14056 13812 14062 13864
rect 14108 13861 14136 13960
rect 17770 13948 17776 14000
rect 17828 13988 17834 14000
rect 17865 13991 17923 13997
rect 17865 13988 17877 13991
rect 17828 13960 17877 13988
rect 17828 13948 17834 13960
rect 17865 13957 17877 13960
rect 17911 13957 17923 13991
rect 17865 13951 17923 13957
rect 17954 13948 17960 14000
rect 18012 13988 18018 14000
rect 18012 13960 20668 13988
rect 18012 13948 18018 13960
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 17552 13892 18184 13920
rect 17552 13880 17558 13892
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 4516 13787 4574 13793
rect 4516 13753 4528 13787
rect 4562 13784 4574 13787
rect 4706 13784 4712 13796
rect 4562 13756 4712 13784
rect 4562 13753 4574 13756
rect 4516 13747 4574 13753
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10220 13787 10278 13793
rect 10220 13784 10232 13787
rect 10100 13756 10232 13784
rect 10100 13744 10106 13756
rect 10220 13753 10232 13756
rect 10266 13753 10278 13787
rect 10220 13747 10278 13753
rect 12437 13787 12495 13793
rect 12437 13753 12449 13787
rect 12483 13784 12495 13787
rect 12710 13784 12716 13796
rect 12483 13756 12716 13784
rect 12483 13753 12495 13756
rect 12437 13747 12495 13753
rect 12710 13744 12716 13756
rect 12768 13744 12774 13796
rect 14108 13784 14136 13815
rect 14182 13812 14188 13864
rect 14240 13812 14246 13864
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 15746 13852 15752 13864
rect 14599 13824 15752 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13852 16543 13855
rect 17034 13852 17040 13864
rect 16531 13824 17040 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17954 13812 17960 13864
rect 18012 13812 18018 13864
rect 18156 13861 18184 13892
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 19242 13920 19248 13932
rect 18472 13892 19248 13920
rect 18472 13880 18478 13892
rect 19242 13880 19248 13892
rect 19300 13880 19306 13932
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13852 18199 13855
rect 19794 13852 19800 13864
rect 18187 13824 19800 13852
rect 18187 13821 18199 13824
rect 18141 13815 18199 13821
rect 19794 13812 19800 13824
rect 19852 13852 19858 13864
rect 20640 13861 20668 13960
rect 20732 13932 20760 14028
rect 20990 14016 20996 14068
rect 21048 14016 21054 14068
rect 21634 14016 21640 14068
rect 21692 14056 21698 14068
rect 22830 14056 22836 14068
rect 21692 14028 22836 14056
rect 21692 14016 21698 14028
rect 22830 14016 22836 14028
rect 22888 14016 22894 14068
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 24578 14056 24584 14068
rect 23523 14028 24584 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 24578 14016 24584 14028
rect 24636 14016 24642 14068
rect 25222 14016 25228 14068
rect 25280 14016 25286 14068
rect 26694 14016 26700 14068
rect 26752 14016 26758 14068
rect 26878 14016 26884 14068
rect 26936 14056 26942 14068
rect 27157 14059 27215 14065
rect 27157 14056 27169 14059
rect 26936 14028 27169 14056
rect 26936 14016 26942 14028
rect 27157 14025 27169 14028
rect 27203 14025 27215 14059
rect 29270 14056 29276 14068
rect 27157 14019 27215 14025
rect 27724 14028 29276 14056
rect 22649 13991 22707 13997
rect 22649 13957 22661 13991
rect 22695 13957 22707 13991
rect 22649 13951 22707 13957
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20772 13892 20913 13920
rect 20772 13880 20778 13892
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 22664 13920 22692 13951
rect 23198 13920 23204 13932
rect 22664 13892 23204 13920
rect 20901 13883 20959 13889
rect 20625 13855 20683 13861
rect 19852 13824 20576 13852
rect 19852 13812 19858 13824
rect 14461 13787 14519 13793
rect 14108 13756 14320 13784
rect 3234 13676 3240 13728
rect 3292 13676 3298 13728
rect 6086 13676 6092 13728
rect 6144 13676 6150 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 7653 13719 7711 13725
rect 7653 13716 7665 13719
rect 7524 13688 7665 13716
rect 7524 13676 7530 13688
rect 7653 13685 7665 13688
rect 7699 13716 7711 13719
rect 7926 13716 7932 13728
rect 7699 13688 7932 13716
rect 7699 13685 7711 13688
rect 7653 13679 7711 13685
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12237 13719 12295 13725
rect 12237 13716 12249 13719
rect 11848 13688 12249 13716
rect 11848 13676 11854 13688
rect 12237 13685 12249 13688
rect 12283 13716 12295 13719
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12283 13688 12633 13716
rect 12283 13685 12295 13688
rect 12237 13679 12295 13685
rect 12621 13685 12633 13688
rect 12667 13685 12679 13719
rect 14292 13716 14320 13756
rect 14461 13753 14473 13787
rect 14507 13784 14519 13787
rect 14798 13787 14856 13793
rect 14798 13784 14810 13787
rect 14507 13756 14810 13784
rect 14507 13753 14519 13756
rect 14461 13747 14519 13753
rect 14798 13753 14810 13756
rect 14844 13753 14856 13787
rect 14798 13747 14856 13753
rect 15194 13744 15200 13796
rect 15252 13784 15258 13796
rect 16025 13787 16083 13793
rect 16025 13784 16037 13787
rect 15252 13756 16037 13784
rect 15252 13744 15258 13756
rect 16025 13753 16037 13756
rect 16071 13784 16083 13787
rect 16114 13784 16120 13796
rect 16071 13756 16120 13784
rect 16071 13753 16083 13756
rect 16025 13747 16083 13753
rect 16114 13744 16120 13756
rect 16172 13744 16178 13796
rect 16752 13787 16810 13793
rect 16224 13756 16528 13784
rect 15470 13716 15476 13728
rect 14292 13688 15476 13716
rect 12621 13679 12679 13685
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 15930 13676 15936 13728
rect 15988 13716 15994 13728
rect 16224 13716 16252 13756
rect 15988 13688 16252 13716
rect 15988 13676 15994 13688
rect 16390 13676 16396 13728
rect 16448 13676 16454 13728
rect 16500 13716 16528 13756
rect 16752 13753 16764 13787
rect 16798 13784 16810 13787
rect 16850 13784 16856 13796
rect 16798 13756 16856 13784
rect 16798 13753 16810 13756
rect 16752 13747 16810 13753
rect 16850 13744 16856 13756
rect 16908 13744 16914 13796
rect 20548 13784 20576 13824
rect 20625 13821 20637 13855
rect 20671 13852 20683 13855
rect 20990 13852 20996 13864
rect 20671 13824 20996 13852
rect 20671 13821 20683 13824
rect 20625 13815 20683 13821
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 22278 13852 22284 13864
rect 21315 13824 22284 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22738 13812 22744 13864
rect 22796 13812 22802 13864
rect 22830 13812 22836 13864
rect 22888 13812 22894 13864
rect 23032 13861 23060 13892
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 23290 13880 23296 13932
rect 23348 13920 23354 13932
rect 26712 13920 26740 14016
rect 27724 13988 27752 14028
rect 29270 14016 29276 14028
rect 29328 14016 29334 14068
rect 29365 14059 29423 14065
rect 29365 14025 29377 14059
rect 29411 14056 29423 14059
rect 30466 14056 30472 14068
rect 29411 14028 30472 14056
rect 29411 14025 29423 14028
rect 29365 14019 29423 14025
rect 30466 14016 30472 14028
rect 30524 14016 30530 14068
rect 30926 14016 30932 14068
rect 30984 14016 30990 14068
rect 29178 13988 29184 14000
rect 27632 13960 27752 13988
rect 28368 13960 29184 13988
rect 27632 13929 27660 13960
rect 27617 13923 27675 13929
rect 23348 13892 23796 13920
rect 26712 13892 27568 13920
rect 23348 13880 23354 13892
rect 23017 13855 23075 13861
rect 23017 13821 23029 13855
rect 23063 13821 23075 13855
rect 23017 13815 23075 13821
rect 23566 13812 23572 13864
rect 23624 13852 23630 13864
rect 23661 13855 23719 13861
rect 23661 13852 23673 13855
rect 23624 13824 23673 13852
rect 23624 13812 23630 13824
rect 23661 13821 23673 13824
rect 23707 13821 23719 13855
rect 23661 13815 23719 13821
rect 21082 13784 21088 13796
rect 20548 13756 21088 13784
rect 21082 13744 21088 13756
rect 21140 13744 21146 13796
rect 21536 13787 21594 13793
rect 21536 13753 21548 13787
rect 21582 13784 21594 13787
rect 21726 13784 21732 13796
rect 21582 13756 21732 13784
rect 21582 13753 21594 13756
rect 21536 13747 21594 13753
rect 21726 13744 21732 13756
rect 21784 13744 21790 13796
rect 22186 13744 22192 13796
rect 22244 13784 22250 13796
rect 23201 13787 23259 13793
rect 23201 13784 23213 13787
rect 22244 13756 23213 13784
rect 22244 13744 22250 13756
rect 23201 13753 23213 13756
rect 23247 13753 23259 13787
rect 23768 13784 23796 13892
rect 23845 13855 23903 13861
rect 23845 13821 23857 13855
rect 23891 13852 23903 13855
rect 24854 13852 24860 13864
rect 23891 13824 24860 13852
rect 23891 13821 23903 13824
rect 23845 13815 23903 13821
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25314 13812 25320 13864
rect 25372 13812 25378 13864
rect 25590 13861 25596 13864
rect 25584 13852 25596 13861
rect 25551 13824 25596 13852
rect 25584 13815 25596 13824
rect 25590 13812 25596 13815
rect 25648 13812 25654 13864
rect 26326 13812 26332 13864
rect 26384 13852 26390 13864
rect 26881 13855 26939 13861
rect 26881 13852 26893 13855
rect 26384 13824 26893 13852
rect 26384 13812 26390 13824
rect 26881 13821 26893 13824
rect 26927 13852 26939 13855
rect 27338 13852 27344 13864
rect 26927 13824 27344 13852
rect 26927 13821 26939 13824
rect 26881 13815 26939 13821
rect 27338 13812 27344 13824
rect 27396 13812 27402 13864
rect 27540 13861 27568 13892
rect 27617 13889 27629 13923
rect 27663 13889 27675 13923
rect 27617 13883 27675 13889
rect 27706 13880 27712 13932
rect 27764 13880 27770 13932
rect 27525 13855 27583 13861
rect 27525 13821 27537 13855
rect 27571 13852 27583 13855
rect 27798 13852 27804 13864
rect 27571 13824 27804 13852
rect 27571 13821 27583 13824
rect 27525 13815 27583 13821
rect 27798 13812 27804 13824
rect 27856 13812 27862 13864
rect 27890 13812 27896 13864
rect 27948 13852 27954 13864
rect 28169 13855 28227 13861
rect 28169 13852 28181 13855
rect 27948 13824 28181 13852
rect 27948 13812 27954 13824
rect 28169 13821 28181 13824
rect 28215 13821 28227 13855
rect 28169 13815 28227 13821
rect 28258 13812 28264 13864
rect 28316 13812 28322 13864
rect 28368 13861 28396 13960
rect 29178 13948 29184 13960
rect 29236 13948 29242 14000
rect 28813 13923 28871 13929
rect 28813 13889 28825 13923
rect 28859 13920 28871 13923
rect 29454 13920 29460 13932
rect 28859 13892 29460 13920
rect 28859 13889 28871 13892
rect 28813 13883 28871 13889
rect 29454 13880 29460 13892
rect 29512 13880 29518 13932
rect 28353 13855 28411 13861
rect 28353 13821 28365 13855
rect 28399 13821 28411 13855
rect 28353 13815 28411 13821
rect 28445 13855 28503 13861
rect 28445 13821 28457 13855
rect 28491 13821 28503 13855
rect 28445 13815 28503 13821
rect 28537 13855 28595 13861
rect 28537 13821 28549 13855
rect 28583 13852 28595 13855
rect 29086 13852 29092 13864
rect 28583 13824 29092 13852
rect 28583 13821 28595 13824
rect 28537 13815 28595 13821
rect 24090 13787 24148 13793
rect 24090 13784 24102 13787
rect 23768 13756 24102 13784
rect 23201 13747 23259 13753
rect 24090 13753 24102 13756
rect 24136 13753 24148 13787
rect 28276 13784 28304 13812
rect 28460 13784 28488 13815
rect 29086 13812 29092 13824
rect 29144 13812 29150 13864
rect 29181 13855 29239 13861
rect 29181 13821 29193 13855
rect 29227 13852 29239 13855
rect 29362 13852 29368 13864
rect 29227 13824 29368 13852
rect 29227 13821 29239 13824
rect 29181 13815 29239 13821
rect 29362 13812 29368 13824
rect 29420 13812 29426 13864
rect 29546 13812 29552 13864
rect 29604 13812 29610 13864
rect 29822 13861 29828 13864
rect 29816 13852 29828 13861
rect 29783 13824 29828 13852
rect 29816 13815 29828 13824
rect 29822 13812 29828 13815
rect 29880 13812 29886 13864
rect 31018 13812 31024 13864
rect 31076 13812 31082 13864
rect 24090 13747 24148 13753
rect 24228 13756 27108 13784
rect 28276 13756 28488 13784
rect 28997 13787 29055 13793
rect 22922 13716 22928 13728
rect 16500 13688 22928 13716
rect 22922 13676 22928 13688
rect 22980 13676 22986 13728
rect 23382 13676 23388 13728
rect 23440 13716 23446 13728
rect 24228 13716 24256 13756
rect 23440 13688 24256 13716
rect 23440 13676 23446 13688
rect 26970 13676 26976 13728
rect 27028 13676 27034 13728
rect 27080 13716 27108 13756
rect 28997 13753 29009 13787
rect 29043 13784 29055 13787
rect 29914 13784 29920 13796
rect 29043 13756 29920 13784
rect 29043 13753 29055 13756
rect 28997 13747 29055 13753
rect 29914 13744 29920 13756
rect 29972 13744 29978 13796
rect 28810 13716 28816 13728
rect 27080 13688 28816 13716
rect 28810 13676 28816 13688
rect 28868 13676 28874 13728
rect 31110 13676 31116 13728
rect 31168 13676 31174 13728
rect 552 13626 31648 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 12096 13626
rect 12148 13574 12160 13626
rect 12212 13574 12224 13626
rect 12276 13574 12288 13626
rect 12340 13574 12352 13626
rect 12404 13574 19870 13626
rect 19922 13574 19934 13626
rect 19986 13574 19998 13626
rect 20050 13574 20062 13626
rect 20114 13574 20126 13626
rect 20178 13574 27644 13626
rect 27696 13574 27708 13626
rect 27760 13574 27772 13626
rect 27824 13574 27836 13626
rect 27888 13574 27900 13626
rect 27952 13574 31648 13626
rect 552 13552 31648 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2832 13484 2881 13512
rect 2832 13472 2838 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 2869 13475 2927 13481
rect 3436 13484 3893 13512
rect 2685 13447 2743 13453
rect 2685 13413 2697 13447
rect 2731 13444 2743 13447
rect 3234 13444 3240 13456
rect 2731 13416 3240 13444
rect 2731 13413 2743 13416
rect 2685 13407 2743 13413
rect 3234 13404 3240 13416
rect 3292 13404 3298 13456
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 3436 13376 3464 13484
rect 3881 13481 3893 13484
rect 3927 13512 3939 13515
rect 4154 13512 4160 13524
rect 3927 13484 4160 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 7248 13484 12434 13512
rect 7248 13472 7254 13484
rect 3697 13447 3755 13453
rect 3697 13413 3709 13447
rect 3743 13444 3755 13447
rect 6264 13447 6322 13453
rect 3743 13416 4016 13444
rect 3743 13413 3755 13416
rect 3697 13407 3755 13413
rect 3988 13385 4016 13416
rect 6264 13413 6276 13447
rect 6310 13444 6322 13447
rect 6638 13444 6644 13456
rect 6310 13416 6644 13444
rect 6310 13413 6322 13416
rect 6264 13407 6322 13413
rect 6638 13404 6644 13416
rect 6696 13404 6702 13456
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 9493 13447 9551 13453
rect 6972 13416 9260 13444
rect 6972 13404 6978 13416
rect 2547 13348 3464 13376
rect 3513 13379 3571 13385
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 3513 13345 3525 13379
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 3789 13379 3847 13385
rect 3789 13345 3801 13379
rect 3835 13345 3847 13379
rect 3789 13339 3847 13345
rect 3973 13379 4031 13385
rect 3973 13345 3985 13379
rect 4019 13376 4031 13379
rect 5997 13379 6055 13385
rect 4019 13348 5948 13376
rect 4019 13345 4031 13348
rect 3973 13339 4031 13345
rect 3528 13308 3556 13339
rect 3804 13308 3832 13339
rect 5718 13308 5724 13320
rect 3528 13280 5724 13308
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 3421 13175 3479 13181
rect 3421 13141 3433 13175
rect 3467 13172 3479 13175
rect 3510 13172 3516 13184
rect 3467 13144 3516 13172
rect 3467 13141 3479 13144
rect 3421 13135 3479 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 5920 13172 5948 13348
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6086 13376 6092 13388
rect 6043 13348 6092 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7834 13376 7840 13388
rect 7156 13348 7840 13376
rect 7156 13336 7162 13348
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8067 13348 9137 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 8036 13308 8064 13339
rect 7524 13280 8064 13308
rect 7524 13268 7530 13280
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8573 13311 8631 13317
rect 8573 13308 8585 13311
rect 8260 13280 8585 13308
rect 8260 13268 8266 13280
rect 8573 13277 8585 13280
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9033 13311 9091 13317
rect 9033 13277 9045 13311
rect 9079 13308 9091 13311
rect 9232 13308 9260 13416
rect 9493 13413 9505 13447
rect 9539 13444 9551 13447
rect 9582 13444 9588 13456
rect 9539 13416 9588 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 9582 13404 9588 13416
rect 9640 13444 9646 13456
rect 12406 13444 12434 13484
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13081 13515 13139 13521
rect 13081 13512 13093 13515
rect 12952 13484 13093 13512
rect 12952 13472 12958 13484
rect 13081 13481 13093 13484
rect 13127 13481 13139 13515
rect 13081 13475 13139 13481
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13906 13512 13912 13524
rect 13320 13484 13912 13512
rect 13320 13472 13326 13484
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 14056 13484 14841 13512
rect 14056 13472 14062 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 14829 13475 14887 13481
rect 15028 13484 15485 13512
rect 15028 13453 15056 13484
rect 15473 13481 15485 13484
rect 15519 13512 15531 13515
rect 15562 13512 15568 13524
rect 15519 13484 15568 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 15746 13472 15752 13524
rect 15804 13472 15810 13524
rect 16850 13472 16856 13524
rect 16908 13472 16914 13524
rect 17034 13472 17040 13524
rect 17092 13472 17098 13524
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 20070 13512 20076 13524
rect 18932 13484 20076 13512
rect 18932 13472 18938 13484
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20530 13472 20536 13524
rect 20588 13512 20594 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 20588 13484 20637 13512
rect 20588 13472 20594 13484
rect 20625 13481 20637 13484
rect 20671 13481 20683 13515
rect 20625 13475 20683 13481
rect 21726 13472 21732 13524
rect 21784 13472 21790 13524
rect 21897 13515 21955 13521
rect 21897 13481 21909 13515
rect 21943 13512 21955 13515
rect 22186 13512 22192 13524
rect 21943 13484 22192 13512
rect 21943 13481 21955 13484
rect 21897 13475 21955 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22278 13472 22284 13524
rect 22336 13472 22342 13524
rect 23750 13472 23756 13524
rect 23808 13472 23814 13524
rect 24394 13472 24400 13524
rect 24452 13512 24458 13524
rect 24489 13515 24547 13521
rect 24489 13512 24501 13515
rect 24452 13484 24501 13512
rect 24452 13472 24458 13484
rect 24489 13481 24501 13484
rect 24535 13481 24547 13515
rect 24489 13475 24547 13481
rect 24854 13472 24860 13524
rect 24912 13472 24918 13524
rect 25130 13472 25136 13524
rect 25188 13472 25194 13524
rect 25314 13472 25320 13524
rect 25372 13512 25378 13524
rect 26053 13515 26111 13521
rect 26053 13512 26065 13515
rect 25372 13484 26065 13512
rect 25372 13472 25378 13484
rect 26053 13481 26065 13484
rect 26099 13481 26111 13515
rect 26053 13475 26111 13481
rect 26786 13472 26792 13524
rect 26844 13472 26850 13524
rect 28537 13515 28595 13521
rect 28537 13512 28549 13515
rect 27356 13484 28549 13512
rect 15013 13447 15071 13453
rect 15013 13444 15025 13447
rect 9640 13416 10088 13444
rect 12406 13416 15025 13444
rect 9640 13404 9646 13416
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13376 9919 13379
rect 9950 13376 9956 13388
rect 9907 13348 9956 13376
rect 9907 13345 9919 13348
rect 9861 13339 9919 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10060 13385 10088 13416
rect 15013 13413 15025 13416
rect 15059 13413 15071 13447
rect 15013 13407 15071 13413
rect 15194 13404 15200 13456
rect 15252 13404 15258 13456
rect 15930 13444 15936 13456
rect 15304 13416 15936 13444
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 10318 13336 10324 13388
rect 10376 13336 10382 13388
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10468 13348 11069 13376
rect 10468 13336 10474 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 13320 13348 13369 13376
rect 13320 13336 13326 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13376 13875 13379
rect 14642 13376 14648 13388
rect 13863 13348 14648 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 9766 13308 9772 13320
rect 9079 13280 9772 13308
rect 9079 13277 9091 13280
rect 9033 13271 9091 13277
rect 8956 13240 8984 13271
rect 9766 13268 9772 13280
rect 9824 13308 9830 13320
rect 11238 13308 11244 13320
rect 9824 13280 11244 13308
rect 9824 13268 9830 13280
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 13832 13308 13860 13339
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 15304 13385 15332 13416
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 17218 13444 17224 13456
rect 16224 13416 17224 13444
rect 16224 13385 16252 13416
rect 17218 13404 17224 13416
rect 17276 13404 17282 13456
rect 19168 13416 21956 13444
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 14976 13348 15301 13376
rect 14976 13336 14982 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13345 15899 13379
rect 15841 13339 15899 13345
rect 16209 13379 16267 13385
rect 16209 13345 16221 13379
rect 16255 13345 16267 13379
rect 16209 13339 16267 13345
rect 11940 13280 13124 13308
rect 11940 13268 11946 13280
rect 12986 13240 12992 13252
rect 6932 13212 7972 13240
rect 8956 13212 12992 13240
rect 6932 13172 6960 13212
rect 5920 13144 6960 13172
rect 7098 13132 7104 13184
rect 7156 13172 7162 13184
rect 7944 13181 7972 13212
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 7377 13175 7435 13181
rect 7377 13172 7389 13175
rect 7156 13144 7389 13172
rect 7156 13132 7162 13144
rect 7377 13141 7389 13144
rect 7423 13141 7435 13175
rect 7377 13135 7435 13141
rect 7929 13175 7987 13181
rect 7929 13141 7941 13175
rect 7975 13172 7987 13175
rect 9030 13172 9036 13184
rect 7975 13144 9036 13172
rect 7975 13141 7987 13144
rect 7929 13135 7987 13141
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13172 10011 13175
rect 10134 13172 10140 13184
rect 9999 13144 10140 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10505 13175 10563 13181
rect 10505 13172 10517 13175
rect 10284 13144 10517 13172
rect 10284 13132 10290 13144
rect 10505 13141 10517 13144
rect 10551 13141 10563 13175
rect 10505 13135 10563 13141
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 12802 13172 12808 13184
rect 11204 13144 12808 13172
rect 11204 13132 11210 13144
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13096 13172 13124 13280
rect 13280 13280 13860 13308
rect 13280 13172 13308 13280
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13964 13280 14105 13308
rect 13964 13268 13970 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14660 13308 14688 13336
rect 15856 13308 15884 13339
rect 16390 13336 16396 13388
rect 16448 13336 16454 13388
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 16577 13379 16635 13385
rect 16577 13345 16589 13379
rect 16623 13376 16635 13379
rect 16758 13376 16764 13388
rect 16623 13348 16764 13376
rect 16623 13345 16635 13348
rect 16577 13339 16635 13345
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 16960 13308 16988 13339
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 19168 13385 19196 13416
rect 21928 13388 21956 13416
rect 22094 13404 22100 13456
rect 22152 13404 22158 13456
rect 24578 13444 24584 13456
rect 24044 13416 24584 13444
rect 19153 13379 19211 13385
rect 19153 13376 19165 13379
rect 17920 13348 19165 13376
rect 17920 13336 17926 13348
rect 19153 13345 19165 13348
rect 19199 13345 19211 13379
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19153 13339 19211 13345
rect 19352 13348 19625 13376
rect 17034 13308 17040 13320
rect 14660 13280 17040 13308
rect 14093 13271 14151 13277
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 16022 13200 16028 13252
rect 16080 13240 16086 13252
rect 19352 13240 19380 13348
rect 19613 13345 19625 13348
rect 19659 13376 19671 13379
rect 19702 13376 19708 13388
rect 19659 13348 19708 13376
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 19702 13336 19708 13348
rect 19760 13336 19766 13388
rect 20070 13336 20076 13388
rect 20128 13336 20134 13388
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 20395 13348 20852 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 20165 13311 20223 13317
rect 20165 13308 20177 13311
rect 19843 13280 20177 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 20165 13277 20177 13280
rect 20211 13308 20223 13311
rect 20438 13308 20444 13320
rect 20211 13280 20444 13308
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 16080 13212 19380 13240
rect 19429 13243 19487 13249
rect 16080 13200 16086 13212
rect 19429 13209 19441 13243
rect 19475 13240 19487 13243
rect 19475 13212 19748 13240
rect 19475 13209 19487 13212
rect 19429 13203 19487 13209
rect 19720 13184 19748 13212
rect 20714 13200 20720 13252
rect 20772 13200 20778 13252
rect 20824 13240 20852 13348
rect 21634 13336 21640 13388
rect 21692 13336 21698 13388
rect 21910 13336 21916 13388
rect 21968 13336 21974 13388
rect 22373 13379 22431 13385
rect 22373 13376 22385 13379
rect 22020 13348 22385 13376
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 21048 13280 21097 13308
rect 21048 13268 21054 13280
rect 21085 13277 21097 13280
rect 21131 13308 21143 13311
rect 21131 13280 21496 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 21269 13243 21327 13249
rect 21269 13240 21281 13243
rect 20824 13212 21281 13240
rect 21269 13209 21281 13212
rect 21315 13209 21327 13243
rect 21468 13240 21496 13280
rect 21542 13268 21548 13320
rect 21600 13268 21606 13320
rect 21928 13308 21956 13336
rect 22020 13320 22048 13348
rect 22373 13345 22385 13348
rect 22419 13345 22431 13379
rect 22373 13339 22431 13345
rect 23934 13336 23940 13388
rect 23992 13336 23998 13388
rect 24044 13385 24072 13416
rect 24578 13404 24584 13416
rect 24636 13404 24642 13456
rect 24688 13416 24900 13444
rect 24029 13379 24087 13385
rect 24029 13345 24041 13379
rect 24075 13345 24087 13379
rect 24029 13339 24087 13345
rect 24210 13336 24216 13388
rect 24268 13336 24274 13388
rect 24688 13385 24716 13416
rect 24305 13379 24363 13385
rect 24305 13345 24317 13379
rect 24351 13345 24363 13379
rect 24305 13339 24363 13345
rect 24673 13379 24731 13385
rect 24673 13345 24685 13379
rect 24719 13345 24731 13379
rect 24673 13339 24731 13345
rect 24765 13379 24823 13385
rect 24765 13345 24777 13379
rect 24811 13345 24823 13379
rect 24872 13376 24900 13416
rect 25222 13404 25228 13456
rect 25280 13444 25286 13456
rect 25501 13447 25559 13453
rect 25501 13444 25513 13447
rect 25280 13416 25513 13444
rect 25280 13404 25286 13416
rect 25501 13413 25513 13416
rect 25547 13413 25559 13447
rect 25501 13407 25559 13413
rect 25593 13447 25651 13453
rect 25593 13413 25605 13447
rect 25639 13444 25651 13447
rect 26605 13447 26663 13453
rect 26605 13444 26617 13447
rect 25639 13416 26617 13444
rect 25639 13413 25651 13416
rect 25593 13407 25651 13413
rect 26605 13413 26617 13416
rect 26651 13444 26663 13447
rect 27356 13444 27384 13484
rect 28537 13481 28549 13484
rect 28583 13512 28595 13515
rect 28626 13512 28632 13524
rect 28583 13484 28632 13512
rect 28583 13481 28595 13484
rect 28537 13475 28595 13481
rect 28626 13472 28632 13484
rect 28684 13472 28690 13524
rect 28997 13515 29055 13521
rect 28997 13481 29009 13515
rect 29043 13512 29055 13515
rect 29546 13512 29552 13524
rect 29043 13484 29552 13512
rect 29043 13481 29055 13484
rect 28997 13475 29055 13481
rect 29546 13472 29552 13484
rect 29604 13472 29610 13524
rect 30834 13472 30840 13524
rect 30892 13512 30898 13524
rect 31297 13515 31355 13521
rect 31297 13512 31309 13515
rect 30892 13484 31309 13512
rect 30892 13472 30898 13484
rect 31297 13481 31309 13484
rect 31343 13481 31355 13515
rect 31297 13475 31355 13481
rect 26651 13416 27384 13444
rect 27424 13447 27482 13453
rect 26651 13413 26663 13416
rect 26605 13407 26663 13413
rect 27424 13413 27436 13447
rect 27470 13444 27482 13447
rect 27982 13444 27988 13456
rect 27470 13416 27988 13444
rect 27470 13413 27482 13416
rect 27424 13407 27482 13413
rect 27982 13404 27988 13416
rect 28040 13404 28046 13456
rect 29454 13404 29460 13456
rect 29512 13444 29518 13456
rect 30294 13447 30352 13453
rect 30294 13444 30306 13447
rect 29512 13416 30306 13444
rect 29512 13404 29518 13416
rect 30294 13413 30306 13416
rect 30340 13413 30352 13447
rect 30294 13407 30352 13413
rect 26050 13376 26056 13388
rect 24872 13348 26056 13376
rect 24765 13339 24823 13345
rect 22002 13308 22008 13320
rect 21928 13280 22008 13308
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 21726 13240 21732 13252
rect 21468 13212 21732 13240
rect 21269 13203 21327 13209
rect 21726 13200 21732 13212
rect 21784 13200 21790 13252
rect 24320 13240 24348 13339
rect 24394 13268 24400 13320
rect 24452 13308 24458 13320
rect 24780 13308 24808 13339
rect 26050 13336 26056 13348
rect 26108 13336 26114 13388
rect 26145 13379 26203 13385
rect 26145 13345 26157 13379
rect 26191 13376 26203 13379
rect 26326 13376 26332 13388
rect 26191 13348 26332 13376
rect 26191 13345 26203 13348
rect 26145 13339 26203 13345
rect 26326 13336 26332 13348
rect 26384 13336 26390 13388
rect 26421 13379 26479 13385
rect 26421 13345 26433 13379
rect 26467 13345 26479 13379
rect 26421 13339 26479 13345
rect 24452 13280 24808 13308
rect 24452 13268 24458 13280
rect 25682 13268 25688 13320
rect 25740 13268 25746 13320
rect 26436 13308 26464 13339
rect 26970 13336 26976 13388
rect 27028 13376 27034 13388
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 27028 13348 27169 13376
rect 27028 13336 27034 13348
rect 27157 13345 27169 13348
rect 27203 13345 27215 13379
rect 28166 13376 28172 13388
rect 27157 13339 27215 13345
rect 27264 13348 28172 13376
rect 27264 13308 27292 13348
rect 28166 13336 28172 13348
rect 28224 13336 28230 13388
rect 28902 13336 28908 13388
rect 28960 13336 28966 13388
rect 30561 13379 30619 13385
rect 30561 13345 30573 13379
rect 30607 13376 30619 13379
rect 31110 13376 31116 13388
rect 30607 13348 31116 13376
rect 30607 13345 30619 13348
rect 30561 13339 30619 13345
rect 31110 13336 31116 13348
rect 31168 13336 31174 13388
rect 26436 13280 27292 13308
rect 30745 13311 30803 13317
rect 30745 13277 30757 13311
rect 30791 13308 30803 13311
rect 30926 13308 30932 13320
rect 30791 13280 30932 13308
rect 30791 13277 30803 13280
rect 30745 13271 30803 13277
rect 30926 13268 30932 13280
rect 30984 13268 30990 13320
rect 24946 13240 24952 13252
rect 24320 13212 24952 13240
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 29181 13243 29239 13249
rect 29181 13209 29193 13243
rect 29227 13240 29239 13243
rect 29270 13240 29276 13252
rect 29227 13212 29276 13240
rect 29227 13209 29239 13212
rect 29181 13203 29239 13209
rect 29270 13200 29276 13212
rect 29328 13200 29334 13252
rect 13096 13144 13308 13172
rect 13538 13132 13544 13184
rect 13596 13172 13602 13184
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13596 13144 13737 13172
rect 13596 13132 13602 13144
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 13725 13135 13783 13141
rect 14734 13132 14740 13184
rect 14792 13132 14798 13184
rect 16666 13132 16672 13184
rect 16724 13172 16730 13184
rect 17678 13172 17684 13184
rect 16724 13144 17684 13172
rect 16724 13132 16730 13144
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19061 13175 19119 13181
rect 19061 13172 19073 13175
rect 18932 13144 19073 13172
rect 18932 13132 18938 13144
rect 19061 13141 19073 13144
rect 19107 13141 19119 13175
rect 19061 13135 19119 13141
rect 19702 13132 19708 13184
rect 19760 13132 19766 13184
rect 19794 13132 19800 13184
rect 19852 13132 19858 13184
rect 20990 13132 20996 13184
rect 21048 13172 21054 13184
rect 21450 13172 21456 13184
rect 21048 13144 21456 13172
rect 21048 13132 21054 13144
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 21913 13175 21971 13181
rect 21913 13141 21925 13175
rect 21959 13172 21971 13175
rect 22462 13172 22468 13184
rect 21959 13144 22468 13172
rect 21959 13141 21971 13144
rect 21913 13135 21971 13141
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 552 13082 31648 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 11436 13082
rect 11488 13030 11500 13082
rect 11552 13030 11564 13082
rect 11616 13030 11628 13082
rect 11680 13030 11692 13082
rect 11744 13030 19210 13082
rect 19262 13030 19274 13082
rect 19326 13030 19338 13082
rect 19390 13030 19402 13082
rect 19454 13030 19466 13082
rect 19518 13030 26984 13082
rect 27036 13030 27048 13082
rect 27100 13030 27112 13082
rect 27164 13030 27176 13082
rect 27228 13030 27240 13082
rect 27292 13030 31648 13082
rect 552 13008 31648 13030
rect 10229 12971 10287 12977
rect 10229 12937 10241 12971
rect 10275 12968 10287 12971
rect 10410 12968 10416 12980
rect 10275 12940 10416 12968
rect 10275 12937 10287 12940
rect 10229 12931 10287 12937
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 14550 12968 14556 12980
rect 13188 12940 14556 12968
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 9398 12900 9404 12912
rect 5132 12872 9404 12900
rect 5132 12860 5138 12872
rect 9398 12860 9404 12872
rect 9456 12900 9462 12912
rect 10594 12900 10600 12912
rect 9456 12872 10600 12900
rect 9456 12860 9462 12872
rect 10594 12860 10600 12872
rect 10652 12860 10658 12912
rect 5534 12792 5540 12844
rect 5592 12792 5598 12844
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5960 12804 6009 12832
rect 5960 12792 5966 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6086 12792 6092 12844
rect 6144 12792 6150 12844
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 7484 12804 8861 12832
rect 7484 12776 7512 12804
rect 8849 12801 8861 12804
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12832 8999 12835
rect 8987 12804 10640 12832
rect 8987 12801 8999 12804
rect 8941 12795 8999 12801
rect 2038 12724 2044 12776
rect 2096 12764 2102 12776
rect 2225 12767 2283 12773
rect 2225 12764 2237 12767
rect 2096 12736 2237 12764
rect 2096 12724 2102 12736
rect 2225 12733 2237 12736
rect 2271 12733 2283 12767
rect 2225 12727 2283 12733
rect 2593 12767 2651 12773
rect 2593 12733 2605 12767
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 1854 12656 1860 12708
rect 1912 12696 1918 12708
rect 2409 12699 2467 12705
rect 2409 12696 2421 12699
rect 1912 12668 2421 12696
rect 1912 12656 1918 12668
rect 2409 12665 2421 12668
rect 2455 12665 2467 12699
rect 2608 12696 2636 12727
rect 2774 12724 2780 12776
rect 2832 12724 2838 12776
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12764 7251 12767
rect 7466 12764 7472 12776
rect 7239 12736 7472 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 7742 12764 7748 12776
rect 7699 12736 7748 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 8202 12764 8208 12776
rect 7883 12736 8208 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 3510 12696 3516 12708
rect 2608 12668 3516 12696
rect 2409 12659 2467 12665
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 7098 12656 7104 12708
rect 7156 12696 7162 12708
rect 7852 12696 7880 12727
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8260 12736 8585 12764
rect 8260 12724 8266 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 9585 12767 9643 12773
rect 9585 12764 9597 12767
rect 9088 12736 9597 12764
rect 9088 12724 9094 12736
rect 9585 12733 9597 12736
rect 9631 12733 9643 12767
rect 9585 12727 9643 12733
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 9861 12767 9919 12773
rect 9861 12764 9873 12767
rect 9824 12736 9873 12764
rect 9824 12724 9830 12736
rect 9861 12733 9873 12736
rect 9907 12733 9919 12767
rect 10612 12764 10640 12804
rect 11514 12764 11520 12776
rect 10612 12736 11520 12764
rect 9861 12727 9919 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 11609 12767 11667 12773
rect 11609 12733 11621 12767
rect 11655 12764 11667 12767
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11655 12736 11805 12764
rect 11655 12733 11667 12736
rect 11609 12727 11667 12733
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 11882 12724 11888 12776
rect 11940 12764 11946 12776
rect 13188 12773 13216 12940
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 14918 12928 14924 12980
rect 14976 12928 14982 12980
rect 15470 12928 15476 12980
rect 15528 12968 15534 12980
rect 16482 12968 16488 12980
rect 15528 12940 16488 12968
rect 15528 12928 15534 12940
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 18877 12971 18935 12977
rect 18877 12937 18889 12971
rect 18923 12968 18935 12971
rect 19058 12968 19064 12980
rect 18923 12940 19064 12968
rect 18923 12937 18935 12940
rect 18877 12931 18935 12937
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19610 12928 19616 12980
rect 19668 12928 19674 12980
rect 21634 12928 21640 12980
rect 21692 12928 21698 12980
rect 28997 12971 29055 12977
rect 28997 12937 29009 12971
rect 29043 12968 29055 12971
rect 29178 12968 29184 12980
rect 29043 12940 29184 12968
rect 29043 12937 29055 12940
rect 28997 12931 29055 12937
rect 29178 12928 29184 12940
rect 29236 12928 29242 12980
rect 19153 12903 19211 12909
rect 19153 12869 19165 12903
rect 19199 12869 19211 12903
rect 19153 12863 19211 12869
rect 13538 12792 13544 12844
rect 13596 12792 13602 12844
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 19061 12835 19119 12841
rect 15436 12804 18460 12832
rect 15436 12792 15442 12804
rect 12713 12767 12771 12773
rect 12713 12764 12725 12767
rect 11940 12736 12725 12764
rect 11940 12724 11946 12736
rect 12713 12733 12725 12736
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 13172 12767 13230 12773
rect 13172 12733 13184 12767
rect 13218 12733 13230 12767
rect 13172 12727 13230 12733
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 14090 12764 14096 12776
rect 13311 12736 14096 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 16025 12767 16083 12773
rect 16025 12764 16037 12767
rect 15896 12736 16037 12764
rect 15896 12724 15902 12736
rect 16025 12733 16037 12736
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16390 12764 16396 12776
rect 16347 12736 16396 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16390 12724 16396 12736
rect 16448 12724 16454 12776
rect 16482 12724 16488 12776
rect 16540 12724 16546 12776
rect 16666 12724 16672 12776
rect 16724 12724 16730 12776
rect 17034 12724 17040 12776
rect 17092 12724 17098 12776
rect 7156 12668 7880 12696
rect 7156 12656 7162 12668
rect 11054 12656 11060 12708
rect 11112 12696 11118 12708
rect 11342 12699 11400 12705
rect 11342 12696 11354 12699
rect 11112 12668 11354 12696
rect 11112 12656 11118 12668
rect 11342 12665 11354 12668
rect 11388 12665 11400 12699
rect 11342 12659 11400 12665
rect 12986 12656 12992 12708
rect 13044 12696 13050 12708
rect 13814 12705 13820 12708
rect 13044 12668 13768 12696
rect 13044 12656 13050 12668
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 2004 12600 2145 12628
rect 2004 12588 2010 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 2133 12591 2191 12597
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 6914 12628 6920 12640
rect 5776 12600 6920 12628
rect 5776 12588 5782 12600
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7650 12588 7656 12640
rect 7708 12588 7714 12640
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10962 12628 10968 12640
rect 10091 12600 10968 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12492 12600 12633 12628
rect 12492 12588 12498 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13446 12628 13452 12640
rect 12943 12600 13452 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 13740 12628 13768 12668
rect 13808 12659 13820 12705
rect 13814 12656 13820 12659
rect 13872 12656 13878 12708
rect 16684 12696 16712 12724
rect 16316 12668 16712 12696
rect 16853 12699 16911 12705
rect 14642 12628 14648 12640
rect 13740 12600 14648 12628
rect 14642 12588 14648 12600
rect 14700 12628 14706 12640
rect 15378 12628 15384 12640
rect 14700 12600 15384 12628
rect 14700 12588 14706 12600
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 16316 12637 16344 12668
rect 16853 12665 16865 12699
rect 16899 12696 16911 12699
rect 18138 12696 18144 12708
rect 16899 12668 18144 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 18138 12656 18144 12668
rect 18196 12656 18202 12708
rect 18432 12696 18460 12804
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 19168 12832 19196 12863
rect 20070 12860 20076 12912
rect 20128 12900 20134 12912
rect 20165 12903 20223 12909
rect 20165 12900 20177 12903
rect 20128 12872 20177 12900
rect 20128 12860 20134 12872
rect 20165 12869 20177 12872
rect 20211 12869 20223 12903
rect 21652 12900 21680 12928
rect 20165 12863 20223 12869
rect 20824 12872 21680 12900
rect 19107 12804 19196 12832
rect 19429 12835 19487 12841
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 19429 12801 19441 12835
rect 19475 12832 19487 12835
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19475 12804 19809 12832
rect 19475 12801 19487 12804
rect 19429 12795 19487 12801
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12764 18843 12767
rect 19702 12764 19708 12776
rect 18831 12736 19708 12764
rect 18831 12733 18843 12736
rect 18785 12727 18843 12733
rect 19702 12724 19708 12736
rect 19760 12724 19766 12776
rect 19978 12724 19984 12776
rect 20036 12724 20042 12776
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 20257 12767 20315 12773
rect 20257 12733 20269 12767
rect 20303 12764 20315 12767
rect 20530 12764 20536 12776
rect 20303 12736 20536 12764
rect 20303 12733 20315 12736
rect 20257 12727 20315 12733
rect 19794 12696 19800 12708
rect 18432 12668 19800 12696
rect 19794 12656 19800 12668
rect 19852 12696 19858 12708
rect 20088 12696 20116 12727
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 20824 12773 20852 12872
rect 20898 12792 20904 12844
rect 20956 12832 20962 12844
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 20956 12804 21373 12832
rect 20956 12792 20962 12804
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 23750 12792 23756 12844
rect 23808 12832 23814 12844
rect 24394 12832 24400 12844
rect 23808 12804 24400 12832
rect 23808 12792 23814 12804
rect 24394 12792 24400 12804
rect 24452 12792 24458 12844
rect 28442 12792 28448 12844
rect 28500 12832 28506 12844
rect 30098 12832 30104 12844
rect 28500 12804 29316 12832
rect 28500 12792 28506 12804
rect 20809 12767 20867 12773
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 21140 12736 21465 12764
rect 21140 12724 21146 12736
rect 21453 12733 21465 12736
rect 21499 12733 21511 12767
rect 21453 12727 21511 12733
rect 21637 12767 21695 12773
rect 21637 12733 21649 12767
rect 21683 12764 21695 12767
rect 21726 12764 21732 12776
rect 21683 12736 21732 12764
rect 21683 12733 21695 12736
rect 21637 12727 21695 12733
rect 20622 12696 20628 12708
rect 19852 12668 20628 12696
rect 19852 12656 19858 12668
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 21468 12696 21496 12727
rect 21726 12724 21732 12736
rect 21784 12764 21790 12776
rect 23106 12764 23112 12776
rect 21784 12736 23112 12764
rect 21784 12724 21790 12736
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 28994 12724 29000 12776
rect 29052 12764 29058 12776
rect 29288 12773 29316 12804
rect 29472 12804 30104 12832
rect 29472 12773 29500 12804
rect 30098 12792 30104 12804
rect 30156 12792 30162 12844
rect 29181 12767 29239 12773
rect 29181 12764 29193 12767
rect 29052 12736 29193 12764
rect 29052 12724 29058 12736
rect 29181 12733 29193 12736
rect 29227 12733 29239 12767
rect 29181 12727 29239 12733
rect 29273 12767 29331 12773
rect 29273 12733 29285 12767
rect 29319 12733 29331 12767
rect 29273 12727 29331 12733
rect 29457 12767 29515 12773
rect 29457 12733 29469 12767
rect 29503 12733 29515 12767
rect 29457 12727 29515 12733
rect 29549 12767 29607 12773
rect 29549 12733 29561 12767
rect 29595 12733 29607 12767
rect 29549 12727 29607 12733
rect 21468 12668 21680 12696
rect 21652 12640 21680 12668
rect 28810 12656 28816 12708
rect 28868 12696 28874 12708
rect 29564 12696 29592 12727
rect 28868 12668 29592 12696
rect 28868 12656 28874 12668
rect 16301 12631 16359 12637
rect 16301 12597 16313 12631
rect 16347 12597 16359 12631
rect 16301 12591 16359 12597
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 17129 12631 17187 12637
rect 17129 12628 17141 12631
rect 16724 12600 17141 12628
rect 16724 12588 16730 12600
rect 17129 12597 17141 12600
rect 17175 12597 17187 12631
rect 17129 12591 17187 12597
rect 19058 12588 19064 12640
rect 19116 12588 19122 12640
rect 20714 12588 20720 12640
rect 20772 12588 20778 12640
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12628 21235 12631
rect 21358 12628 21364 12640
rect 21223 12600 21364 12628
rect 21223 12597 21235 12600
rect 21177 12591 21235 12597
rect 21358 12588 21364 12600
rect 21416 12588 21422 12640
rect 21634 12588 21640 12640
rect 21692 12588 21698 12640
rect 22002 12588 22008 12640
rect 22060 12628 22066 12640
rect 23750 12628 23756 12640
rect 22060 12600 23756 12628
rect 22060 12588 22066 12600
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 552 12538 31648 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 12096 12538
rect 12148 12486 12160 12538
rect 12212 12486 12224 12538
rect 12276 12486 12288 12538
rect 12340 12486 12352 12538
rect 12404 12486 19870 12538
rect 19922 12486 19934 12538
rect 19986 12486 19998 12538
rect 20050 12486 20062 12538
rect 20114 12486 20126 12538
rect 20178 12486 27644 12538
rect 27696 12486 27708 12538
rect 27760 12486 27772 12538
rect 27824 12486 27836 12538
rect 27888 12486 27900 12538
rect 27952 12486 31648 12538
rect 552 12464 31648 12486
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 1688 12396 3433 12424
rect 1688 12297 1716 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 5166 12424 5172 12436
rect 3421 12387 3479 12393
rect 3620 12396 5172 12424
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2194 12359 2252 12365
rect 2194 12356 2206 12359
rect 1903 12328 2206 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 2194 12325 2206 12328
rect 2240 12325 2252 12359
rect 2194 12319 2252 12325
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12257 1731 12291
rect 1673 12251 1731 12257
rect 1946 12248 1952 12300
rect 2004 12248 2010 12300
rect 2774 12288 2780 12300
rect 2056 12260 2780 12288
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 2056 12220 2084 12260
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3620 12297 3648 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7742 12424 7748 12436
rect 6972 12396 7748 12424
rect 6972 12384 6978 12396
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 9030 12424 9036 12436
rect 8798 12396 9036 12424
rect 3789 12359 3847 12365
rect 3789 12325 3801 12359
rect 3835 12356 3847 12359
rect 4062 12356 4068 12368
rect 3835 12328 4068 12356
rect 3835 12325 3847 12328
rect 3789 12319 3847 12325
rect 4062 12316 4068 12328
rect 4120 12316 4126 12368
rect 8798 12365 8826 12396
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9582 12384 9588 12436
rect 9640 12384 9646 12436
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 11054 12424 11060 12436
rect 10643 12396 11060 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 13722 12424 13728 12436
rect 12406 12396 13728 12424
rect 8783 12359 8841 12365
rect 8783 12325 8795 12359
rect 8829 12325 8841 12359
rect 9600 12356 9628 12384
rect 12406 12356 12434 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12393 13967 12427
rect 13909 12387 13967 12393
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 14734 12424 14740 12436
rect 14415 12396 14740 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 8783 12319 8841 12325
rect 8956 12328 9628 12356
rect 9968 12328 12434 12356
rect 12704 12359 12762 12365
rect 3605 12291 3663 12297
rect 3605 12288 3617 12291
rect 3476 12260 3617 12288
rect 3476 12248 3482 12260
rect 3605 12257 3617 12260
rect 3651 12257 3663 12291
rect 3605 12251 3663 12257
rect 3697 12291 3755 12297
rect 3697 12257 3709 12291
rect 3743 12257 3755 12291
rect 3697 12251 3755 12257
rect 3927 12291 3985 12297
rect 3927 12257 3939 12291
rect 3973 12288 3985 12291
rect 4430 12288 4436 12300
rect 3973 12260 4436 12288
rect 3973 12257 3985 12260
rect 3927 12251 3985 12257
rect 3712 12220 3740 12251
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 6914 12248 6920 12300
rect 6972 12248 6978 12300
rect 7098 12248 7104 12300
rect 7156 12248 7162 12300
rect 7466 12248 7472 12300
rect 7524 12248 7530 12300
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12257 8079 12291
rect 8021 12251 8079 12257
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 8251 12260 8309 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 1535 12192 2084 12220
rect 3344 12192 3740 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 3344 12161 3372 12192
rect 3329 12155 3387 12161
rect 3329 12121 3341 12155
rect 3375 12121 3387 12155
rect 3712 12152 3740 12192
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 4798 12220 4804 12232
rect 4111 12192 4804 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 6656 12192 7144 12220
rect 6656 12152 6684 12192
rect 7116 12164 7144 12192
rect 3712 12124 6684 12152
rect 3329 12115 3387 12121
rect 7006 12112 7012 12164
rect 7064 12112 7070 12164
rect 7098 12112 7104 12164
rect 7156 12112 7162 12164
rect 7374 12112 7380 12164
rect 7432 12152 7438 12164
rect 8036 12152 8064 12251
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 8481 12291 8539 12297
rect 8481 12288 8493 12291
rect 8444 12260 8493 12288
rect 8444 12248 8450 12260
rect 8481 12257 8493 12260
rect 8527 12257 8539 12291
rect 8481 12251 8539 12257
rect 8570 12248 8576 12300
rect 8628 12248 8634 12300
rect 8662 12248 8668 12300
rect 8720 12248 8726 12300
rect 8956 12297 8984 12328
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12257 8999 12291
rect 8941 12251 8999 12257
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9490 12288 9496 12300
rect 9263 12260 9496 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 9968 12297 9996 12328
rect 12704 12325 12716 12359
rect 12750 12356 12762 12359
rect 13924 12356 13952 12387
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 17957 12427 18015 12433
rect 17957 12393 17969 12427
rect 18003 12424 18015 12427
rect 18138 12424 18144 12436
rect 18003 12396 18144 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 19058 12384 19064 12436
rect 19116 12424 19122 12436
rect 19116 12396 19196 12424
rect 19116 12384 19122 12396
rect 12750 12328 13952 12356
rect 12750 12325 12762 12328
rect 12704 12319 12762 12325
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 17862 12356 17868 12368
rect 14240 12328 15056 12356
rect 14240 12316 14246 12328
rect 9585 12291 9643 12297
rect 9585 12257 9597 12291
rect 9631 12288 9643 12291
rect 9953 12291 10011 12297
rect 9631 12260 9904 12288
rect 9631 12257 9643 12260
rect 9585 12251 9643 12257
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8168 12192 9812 12220
rect 8168 12180 8174 12192
rect 9033 12155 9091 12161
rect 9033 12152 9045 12155
rect 7432 12124 9045 12152
rect 7432 12112 7438 12124
rect 9033 12121 9045 12124
rect 9079 12121 9091 12155
rect 9033 12115 9091 12121
rect 8113 12087 8171 12093
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8478 12084 8484 12096
rect 8159 12056 8484 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 9490 12084 9496 12096
rect 9447 12056 9496 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 9784 12084 9812 12192
rect 9876 12152 9904 12260
rect 9953 12257 9965 12291
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 10134 12248 10140 12300
rect 10192 12248 10198 12300
rect 10226 12248 10232 12300
rect 10284 12248 10290 12300
rect 10318 12248 10324 12300
rect 10376 12288 10382 12300
rect 11146 12288 11152 12300
rect 10376 12260 11152 12288
rect 10376 12248 10382 12260
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 11238 12248 11244 12300
rect 11296 12248 11302 12300
rect 11514 12248 11520 12300
rect 11572 12248 11578 12300
rect 12434 12248 12440 12300
rect 12492 12248 12498 12300
rect 14274 12248 14280 12300
rect 14332 12248 14338 12300
rect 15028 12297 15056 12328
rect 16408 12328 17868 12356
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 14384 12260 14749 12288
rect 11238 12152 11244 12164
rect 9876 12124 11244 12152
rect 11238 12112 11244 12124
rect 11296 12112 11302 12164
rect 11532 12152 11560 12248
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12220 11759 12223
rect 11882 12220 11888 12232
rect 11747 12192 11888 12220
rect 11747 12189 11759 12192
rect 11701 12183 11759 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 14384 12220 14412 12260
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 15013 12291 15071 12297
rect 15013 12257 15025 12291
rect 15059 12288 15071 12291
rect 15286 12288 15292 12300
rect 15059 12260 15292 12288
rect 15059 12257 15071 12260
rect 15013 12251 15071 12257
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 15470 12248 15476 12300
rect 15528 12248 15534 12300
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 13504 12192 14412 12220
rect 14553 12223 14611 12229
rect 13504 12180 13510 12192
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 12434 12152 12440 12164
rect 11532 12124 12440 12152
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 14568 12152 14596 12183
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14700 12192 14841 12220
rect 14700 12180 14706 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 15672 12220 15700 12251
rect 15746 12248 15752 12300
rect 15804 12248 15810 12300
rect 16408 12297 16436 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 19168 12365 19196 12396
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 21048 12396 23244 12424
rect 21048 12384 21054 12396
rect 19144 12359 19202 12365
rect 19144 12325 19156 12359
rect 19190 12325 19202 12359
rect 19144 12319 19202 12325
rect 19610 12316 19616 12368
rect 19668 12356 19674 12368
rect 19978 12356 19984 12368
rect 19668 12328 19984 12356
rect 19668 12316 19674 12328
rect 19978 12316 19984 12328
rect 20036 12356 20042 12368
rect 20533 12359 20591 12365
rect 20533 12356 20545 12359
rect 20036 12328 20545 12356
rect 20036 12316 20042 12328
rect 20533 12325 20545 12328
rect 20579 12325 20591 12359
rect 20533 12319 20591 12325
rect 21358 12316 21364 12368
rect 21416 12356 21422 12368
rect 21818 12356 21824 12368
rect 21416 12328 21824 12356
rect 21416 12316 21422 12328
rect 21818 12316 21824 12328
rect 21876 12316 21882 12368
rect 16393 12291 16451 12297
rect 16393 12257 16405 12291
rect 16439 12257 16451 12291
rect 16393 12251 16451 12257
rect 16577 12291 16635 12297
rect 16577 12257 16589 12291
rect 16623 12288 16635 12291
rect 16666 12288 16672 12300
rect 16623 12260 16672 12288
rect 16623 12257 16635 12260
rect 16577 12251 16635 12257
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 16850 12297 16856 12300
rect 16844 12251 16856 12297
rect 16850 12248 16856 12251
rect 16908 12248 16914 12300
rect 18690 12248 18696 12300
rect 18748 12248 18754 12300
rect 18874 12248 18880 12300
rect 18932 12248 18938 12300
rect 20162 12288 20168 12300
rect 18984 12260 20168 12288
rect 15672 12192 15884 12220
rect 14829 12183 14887 12189
rect 15856 12161 15884 12192
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18984 12220 19012 12260
rect 20162 12248 20168 12260
rect 20220 12288 20226 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 20220 12260 20361 12288
rect 20220 12248 20226 12260
rect 20349 12257 20361 12260
rect 20395 12257 20407 12291
rect 20349 12251 20407 12257
rect 20622 12248 20628 12300
rect 20680 12288 20686 12300
rect 22373 12291 22431 12297
rect 22373 12288 22385 12291
rect 20680 12260 22385 12288
rect 20680 12248 20686 12260
rect 22373 12257 22385 12260
rect 22419 12288 22431 12291
rect 22830 12288 22836 12300
rect 22419 12260 22836 12288
rect 22419 12257 22431 12260
rect 22373 12251 22431 12257
rect 22830 12248 22836 12260
rect 22888 12248 22894 12300
rect 23014 12248 23020 12300
rect 23072 12248 23078 12300
rect 23216 12297 23244 12396
rect 27338 12316 27344 12368
rect 27396 12356 27402 12368
rect 30285 12359 30343 12365
rect 30285 12356 30297 12359
rect 27396 12328 28948 12356
rect 27396 12316 27402 12328
rect 28920 12300 28948 12328
rect 29748 12328 30297 12356
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12257 23167 12291
rect 23109 12251 23167 12257
rect 23201 12291 23259 12297
rect 23201 12257 23213 12291
rect 23247 12257 23259 12291
rect 23201 12251 23259 12257
rect 23124 12220 23152 12251
rect 23750 12248 23756 12300
rect 23808 12288 23814 12300
rect 24121 12291 24179 12297
rect 24121 12288 24133 12291
rect 23808 12260 24133 12288
rect 23808 12248 23814 12260
rect 24121 12257 24133 12260
rect 24167 12257 24179 12291
rect 24121 12251 24179 12257
rect 28261 12291 28319 12297
rect 28261 12257 28273 12291
rect 28307 12288 28319 12291
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 28307 12260 28549 12288
rect 28307 12257 28319 12260
rect 28261 12251 28319 12257
rect 28537 12257 28549 12260
rect 28583 12257 28595 12291
rect 28537 12251 28595 12257
rect 28902 12248 28908 12300
rect 28960 12288 28966 12300
rect 29457 12291 29515 12297
rect 29457 12288 29469 12291
rect 28960 12260 29469 12288
rect 28960 12248 28966 12260
rect 29457 12257 29469 12260
rect 29503 12257 29515 12291
rect 29457 12251 29515 12257
rect 18012 12192 19012 12220
rect 21468 12192 23152 12220
rect 18012 12180 18018 12192
rect 21468 12164 21496 12192
rect 28810 12180 28816 12232
rect 28868 12220 28874 12232
rect 29089 12223 29147 12229
rect 29089 12220 29101 12223
rect 28868 12192 29101 12220
rect 28868 12180 28874 12192
rect 29089 12189 29101 12192
rect 29135 12189 29147 12223
rect 29472 12220 29500 12251
rect 29546 12248 29552 12300
rect 29604 12248 29610 12300
rect 29748 12297 29776 12328
rect 30285 12325 30297 12328
rect 30331 12325 30343 12359
rect 30285 12319 30343 12325
rect 29733 12291 29791 12297
rect 29733 12257 29745 12291
rect 29779 12257 29791 12291
rect 29733 12251 29791 12257
rect 29825 12291 29883 12297
rect 29825 12257 29837 12291
rect 29871 12288 29883 12291
rect 31018 12288 31024 12300
rect 29871 12260 31024 12288
rect 29871 12257 29883 12260
rect 29825 12251 29883 12257
rect 29840 12220 29868 12251
rect 31018 12248 31024 12260
rect 31076 12248 31082 12300
rect 29472 12192 29868 12220
rect 29089 12183 29147 12189
rect 30926 12180 30932 12232
rect 30984 12180 30990 12232
rect 15197 12155 15255 12161
rect 15197 12152 15209 12155
rect 14568 12124 15209 12152
rect 15197 12121 15209 12124
rect 15243 12121 15255 12155
rect 15197 12115 15255 12121
rect 15841 12155 15899 12161
rect 15841 12121 15853 12155
rect 15887 12152 15899 12155
rect 16482 12152 16488 12164
rect 15887 12124 16488 12152
rect 15887 12121 15899 12124
rect 15841 12115 15899 12121
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 20717 12155 20775 12161
rect 20717 12121 20729 12155
rect 20763 12152 20775 12155
rect 21450 12152 21456 12164
rect 20763 12124 21456 12152
rect 20763 12121 20775 12124
rect 20717 12115 20775 12121
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 26418 12152 26424 12164
rect 21560 12124 26424 12152
rect 10318 12084 10324 12096
rect 9784 12056 10324 12084
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 10652 12056 13829 12084
rect 10652 12044 10658 12056
rect 13817 12053 13829 12056
rect 13863 12084 13875 12087
rect 13906 12084 13912 12096
rect 13863 12056 13912 12084
rect 13863 12053 13875 12056
rect 13817 12047 13875 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 14056 12056 14749 12084
rect 14056 12044 14062 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 14737 12047 14795 12053
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12084 15623 12087
rect 15746 12084 15752 12096
rect 15611 12056 15752 12084
rect 15611 12053 15623 12056
rect 15565 12047 15623 12053
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 16172 12056 16313 12084
rect 16172 12044 16178 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16301 12047 16359 12053
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 18506 12084 18512 12096
rect 16448 12056 18512 12084
rect 16448 12044 16454 12056
rect 18506 12044 18512 12056
rect 18564 12084 18570 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18564 12056 18613 12084
rect 18564 12044 18570 12056
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 18601 12047 18659 12053
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 20257 12087 20315 12093
rect 20257 12084 20269 12087
rect 18748 12056 20269 12084
rect 18748 12044 18754 12056
rect 20257 12053 20269 12056
rect 20303 12053 20315 12087
rect 20257 12047 20315 12053
rect 20346 12044 20352 12096
rect 20404 12084 20410 12096
rect 21560 12084 21588 12124
rect 26418 12112 26424 12124
rect 26476 12112 26482 12164
rect 20404 12056 21588 12084
rect 20404 12044 20410 12056
rect 21726 12044 21732 12096
rect 21784 12084 21790 12096
rect 21910 12084 21916 12096
rect 21784 12056 21916 12084
rect 21784 12044 21790 12056
rect 21910 12044 21916 12056
rect 21968 12084 21974 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 21968 12056 22293 12084
rect 21968 12044 21974 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22281 12047 22339 12053
rect 23474 12044 23480 12096
rect 23532 12044 23538 12096
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 23661 12087 23719 12093
rect 23661 12084 23673 12087
rect 23624 12056 23673 12084
rect 23624 12044 23630 12056
rect 23661 12053 23673 12056
rect 23707 12053 23719 12087
rect 23661 12047 23719 12053
rect 23842 12044 23848 12096
rect 23900 12084 23906 12096
rect 24029 12087 24087 12093
rect 24029 12084 24041 12087
rect 23900 12056 24041 12084
rect 23900 12044 23906 12056
rect 24029 12053 24041 12056
rect 24075 12053 24087 12087
rect 24029 12047 24087 12053
rect 28166 12044 28172 12096
rect 28224 12044 28230 12096
rect 29178 12044 29184 12096
rect 29236 12084 29242 12096
rect 29365 12087 29423 12093
rect 29365 12084 29377 12087
rect 29236 12056 29377 12084
rect 29236 12044 29242 12056
rect 29365 12053 29377 12056
rect 29411 12053 29423 12087
rect 29365 12047 29423 12053
rect 29730 12044 29736 12096
rect 29788 12044 29794 12096
rect 29914 12044 29920 12096
rect 29972 12044 29978 12096
rect 552 11994 31648 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 11436 11994
rect 11488 11942 11500 11994
rect 11552 11942 11564 11994
rect 11616 11942 11628 11994
rect 11680 11942 11692 11994
rect 11744 11942 19210 11994
rect 19262 11942 19274 11994
rect 19326 11942 19338 11994
rect 19390 11942 19402 11994
rect 19454 11942 19466 11994
rect 19518 11942 26984 11994
rect 27036 11942 27048 11994
rect 27100 11942 27112 11994
rect 27164 11942 27176 11994
rect 27228 11942 27240 11994
rect 27292 11942 31648 11994
rect 552 11920 31648 11942
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3568 11852 3985 11880
rect 3568 11840 3574 11852
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 3973 11843 4031 11849
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 7800 11852 9352 11880
rect 7800 11840 7806 11852
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 9324 11812 9352 11852
rect 10042 11840 10048 11892
rect 10100 11840 10106 11892
rect 10152 11852 11468 11880
rect 10152 11812 10180 11852
rect 3476 11784 4016 11812
rect 9324 11784 10180 11812
rect 11440 11812 11468 11852
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12492 11852 13768 11880
rect 12492 11840 12498 11852
rect 13630 11812 13636 11824
rect 11440 11784 13636 11812
rect 3476 11772 3482 11784
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1535 11716 1685 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 3878 11744 3884 11756
rect 1673 11707 1731 11713
rect 3344 11716 3884 11744
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 1627 11648 2084 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 2056 11620 2084 11648
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 3344 11676 3372 11716
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 3988 11744 4016 11784
rect 13630 11772 13636 11784
rect 13688 11772 13694 11824
rect 13740 11812 13768 11852
rect 13814 11840 13820 11892
rect 13872 11840 13878 11892
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 15654 11880 15660 11892
rect 14332 11852 15660 11880
rect 14332 11840 14338 11852
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 16850 11880 16856 11892
rect 16255 11852 16856 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 18046 11840 18052 11892
rect 18104 11880 18110 11892
rect 28074 11880 28080 11892
rect 18104 11852 28080 11880
rect 18104 11840 18110 11852
rect 28074 11840 28080 11852
rect 28132 11840 28138 11892
rect 28810 11840 28816 11892
rect 28868 11840 28874 11892
rect 17954 11812 17960 11824
rect 13740 11784 17960 11812
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 21726 11812 21732 11824
rect 18340 11784 21732 11812
rect 3988 11716 4108 11744
rect 2556 11648 3372 11676
rect 2556 11636 2562 11648
rect 3418 11636 3424 11688
rect 3476 11636 3482 11688
rect 3786 11685 3792 11688
rect 3743 11679 3792 11685
rect 3743 11645 3755 11679
rect 3789 11645 3792 11679
rect 3743 11639 3792 11645
rect 3786 11636 3792 11639
rect 3844 11636 3850 11688
rect 3970 11636 3976 11688
rect 4028 11636 4034 11688
rect 4080 11654 4108 11716
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 4212 11716 4292 11744
rect 4212 11704 4218 11716
rect 4264 11676 4292 11716
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4396 11716 4629 11744
rect 4396 11704 4402 11716
rect 4617 11713 4629 11716
rect 4663 11744 4675 11747
rect 4890 11744 4896 11756
rect 4663 11716 4896 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6328 11716 6837 11744
rect 6328 11704 6334 11716
rect 6825 11713 6837 11716
rect 6871 11744 6883 11747
rect 7374 11744 7380 11756
rect 6871 11716 7380 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 15194 11744 15200 11756
rect 13740 11716 15200 11744
rect 4158 11657 4216 11663
rect 4158 11654 4170 11657
rect 1946 11617 1952 11620
rect 1940 11571 1952 11617
rect 1946 11568 1952 11571
rect 2004 11568 2010 11620
rect 2038 11568 2044 11620
rect 2096 11568 2102 11620
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 3237 11611 3295 11617
rect 3237 11608 3249 11611
rect 2832 11580 3249 11608
rect 2832 11568 2838 11580
rect 3237 11577 3249 11580
rect 3283 11577 3295 11611
rect 3237 11571 3295 11577
rect 3510 11568 3516 11620
rect 3568 11568 3574 11620
rect 3602 11568 3608 11620
rect 3660 11608 3666 11620
rect 3988 11608 4016 11636
rect 4080 11626 4170 11654
rect 4158 11623 4170 11626
rect 4204 11623 4216 11657
rect 4264 11648 4384 11676
rect 4158 11617 4216 11623
rect 4356 11617 4384 11648
rect 4430 11636 4436 11688
rect 4488 11685 4494 11688
rect 4488 11679 4537 11685
rect 4488 11645 4491 11679
rect 4525 11645 4537 11679
rect 4488 11639 4537 11645
rect 4488 11636 4522 11639
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 6089 11679 6147 11685
rect 6089 11676 6101 11679
rect 5592 11648 6101 11676
rect 5592 11636 5598 11648
rect 6089 11645 6101 11648
rect 6135 11645 6147 11679
rect 6089 11639 6147 11645
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7190 11676 7196 11688
rect 7055 11648 7196 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7466 11636 7472 11688
rect 7524 11636 7530 11688
rect 7650 11636 7656 11688
rect 7708 11676 7714 11688
rect 7708 11648 7788 11676
rect 7708 11636 7714 11648
rect 3660 11580 4016 11608
rect 4249 11611 4307 11617
rect 3660 11568 3666 11580
rect 4249 11577 4261 11611
rect 4295 11577 4307 11611
rect 4249 11571 4307 11577
rect 4341 11611 4399 11617
rect 4341 11577 4353 11611
rect 4387 11577 4399 11611
rect 4494 11608 4522 11636
rect 5718 11608 5724 11620
rect 4494 11580 5724 11608
rect 4341 11571 4399 11577
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 4264 11540 4292 11571
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 7760 11608 7788 11648
rect 8018 11636 8024 11688
rect 8076 11636 8082 11688
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8159 11648 8401 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8645 11679 8703 11685
rect 8645 11676 8657 11679
rect 8536 11648 8657 11676
rect 8536 11636 8542 11648
rect 8645 11645 8657 11648
rect 8691 11645 8703 11679
rect 8645 11639 8703 11645
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10778 11676 10784 11688
rect 10008 11648 10784 11676
rect 10008 11636 10014 11648
rect 10778 11636 10784 11648
rect 10836 11676 10842 11688
rect 11425 11679 11483 11685
rect 10836 11648 11284 11676
rect 10836 11636 10842 11648
rect 9030 11608 9036 11620
rect 7760 11580 9036 11608
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 11158 11611 11216 11617
rect 11158 11608 11170 11611
rect 10376 11580 11170 11608
rect 10376 11568 10382 11580
rect 11158 11577 11170 11580
rect 11204 11577 11216 11611
rect 11256 11608 11284 11648
rect 11425 11645 11437 11679
rect 11471 11676 11483 11679
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 11471 11648 11621 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11676 11759 11679
rect 11790 11676 11796 11688
rect 11747 11648 11796 11676
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 12986 11636 12992 11688
rect 13044 11636 13050 11688
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 13740 11685 13768 11716
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 15528 11716 18184 11744
rect 15528 11704 15534 11716
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 14090 11636 14096 11688
rect 14148 11636 14154 11688
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 15289 11611 15347 11617
rect 15289 11608 15301 11611
rect 11256 11580 15301 11608
rect 11158 11571 11216 11577
rect 15289 11577 15301 11580
rect 15335 11577 15347 11611
rect 15289 11571 15347 11577
rect 4890 11540 4896 11552
rect 3099 11512 4896 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5868 11512 6009 11540
rect 5868 11500 5874 11512
rect 5997 11509 6009 11512
rect 6043 11509 6055 11543
rect 5997 11503 6055 11509
rect 7193 11543 7251 11549
rect 7193 11509 7205 11543
rect 7239 11540 7251 11543
rect 7558 11540 7564 11552
rect 7239 11512 7564 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 7653 11543 7711 11549
rect 7653 11509 7665 11543
rect 7699 11540 7711 11543
rect 8386 11540 8392 11552
rect 7699 11512 8392 11540
rect 7699 11509 7711 11512
rect 7653 11503 7711 11509
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9364 11512 9781 11540
rect 9364 11500 9370 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 13081 11543 13139 11549
rect 13081 11509 13093 11543
rect 13127 11540 13139 11543
rect 13998 11540 14004 11552
rect 13127 11512 14004 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 15378 11500 15384 11552
rect 15436 11500 15442 11552
rect 15580 11540 15608 11639
rect 15746 11636 15752 11688
rect 15804 11636 15810 11688
rect 15856 11685 15884 11716
rect 15841 11679 15899 11685
rect 15841 11645 15853 11679
rect 15887 11645 15899 11679
rect 15841 11639 15899 11645
rect 15930 11636 15936 11688
rect 15988 11636 15994 11688
rect 16485 11679 16543 11685
rect 16485 11645 16497 11679
rect 16531 11676 16543 11679
rect 16574 11676 16580 11688
rect 16531 11648 16580 11676
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 18156 11685 18184 11716
rect 18340 11685 18368 11784
rect 18598 11704 18604 11756
rect 18656 11744 18662 11756
rect 19242 11744 19248 11756
rect 18656 11716 19248 11744
rect 18656 11704 18662 11716
rect 19242 11704 19248 11716
rect 19300 11744 19306 11756
rect 19337 11747 19395 11753
rect 19337 11744 19349 11747
rect 19300 11716 19349 11744
rect 19300 11704 19306 11716
rect 19337 11713 19349 11716
rect 19383 11713 19395 11747
rect 20622 11744 20628 11756
rect 19337 11707 19395 11713
rect 19536 11716 20628 11744
rect 18141 11679 18199 11685
rect 18141 11645 18153 11679
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11645 18383 11679
rect 18325 11639 18383 11645
rect 17678 11568 17684 11620
rect 17736 11608 17742 11620
rect 18233 11611 18291 11617
rect 18233 11608 18245 11611
rect 17736 11580 18245 11608
rect 17736 11568 17742 11580
rect 18233 11577 18245 11580
rect 18279 11577 18291 11611
rect 18233 11571 18291 11577
rect 18340 11540 18368 11639
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 19536 11685 19564 11716
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18564 11648 18981 11676
rect 18564 11636 18570 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19521 11679 19579 11685
rect 19521 11645 19533 11679
rect 19567 11645 19579 11679
rect 19705 11679 19763 11685
rect 19705 11676 19717 11679
rect 19521 11639 19579 11645
rect 19628 11648 19717 11676
rect 19628 11608 19656 11648
rect 19705 11645 19717 11648
rect 19751 11645 19763 11679
rect 19705 11639 19763 11645
rect 19794 11636 19800 11688
rect 19852 11676 19858 11688
rect 19889 11679 19947 11685
rect 19889 11676 19901 11679
rect 19852 11648 19901 11676
rect 19852 11636 19858 11648
rect 19889 11645 19901 11648
rect 19935 11645 19947 11679
rect 19889 11639 19947 11645
rect 19978 11636 19984 11688
rect 20036 11636 20042 11688
rect 20162 11636 20168 11688
rect 20220 11636 20226 11688
rect 21008 11685 21036 11784
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 23014 11772 23020 11824
rect 23072 11812 23078 11824
rect 23293 11815 23351 11821
rect 23293 11812 23305 11815
rect 23072 11784 23305 11812
rect 23072 11772 23078 11784
rect 23293 11781 23305 11784
rect 23339 11781 23351 11815
rect 23293 11775 23351 11781
rect 23474 11772 23480 11824
rect 23532 11812 23538 11824
rect 23532 11784 23796 11812
rect 23532 11772 23538 11784
rect 21450 11744 21456 11756
rect 21284 11716 21456 11744
rect 20993 11679 21051 11685
rect 20993 11645 21005 11679
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 21174 11636 21180 11688
rect 21232 11636 21238 11688
rect 21284 11685 21312 11716
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 21269 11679 21327 11685
rect 21269 11645 21281 11679
rect 21315 11645 21327 11679
rect 21269 11639 21327 11645
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 21542 11676 21548 11688
rect 21416 11648 21548 11676
rect 21416 11636 21422 11648
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 21726 11636 21732 11688
rect 21784 11636 21790 11688
rect 23768 11676 23796 11784
rect 26418 11772 26424 11824
rect 26476 11772 26482 11824
rect 26605 11815 26663 11821
rect 26605 11781 26617 11815
rect 26651 11812 26663 11815
rect 26651 11784 27476 11812
rect 26651 11781 26663 11784
rect 26605 11775 26663 11781
rect 23842 11704 23848 11756
rect 23900 11704 23906 11756
rect 26620 11744 26648 11775
rect 27338 11744 27344 11756
rect 26436 11716 26648 11744
rect 27172 11716 27344 11744
rect 24101 11679 24159 11685
rect 24101 11676 24113 11679
rect 23768 11648 24113 11676
rect 24101 11645 24113 11648
rect 24147 11645 24159 11679
rect 25314 11676 25320 11688
rect 24101 11639 24159 11645
rect 24412 11648 25320 11676
rect 19168 11580 19656 11608
rect 15580 11512 18368 11540
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 19168 11549 19196 11580
rect 20714 11568 20720 11620
rect 20772 11608 20778 11620
rect 21376 11608 21404 11636
rect 20772 11580 21404 11608
rect 21637 11611 21695 11617
rect 20772 11568 20778 11580
rect 21637 11577 21649 11611
rect 21683 11608 21695 11611
rect 21974 11611 22032 11617
rect 21974 11608 21986 11611
rect 21683 11580 21986 11608
rect 21683 11577 21695 11580
rect 21637 11571 21695 11577
rect 21974 11577 21986 11580
rect 22020 11577 22032 11611
rect 21974 11571 22032 11577
rect 23474 11568 23480 11620
rect 23532 11568 23538 11620
rect 23661 11611 23719 11617
rect 23661 11577 23673 11611
rect 23707 11608 23719 11611
rect 24210 11608 24216 11620
rect 23707 11580 24216 11608
rect 23707 11577 23719 11580
rect 23661 11571 23719 11577
rect 24210 11568 24216 11580
rect 24268 11568 24274 11620
rect 19153 11543 19211 11549
rect 19153 11540 19165 11543
rect 18472 11512 19165 11540
rect 18472 11500 18478 11512
rect 19153 11509 19165 11512
rect 19199 11509 19211 11543
rect 19153 11503 19211 11509
rect 19242 11500 19248 11552
rect 19300 11540 19306 11552
rect 19702 11540 19708 11552
rect 19300 11512 19708 11540
rect 19300 11500 19306 11512
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 19886 11540 19892 11552
rect 19852 11512 19892 11540
rect 19852 11500 19858 11512
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 20073 11543 20131 11549
rect 20073 11509 20085 11543
rect 20119 11540 20131 11543
rect 21266 11540 21272 11552
rect 20119 11512 21272 11540
rect 20119 11509 20131 11512
rect 20073 11503 20131 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 23109 11543 23167 11549
rect 23109 11509 23121 11543
rect 23155 11540 23167 11543
rect 23290 11540 23296 11552
rect 23155 11512 23296 11540
rect 23155 11509 23167 11512
rect 23109 11503 23167 11509
rect 23290 11500 23296 11512
rect 23348 11540 23354 11552
rect 24412 11540 24440 11648
rect 25314 11636 25320 11648
rect 25372 11636 25378 11688
rect 25471 11679 25529 11685
rect 25471 11645 25483 11679
rect 25517 11676 25529 11679
rect 25590 11676 25596 11688
rect 25517 11648 25596 11676
rect 25517 11645 25529 11648
rect 25471 11639 25529 11645
rect 25590 11636 25596 11648
rect 25648 11636 25654 11688
rect 25774 11636 25780 11688
rect 25832 11636 25838 11688
rect 25866 11636 25872 11688
rect 25924 11636 25930 11688
rect 26283 11679 26341 11685
rect 26283 11645 26295 11679
rect 26329 11676 26341 11679
rect 26436 11676 26464 11716
rect 26329 11648 26464 11676
rect 26513 11679 26571 11685
rect 26329 11645 26341 11648
rect 26283 11639 26341 11645
rect 26513 11645 26525 11679
rect 26559 11645 26571 11679
rect 26513 11639 26571 11645
rect 25685 11611 25743 11617
rect 25685 11577 25697 11611
rect 25731 11608 25743 11611
rect 26053 11611 26111 11617
rect 26053 11608 26065 11611
rect 25731 11580 26065 11608
rect 25731 11577 25743 11580
rect 25685 11571 25743 11577
rect 26053 11577 26065 11580
rect 26099 11577 26111 11611
rect 26053 11571 26111 11577
rect 26145 11611 26203 11617
rect 26145 11577 26157 11611
rect 26191 11608 26203 11611
rect 26528 11608 26556 11639
rect 26786 11636 26792 11688
rect 26844 11636 26850 11688
rect 26878 11636 26884 11688
rect 26936 11636 26942 11688
rect 27172 11685 27200 11716
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 27448 11744 27476 11784
rect 27448 11716 27568 11744
rect 27157 11679 27215 11685
rect 27157 11645 27169 11679
rect 27203 11645 27215 11679
rect 27157 11639 27215 11645
rect 27249 11679 27307 11685
rect 27249 11645 27261 11679
rect 27295 11676 27307 11679
rect 27433 11679 27491 11685
rect 27433 11676 27445 11679
rect 27295 11648 27445 11676
rect 27295 11645 27307 11648
rect 27249 11639 27307 11645
rect 27433 11645 27445 11648
rect 27479 11645 27491 11679
rect 27540 11676 27568 11716
rect 29178 11704 29184 11756
rect 29236 11704 29242 11756
rect 28166 11676 28172 11688
rect 27540 11648 28172 11676
rect 27433 11639 27491 11645
rect 28166 11636 28172 11648
rect 28224 11636 28230 11688
rect 29448 11679 29506 11685
rect 29448 11645 29460 11679
rect 29494 11676 29506 11679
rect 29730 11676 29736 11688
rect 29494 11648 29736 11676
rect 29494 11645 29506 11648
rect 29448 11639 29506 11645
rect 29730 11636 29736 11648
rect 29788 11636 29794 11688
rect 31110 11636 31116 11688
rect 31168 11676 31174 11688
rect 31205 11679 31263 11685
rect 31205 11676 31217 11679
rect 31168 11648 31217 11676
rect 31168 11636 31174 11648
rect 31205 11645 31217 11648
rect 31251 11645 31263 11679
rect 31205 11639 31263 11645
rect 26191 11580 26556 11608
rect 26191 11577 26203 11580
rect 26145 11571 26203 11577
rect 23348 11512 24440 11540
rect 23348 11500 23354 11512
rect 25222 11500 25228 11552
rect 25280 11540 25286 11552
rect 26160 11540 26188 11571
rect 27062 11568 27068 11620
rect 27120 11568 27126 11620
rect 27522 11568 27528 11620
rect 27580 11608 27586 11620
rect 27678 11611 27736 11617
rect 27678 11608 27690 11611
rect 27580 11580 27690 11608
rect 27580 11568 27586 11580
rect 27678 11577 27690 11580
rect 27724 11577 27736 11611
rect 27678 11571 27736 11577
rect 29086 11568 29092 11620
rect 29144 11608 29150 11620
rect 30653 11611 30711 11617
rect 30653 11608 30665 11611
rect 29144 11580 30665 11608
rect 29144 11568 29150 11580
rect 30653 11577 30665 11580
rect 30699 11577 30711 11611
rect 30653 11571 30711 11577
rect 25280 11512 26188 11540
rect 25280 11500 25286 11512
rect 28534 11500 28540 11552
rect 28592 11540 28598 11552
rect 30561 11543 30619 11549
rect 30561 11540 30573 11543
rect 28592 11512 30573 11540
rect 28592 11500 28598 11512
rect 30561 11509 30573 11512
rect 30607 11540 30619 11543
rect 30742 11540 30748 11552
rect 30607 11512 30748 11540
rect 30607 11509 30619 11512
rect 30561 11503 30619 11509
rect 30742 11500 30748 11512
rect 30800 11500 30806 11552
rect 552 11450 31648 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 12096 11450
rect 12148 11398 12160 11450
rect 12212 11398 12224 11450
rect 12276 11398 12288 11450
rect 12340 11398 12352 11450
rect 12404 11398 19870 11450
rect 19922 11398 19934 11450
rect 19986 11398 19998 11450
rect 20050 11398 20062 11450
rect 20114 11398 20126 11450
rect 20178 11398 27644 11450
rect 27696 11398 27708 11450
rect 27760 11398 27772 11450
rect 27824 11398 27836 11450
rect 27888 11398 27900 11450
rect 27952 11398 31648 11450
rect 552 11376 31648 11398
rect 3510 11296 3516 11348
rect 3568 11336 3574 11348
rect 3697 11339 3755 11345
rect 3697 11336 3709 11339
rect 3568 11308 3709 11336
rect 3568 11296 3574 11308
rect 3697 11305 3709 11308
rect 3743 11305 3755 11339
rect 3697 11299 3755 11305
rect 2038 11160 2044 11212
rect 2096 11160 2102 11212
rect 2590 11209 2596 11212
rect 2584 11163 2596 11209
rect 2590 11160 2596 11163
rect 2648 11160 2654 11212
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2179 11104 2329 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 3712 11064 3740 11299
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 6546 11336 6552 11348
rect 5224 11308 6552 11336
rect 5224 11296 5230 11308
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 5184 11209 5212 11296
rect 5261 11271 5319 11277
rect 5261 11237 5273 11271
rect 5307 11268 5319 11271
rect 5902 11268 5908 11280
rect 5307 11240 5908 11268
rect 5307 11237 5319 11240
rect 5261 11231 5319 11237
rect 5902 11228 5908 11240
rect 5960 11228 5966 11280
rect 6086 11277 6092 11280
rect 6080 11231 6092 11277
rect 6086 11228 6092 11231
rect 6144 11228 6150 11280
rect 6178 11228 6184 11280
rect 6236 11268 6242 11280
rect 7208 11268 7236 11299
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 7616 11308 8524 11336
rect 7616 11296 7622 11308
rect 7650 11268 7656 11280
rect 6236 11240 7656 11268
rect 6236 11228 6242 11240
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 8496 11268 8524 11308
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 8628 11308 9229 11336
rect 8628 11296 8634 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 10163 11339 10221 11345
rect 10163 11305 10175 11339
rect 10209 11336 10221 11339
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10209 11308 10977 11336
rect 10209 11305 10221 11308
rect 10163 11299 10221 11305
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 19610 11336 19616 11348
rect 13688 11308 19616 11336
rect 13688 11296 13694 11308
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 19794 11296 19800 11348
rect 19852 11336 19858 11348
rect 20530 11336 20536 11348
rect 19852 11308 20536 11336
rect 19852 11296 19858 11308
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 21726 11296 21732 11348
rect 21784 11336 21790 11348
rect 21913 11339 21971 11345
rect 21913 11336 21925 11339
rect 21784 11308 21925 11336
rect 21784 11296 21790 11308
rect 21913 11305 21925 11308
rect 21959 11305 21971 11339
rect 21913 11299 21971 11305
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 25222 11336 25228 11348
rect 23532 11308 25228 11336
rect 23532 11296 23538 11308
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 25774 11336 25780 11348
rect 25547 11308 25780 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 25774 11296 25780 11308
rect 25832 11296 25838 11348
rect 26786 11296 26792 11348
rect 26844 11336 26850 11348
rect 28353 11339 28411 11345
rect 28353 11336 28365 11339
rect 26844 11308 28365 11336
rect 26844 11296 26850 11308
rect 28353 11305 28365 11308
rect 28399 11305 28411 11339
rect 28353 11299 28411 11305
rect 28810 11296 28816 11348
rect 28868 11296 28874 11348
rect 29181 11339 29239 11345
rect 29181 11305 29193 11339
rect 29227 11336 29239 11339
rect 31110 11336 31116 11348
rect 29227 11308 31116 11336
rect 29227 11305 29239 11308
rect 29181 11299 29239 11305
rect 8496 11240 9076 11268
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5350 11160 5356 11212
rect 5408 11160 5414 11212
rect 5491 11203 5549 11209
rect 5491 11169 5503 11203
rect 5537 11200 5549 11203
rect 5718 11200 5724 11212
rect 5537 11172 5724 11200
rect 5537 11169 5549 11172
rect 5491 11163 5549 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 8294 11200 8300 11212
rect 5920 11172 8300 11200
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 5629 11135 5687 11141
rect 5629 11132 5641 11135
rect 5316 11104 5641 11132
rect 5316 11092 5322 11104
rect 5629 11101 5641 11104
rect 5675 11101 5687 11135
rect 5920 11132 5948 11172
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8570 11160 8576 11212
rect 8628 11160 8634 11212
rect 8662 11160 8668 11212
rect 8720 11160 8726 11212
rect 8754 11160 8760 11212
rect 8812 11160 8818 11212
rect 9048 11209 9076 11240
rect 9950 11228 9956 11280
rect 10008 11228 10014 11280
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 10781 11271 10839 11277
rect 10781 11268 10793 11271
rect 10100 11240 10793 11268
rect 10100 11228 10106 11240
rect 10781 11237 10793 11240
rect 10827 11237 10839 11271
rect 10781 11231 10839 11237
rect 8875 11203 8933 11209
rect 8875 11169 8887 11203
rect 8921 11169 8933 11203
rect 8875 11163 8933 11169
rect 9033 11203 9091 11209
rect 9033 11169 9045 11203
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 8890 11132 8918 11163
rect 5629 11095 5687 11101
rect 5828 11104 5948 11132
rect 8496 11104 8918 11132
rect 9048 11132 9076 11163
rect 9306 11160 9312 11212
rect 9364 11160 9370 11212
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 9916 11172 10517 11200
rect 9916 11160 9922 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 10594 11160 10600 11212
rect 10652 11160 10658 11212
rect 10796 11200 10824 11231
rect 11054 11228 11060 11280
rect 11112 11268 11118 11280
rect 15749 11271 15807 11277
rect 11112 11240 11560 11268
rect 11112 11228 11118 11240
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 10796 11172 11345 11200
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 11532 11141 11560 11240
rect 15749 11237 15761 11271
rect 15795 11268 15807 11271
rect 16362 11271 16420 11277
rect 16362 11268 16374 11271
rect 15795 11240 16374 11268
rect 15795 11237 15807 11240
rect 15749 11231 15807 11237
rect 16362 11237 16374 11240
rect 16408 11237 16420 11271
rect 20346 11268 20352 11280
rect 16362 11231 16420 11237
rect 16480 11240 20352 11268
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15436 11172 15669 11200
rect 15436 11160 15442 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 15838 11160 15844 11212
rect 15896 11160 15902 11212
rect 16114 11160 16120 11212
rect 16172 11160 16178 11212
rect 16480 11200 16508 11240
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 22097 11271 22155 11277
rect 22097 11268 22109 11271
rect 21232 11240 22109 11268
rect 21232 11228 21238 11240
rect 22097 11237 22109 11240
rect 22143 11237 22155 11271
rect 22097 11231 22155 11237
rect 22281 11271 22339 11277
rect 22281 11237 22293 11271
rect 22327 11268 22339 11271
rect 22741 11271 22799 11277
rect 22741 11268 22753 11271
rect 22327 11240 22753 11268
rect 22327 11237 22339 11240
rect 22281 11231 22339 11237
rect 22741 11237 22753 11240
rect 22787 11237 22799 11271
rect 24210 11268 24216 11280
rect 22741 11231 22799 11237
rect 23216 11240 24216 11268
rect 16224 11172 16508 11200
rect 17773 11203 17831 11209
rect 11425 11135 11483 11141
rect 9048 11104 10732 11132
rect 5828 11064 5856 11104
rect 8496 11076 8524 11104
rect 3712 11036 5856 11064
rect 8478 11024 8484 11076
rect 8536 11024 8542 11076
rect 8890 11064 8918 11104
rect 9030 11064 9036 11076
rect 8890 11036 9036 11064
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 10318 11024 10324 11076
rect 10376 11024 10382 11076
rect 4985 10999 5043 11005
rect 4985 10965 4997 10999
rect 5031 10996 5043 10999
rect 5258 10996 5264 11008
rect 5031 10968 5264 10996
rect 5031 10965 5043 10968
rect 4985 10959 5043 10965
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 8386 10956 8392 11008
rect 8444 10956 8450 11008
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 10137 10999 10195 11005
rect 10137 10996 10149 10999
rect 8996 10968 10149 10996
rect 8996 10956 9002 10968
rect 10137 10965 10149 10968
rect 10183 10996 10195 10999
rect 10410 10996 10416 11008
rect 10183 10968 10416 10996
rect 10183 10965 10195 10968
rect 10137 10959 10195 10965
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 10704 10996 10732 11104
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 10781 11067 10839 11073
rect 10781 11033 10793 11067
rect 10827 11064 10839 11067
rect 11440 11064 11468 11095
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 16224 11132 16252 11172
rect 17773 11169 17785 11203
rect 17819 11200 17831 11203
rect 18969 11203 19027 11209
rect 18969 11200 18981 11203
rect 17819 11172 18981 11200
rect 17819 11169 17831 11172
rect 17773 11163 17831 11169
rect 18969 11169 18981 11172
rect 19015 11169 19027 11203
rect 18969 11163 19027 11169
rect 21266 11160 21272 11212
rect 21324 11160 21330 11212
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11169 21511 11203
rect 21453 11163 21511 11169
rect 12768 11104 16252 11132
rect 12768 11092 12774 11104
rect 17678 11092 17684 11144
rect 17736 11092 17742 11144
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 19613 11135 19671 11141
rect 18288 11104 19564 11132
rect 18288 11092 18294 11104
rect 10827 11036 11468 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 12802 11064 12808 11076
rect 11940 11036 12808 11064
rect 11940 11024 11946 11036
rect 12802 11024 12808 11036
rect 12860 11024 12866 11076
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13538 11064 13544 11076
rect 13228 11036 13544 11064
rect 13228 11024 13234 11036
rect 13538 11024 13544 11036
rect 13596 11064 13602 11076
rect 16022 11064 16028 11076
rect 13596 11036 16028 11064
rect 13596 11024 13602 11036
rect 16022 11024 16028 11036
rect 16080 11024 16086 11076
rect 18141 11067 18199 11073
rect 18141 11033 18153 11067
rect 18187 11064 18199 11067
rect 18782 11064 18788 11076
rect 18187 11036 18788 11064
rect 18187 11033 18199 11036
rect 18141 11027 18199 11033
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 19536 11064 19564 11104
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 20254 11132 20260 11144
rect 19659 11104 20260 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 19702 11064 19708 11076
rect 19536 11036 19708 11064
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 21284 11064 21312 11160
rect 21468 11132 21496 11163
rect 22002 11160 22008 11212
rect 22060 11160 22066 11212
rect 22465 11203 22523 11209
rect 22465 11169 22477 11203
rect 22511 11200 22523 11203
rect 23216 11200 23244 11240
rect 24210 11228 24216 11240
rect 24268 11228 24274 11280
rect 25590 11228 25596 11280
rect 25648 11268 25654 11280
rect 25961 11271 26019 11277
rect 25961 11268 25973 11271
rect 25648 11240 25973 11268
rect 25648 11228 25654 11240
rect 25961 11237 25973 11240
rect 26007 11237 26019 11271
rect 28828 11268 28856 11296
rect 25961 11231 26019 11237
rect 28552 11240 28856 11268
rect 22511 11172 23244 11200
rect 22511 11169 22523 11172
rect 22465 11163 22523 11169
rect 22094 11132 22100 11144
rect 21468 11104 22100 11132
rect 22094 11092 22100 11104
rect 22152 11092 22158 11144
rect 22480 11064 22508 11163
rect 23290 11160 23296 11212
rect 23348 11160 23354 11212
rect 23477 11203 23535 11209
rect 23477 11169 23489 11203
rect 23523 11200 23535 11203
rect 23566 11200 23572 11212
rect 23523 11172 23572 11200
rect 23523 11169 23535 11172
rect 23477 11163 23535 11169
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 23750 11209 23756 11212
rect 23744 11163 23756 11209
rect 23750 11160 23756 11163
rect 23808 11160 23814 11212
rect 25976 11132 26004 11231
rect 28077 11203 28135 11209
rect 28077 11169 28089 11203
rect 28123 11200 28135 11203
rect 28166 11200 28172 11212
rect 28123 11172 28172 11200
rect 28123 11169 28135 11172
rect 28077 11163 28135 11169
rect 28166 11160 28172 11172
rect 28224 11160 28230 11212
rect 28552 11209 28580 11240
rect 28537 11203 28595 11209
rect 28537 11169 28549 11203
rect 28583 11169 28595 11203
rect 28537 11163 28595 11169
rect 28813 11203 28871 11209
rect 28813 11169 28825 11203
rect 28859 11200 28871 11203
rect 28902 11200 28908 11212
rect 28859 11172 28908 11200
rect 28859 11169 28871 11172
rect 28813 11163 28871 11169
rect 28902 11160 28908 11172
rect 28960 11160 28966 11212
rect 29086 11160 29092 11212
rect 29144 11160 29150 11212
rect 27985 11135 28043 11141
rect 25976 11104 27936 11132
rect 21284 11036 22508 11064
rect 25314 11024 25320 11076
rect 25372 11064 25378 11076
rect 25593 11067 25651 11073
rect 25593 11064 25605 11067
rect 25372 11036 25605 11064
rect 25372 11024 25378 11036
rect 25593 11033 25605 11036
rect 25639 11033 25651 11067
rect 25593 11027 25651 11033
rect 27614 11024 27620 11076
rect 27672 11064 27678 11076
rect 27709 11067 27767 11073
rect 27709 11064 27721 11067
rect 27672 11036 27721 11064
rect 27672 11024 27678 11036
rect 27709 11033 27721 11036
rect 27755 11033 27767 11067
rect 27709 11027 27767 11033
rect 11330 10996 11336 11008
rect 10704 10968 11336 10996
rect 11330 10956 11336 10968
rect 11388 10996 11394 11008
rect 12986 10996 12992 11008
rect 11388 10968 12992 10996
rect 11388 10956 11394 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 16758 10956 16764 11008
rect 16816 10996 16822 11008
rect 17497 10999 17555 11005
rect 17497 10996 17509 10999
rect 16816 10968 17509 10996
rect 16816 10956 16822 10968
rect 17497 10965 17509 10968
rect 17543 10965 17555 10999
rect 17497 10959 17555 10965
rect 21637 10999 21695 11005
rect 21637 10965 21649 10999
rect 21683 10996 21695 10999
rect 21726 10996 21732 11008
rect 21683 10968 21732 10996
rect 21683 10965 21695 10968
rect 21637 10959 21695 10965
rect 21726 10956 21732 10968
rect 21784 10956 21790 11008
rect 24854 10956 24860 11008
rect 24912 10996 24918 11008
rect 26142 10996 26148 11008
rect 24912 10968 26148 10996
rect 24912 10956 24918 10968
rect 26142 10956 26148 10968
rect 26200 10956 26206 11008
rect 27908 10996 27936 11104
rect 27985 11101 27997 11135
rect 28031 11101 28043 11135
rect 27985 11095 28043 11101
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11132 28779 11135
rect 29196 11132 29224 11299
rect 31110 11296 31116 11308
rect 31168 11296 31174 11348
rect 29914 11228 29920 11280
rect 29972 11268 29978 11280
rect 29972 11240 30604 11268
rect 29972 11228 29978 11240
rect 30006 11160 30012 11212
rect 30064 11200 30070 11212
rect 30576 11209 30604 11240
rect 30294 11203 30352 11209
rect 30294 11200 30306 11203
rect 30064 11172 30306 11200
rect 30064 11160 30070 11172
rect 30294 11169 30306 11172
rect 30340 11169 30352 11203
rect 30294 11163 30352 11169
rect 30561 11203 30619 11209
rect 30561 11169 30573 11203
rect 30607 11169 30619 11203
rect 30561 11163 30619 11169
rect 30742 11160 30748 11212
rect 30800 11160 30806 11212
rect 28767 11104 29224 11132
rect 28767 11101 28779 11104
rect 28721 11095 28779 11101
rect 28000 11064 28028 11095
rect 29546 11064 29552 11076
rect 28000 11036 29552 11064
rect 29546 11024 29552 11036
rect 29604 11024 29610 11076
rect 28534 10996 28540 11008
rect 27908 10968 28540 10996
rect 28534 10956 28540 10968
rect 28592 10956 28598 11008
rect 28994 10956 29000 11008
rect 29052 10956 29058 11008
rect 31294 10956 31300 11008
rect 31352 10956 31358 11008
rect 552 10906 31648 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 11436 10906
rect 11488 10854 11500 10906
rect 11552 10854 11564 10906
rect 11616 10854 11628 10906
rect 11680 10854 11692 10906
rect 11744 10854 19210 10906
rect 19262 10854 19274 10906
rect 19326 10854 19338 10906
rect 19390 10854 19402 10906
rect 19454 10854 19466 10906
rect 19518 10854 26984 10906
rect 27036 10854 27048 10906
rect 27100 10854 27112 10906
rect 27164 10854 27176 10906
rect 27228 10854 27240 10906
rect 27292 10854 31648 10906
rect 552 10832 31648 10854
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 2590 10792 2596 10804
rect 2547 10764 2596 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 5166 10792 5172 10804
rect 3108 10764 5172 10792
rect 3108 10752 3114 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 6086 10792 6092 10804
rect 5491 10764 6092 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 6788 10764 7389 10792
rect 6788 10752 6794 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 8754 10752 8760 10804
rect 8812 10752 8818 10804
rect 12618 10752 12624 10804
rect 12676 10792 12682 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12676 10764 13185 10792
rect 12676 10752 12682 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 15838 10752 15844 10804
rect 15896 10752 15902 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 20438 10792 20444 10804
rect 18288 10764 20444 10792
rect 18288 10752 18294 10764
rect 20438 10752 20444 10764
rect 20496 10792 20502 10804
rect 20714 10792 20720 10804
rect 20496 10764 20720 10792
rect 20496 10752 20502 10764
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 22094 10752 22100 10804
rect 22152 10752 22158 10804
rect 23385 10795 23443 10801
rect 23385 10761 23397 10795
rect 23431 10792 23443 10795
rect 23750 10792 23756 10804
rect 23431 10764 23756 10792
rect 23431 10761 23443 10764
rect 23385 10755 23443 10761
rect 23750 10752 23756 10764
rect 23808 10752 23814 10804
rect 25866 10752 25872 10804
rect 25924 10752 25930 10804
rect 29917 10795 29975 10801
rect 29917 10761 29929 10795
rect 29963 10792 29975 10795
rect 30006 10792 30012 10804
rect 29963 10764 30012 10792
rect 29963 10761 29975 10764
rect 29917 10755 29975 10761
rect 30006 10752 30012 10764
rect 30064 10752 30070 10804
rect 30653 10795 30711 10801
rect 30653 10761 30665 10795
rect 30699 10761 30711 10795
rect 30653 10755 30711 10761
rect 7190 10684 7196 10736
rect 7248 10724 7254 10736
rect 8846 10724 8852 10736
rect 7248 10696 8852 10724
rect 7248 10684 7254 10696
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 18690 10724 18696 10736
rect 12268 10696 18696 10724
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 2924 10628 5089 10656
rect 2924 10616 2930 10628
rect 5077 10625 5089 10628
rect 5123 10656 5135 10659
rect 8938 10656 8944 10668
rect 5123 10628 5948 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 2038 10548 2044 10600
rect 2096 10588 2102 10600
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 2096 10560 2237 10588
rect 2096 10548 2102 10560
rect 2225 10557 2237 10560
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10588 2743 10591
rect 2774 10588 2780 10600
rect 2731 10560 2780 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 5258 10548 5264 10600
rect 5316 10548 5322 10600
rect 5534 10548 5540 10600
rect 5592 10548 5598 10600
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10588 5687 10591
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5675 10560 5825 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 5813 10557 5825 10560
rect 5859 10557 5871 10591
rect 5920 10588 5948 10628
rect 7576 10628 8944 10656
rect 7576 10597 7604 10628
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 5920 10560 6316 10588
rect 5813 10551 5871 10557
rect 6288 10532 6316 10560
rect 6472 10560 7573 10588
rect 6472 10532 6500 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8018 10588 8024 10600
rect 7883 10560 8024 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 4154 10480 4160 10532
rect 4212 10520 4218 10532
rect 4798 10520 4804 10532
rect 4212 10492 4804 10520
rect 4212 10480 4218 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 5902 10480 5908 10532
rect 5960 10520 5966 10532
rect 6058 10523 6116 10529
rect 6058 10520 6070 10523
rect 5960 10492 6070 10520
rect 5960 10480 5966 10492
rect 6058 10489 6070 10492
rect 6104 10489 6116 10523
rect 6058 10483 6116 10489
rect 6270 10480 6276 10532
rect 6328 10480 6334 10532
rect 6454 10480 6460 10532
rect 6512 10480 6518 10532
rect 7852 10520 7880 10551
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 9490 10548 9496 10600
rect 9548 10548 9554 10600
rect 9674 10548 9680 10600
rect 9732 10548 9738 10600
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 11790 10588 11796 10600
rect 10284 10560 11796 10588
rect 10284 10548 10290 10560
rect 11790 10548 11796 10560
rect 11848 10588 11854 10600
rect 12158 10588 12164 10600
rect 11848 10560 12164 10588
rect 11848 10548 11854 10560
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 12268 10597 12296 10696
rect 18690 10684 18696 10696
rect 18748 10684 18754 10736
rect 22112 10724 22140 10752
rect 22112 10696 26004 10724
rect 15378 10616 15384 10668
rect 15436 10616 15442 10668
rect 15930 10616 15936 10668
rect 15988 10656 15994 10668
rect 16390 10656 16396 10668
rect 15988 10628 16396 10656
rect 15988 10616 15994 10628
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12526 10548 12532 10600
rect 12584 10548 12590 10600
rect 12802 10548 12808 10600
rect 12860 10597 12866 10600
rect 12860 10591 12889 10597
rect 12877 10557 12889 10591
rect 12860 10551 12889 10557
rect 12860 10548 12866 10551
rect 12986 10548 12992 10600
rect 13044 10548 13050 10600
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 7208 10492 7880 10520
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 2004 10424 2145 10452
rect 2004 10412 2010 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 7208 10452 7236 10492
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12345 10523 12403 10529
rect 12345 10520 12357 10523
rect 12032 10492 12357 10520
rect 12032 10480 12038 10492
rect 12345 10489 12357 10492
rect 12391 10489 12403 10523
rect 12345 10483 12403 10489
rect 12434 10480 12440 10532
rect 12492 10520 12498 10532
rect 12621 10523 12679 10529
rect 12621 10520 12633 10523
rect 12492 10492 12633 10520
rect 12492 10480 12498 10492
rect 12621 10489 12633 10492
rect 12667 10489 12679 10523
rect 12621 10483 12679 10489
rect 12710 10480 12716 10532
rect 12768 10480 12774 10532
rect 13280 10520 13308 10551
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 14056 10560 14105 10588
rect 14056 10548 14062 10560
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 13722 10520 13728 10532
rect 13280 10492 13728 10520
rect 5592 10424 7236 10452
rect 5592 10412 5598 10424
rect 7742 10412 7748 10464
rect 7800 10412 7806 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9824 10424 9873 10452
rect 9824 10412 9830 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 9861 10415 9919 10421
rect 10042 10412 10048 10464
rect 10100 10452 10106 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 10100 10424 10149 10452
rect 10100 10412 10106 10424
rect 10137 10421 10149 10424
rect 10183 10421 10195 10455
rect 10137 10415 10195 10421
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 11698 10452 11704 10464
rect 10468 10424 11704 10452
rect 10468 10412 10474 10424
rect 11698 10412 11704 10424
rect 11756 10452 11762 10464
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 11756 10424 12081 10452
rect 11756 10412 11762 10424
rect 12069 10421 12081 10424
rect 12115 10421 12127 10455
rect 12069 10415 12127 10421
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 13280 10452 13308 10492
rect 13722 10480 13728 10492
rect 13780 10520 13786 10532
rect 14660 10520 14688 10551
rect 15194 10548 15200 10600
rect 15252 10548 15258 10600
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16224 10597 16252 10628
rect 16390 10616 16396 10628
rect 16448 10616 16454 10668
rect 16482 10616 16488 10668
rect 16540 10616 16546 10668
rect 23845 10659 23903 10665
rect 23845 10656 23857 10659
rect 22940 10628 23857 10656
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16758 10548 16764 10600
rect 16816 10548 16822 10600
rect 18230 10548 18236 10600
rect 18288 10548 18294 10600
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 13780 10492 14688 10520
rect 16117 10523 16175 10529
rect 13780 10480 13786 10492
rect 16117 10489 16129 10523
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 12216 10424 13308 10452
rect 12216 10412 12222 10424
rect 13538 10412 13544 10464
rect 13596 10412 13602 10464
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 14608 10424 14749 10452
rect 14608 10412 14614 10424
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 14737 10415 14795 10421
rect 15010 10412 15016 10464
rect 15068 10412 15074 10464
rect 16132 10452 16160 10483
rect 16298 10480 16304 10532
rect 16356 10529 16362 10532
rect 16356 10523 16385 10529
rect 16373 10520 16385 10523
rect 18322 10520 18328 10532
rect 16373 10492 18328 10520
rect 16373 10489 16385 10492
rect 16356 10483 16385 10489
rect 16356 10480 16362 10483
rect 18322 10480 18328 10492
rect 18380 10520 18386 10532
rect 18432 10520 18460 10551
rect 18690 10548 18696 10600
rect 18748 10548 18754 10600
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 18949 10591 19007 10597
rect 18949 10588 18961 10591
rect 18840 10560 18961 10588
rect 18840 10548 18846 10560
rect 18949 10557 18961 10560
rect 18995 10557 19007 10591
rect 18949 10551 19007 10557
rect 20438 10548 20444 10600
rect 20496 10548 20502 10600
rect 20533 10591 20591 10597
rect 20533 10557 20545 10591
rect 20579 10588 20591 10591
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20579 10560 20729 10588
rect 20579 10557 20591 10560
rect 20533 10551 20591 10557
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 22741 10591 22799 10597
rect 22741 10557 22753 10591
rect 22787 10588 22799 10591
rect 22830 10588 22836 10600
rect 22787 10560 22836 10588
rect 22787 10557 22799 10560
rect 22741 10551 22799 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 22940 10597 22968 10628
rect 23845 10625 23857 10628
rect 23891 10625 23903 10659
rect 23845 10619 23903 10625
rect 22925 10591 22983 10597
rect 22925 10557 22937 10591
rect 22971 10557 22983 10591
rect 22925 10551 22983 10557
rect 23017 10591 23075 10597
rect 23017 10557 23029 10591
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 19058 10520 19064 10532
rect 18380 10492 19064 10520
rect 18380 10480 18386 10492
rect 19058 10480 19064 10492
rect 19116 10480 19122 10532
rect 20984 10523 21042 10529
rect 20984 10489 20996 10523
rect 21030 10520 21042 10523
rect 21266 10520 21272 10532
rect 21030 10492 21272 10520
rect 21030 10489 21042 10492
rect 20984 10483 21042 10489
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 21450 10480 21456 10532
rect 21508 10520 21514 10532
rect 22002 10520 22008 10532
rect 21508 10492 22008 10520
rect 21508 10480 21514 10492
rect 22002 10480 22008 10492
rect 22060 10520 22066 10532
rect 23032 10520 23060 10551
rect 23106 10548 23112 10600
rect 23164 10548 23170 10600
rect 24029 10591 24087 10597
rect 24029 10557 24041 10591
rect 24075 10588 24087 10591
rect 24854 10588 24860 10600
rect 24075 10560 24860 10588
rect 24075 10557 24087 10560
rect 24029 10551 24087 10557
rect 24854 10548 24860 10560
rect 24912 10548 24918 10600
rect 25317 10591 25375 10597
rect 25317 10557 25329 10591
rect 25363 10557 25375 10591
rect 25317 10551 25375 10557
rect 22060 10492 23060 10520
rect 22060 10480 22066 10492
rect 24210 10480 24216 10532
rect 24268 10480 24274 10532
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16132 10424 16681 10452
rect 16669 10421 16681 10424
rect 16715 10452 16727 10455
rect 16758 10452 16764 10464
rect 16715 10424 16764 10452
rect 16715 10421 16727 10424
rect 16669 10415 16727 10421
rect 16758 10412 16764 10424
rect 16816 10412 16822 10464
rect 17954 10412 17960 10464
rect 18012 10452 18018 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 18012 10424 18245 10452
rect 18012 10412 18018 10424
rect 18233 10421 18245 10424
rect 18279 10452 18291 10455
rect 18966 10452 18972 10464
rect 18279 10424 18972 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 20073 10455 20131 10461
rect 20073 10421 20085 10455
rect 20119 10452 20131 10455
rect 20254 10452 20260 10464
rect 20119 10424 20260 10452
rect 20119 10421 20131 10424
rect 20073 10415 20131 10421
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 25332 10452 25360 10551
rect 25424 10520 25452 10696
rect 25866 10656 25872 10668
rect 25516 10628 25872 10656
rect 25516 10597 25544 10628
rect 25866 10616 25872 10628
rect 25924 10616 25930 10668
rect 25976 10597 26004 10696
rect 29546 10684 29552 10736
rect 29604 10724 29610 10736
rect 30469 10727 30527 10733
rect 30469 10724 30481 10727
rect 29604 10696 30481 10724
rect 29604 10684 29610 10696
rect 30469 10693 30481 10696
rect 30515 10693 30527 10727
rect 30668 10724 30696 10755
rect 30926 10752 30932 10804
rect 30984 10792 30990 10804
rect 31205 10795 31263 10801
rect 31205 10792 31217 10795
rect 30984 10764 31217 10792
rect 30984 10752 30990 10764
rect 31205 10761 31217 10764
rect 31251 10761 31263 10795
rect 31205 10755 31263 10761
rect 30668 10696 31064 10724
rect 30469 10687 30527 10693
rect 26053 10659 26111 10665
rect 26053 10625 26065 10659
rect 26099 10656 26111 10659
rect 28994 10656 29000 10668
rect 26099 10628 29000 10656
rect 26099 10625 26111 10628
rect 26053 10619 26111 10625
rect 25501 10591 25559 10597
rect 25501 10557 25513 10591
rect 25547 10557 25559 10591
rect 25501 10551 25559 10557
rect 25685 10591 25743 10597
rect 25685 10557 25697 10591
rect 25731 10557 25743 10591
rect 25685 10551 25743 10557
rect 25961 10591 26019 10597
rect 25961 10557 25973 10591
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 25593 10523 25651 10529
rect 25593 10520 25605 10523
rect 25424 10492 25605 10520
rect 25593 10489 25605 10492
rect 25639 10489 25651 10523
rect 25700 10520 25728 10551
rect 26068 10520 26096 10619
rect 28994 10616 29000 10628
rect 29052 10656 29058 10668
rect 29052 10628 29776 10656
rect 29052 10616 29058 10628
rect 26142 10548 26148 10600
rect 26200 10588 26206 10600
rect 26237 10591 26295 10597
rect 26237 10588 26249 10591
rect 26200 10560 26249 10588
rect 26200 10548 26206 10560
rect 26237 10557 26249 10560
rect 26283 10557 26295 10591
rect 26237 10551 26295 10557
rect 26326 10548 26332 10600
rect 26384 10548 26390 10600
rect 28902 10548 28908 10600
rect 28960 10588 28966 10600
rect 29641 10591 29699 10597
rect 29641 10588 29653 10591
rect 28960 10560 29653 10588
rect 28960 10548 28966 10560
rect 29641 10557 29653 10560
rect 29687 10557 29699 10591
rect 29748 10588 29776 10628
rect 30098 10616 30104 10668
rect 30156 10656 30162 10668
rect 30156 10628 30972 10656
rect 30156 10616 30162 10628
rect 30193 10591 30251 10597
rect 30193 10588 30205 10591
rect 29748 10560 30205 10588
rect 29641 10551 29699 10557
rect 30193 10557 30205 10560
rect 30239 10557 30251 10591
rect 30193 10551 30251 10557
rect 30668 10529 30696 10628
rect 30944 10597 30972 10628
rect 31036 10597 31064 10696
rect 30929 10591 30987 10597
rect 30929 10557 30941 10591
rect 30975 10557 30987 10591
rect 30929 10551 30987 10557
rect 31021 10591 31079 10597
rect 31021 10557 31033 10591
rect 31067 10588 31079 10591
rect 31110 10588 31116 10600
rect 31067 10560 31116 10588
rect 31067 10557 31079 10560
rect 31021 10551 31079 10557
rect 31110 10548 31116 10560
rect 31168 10548 31174 10600
rect 31205 10591 31263 10597
rect 31205 10557 31217 10591
rect 31251 10588 31263 10591
rect 31294 10588 31300 10600
rect 31251 10560 31300 10588
rect 31251 10557 31263 10560
rect 31205 10551 31263 10557
rect 31294 10548 31300 10560
rect 31352 10548 31358 10600
rect 25700 10492 26096 10520
rect 30637 10523 30696 10529
rect 25593 10483 25651 10489
rect 30637 10489 30649 10523
rect 30683 10492 30696 10523
rect 30683 10489 30695 10492
rect 30637 10483 30695 10489
rect 30742 10480 30748 10532
rect 30800 10520 30806 10532
rect 30837 10523 30895 10529
rect 30837 10520 30849 10523
rect 30800 10492 30849 10520
rect 30800 10480 30806 10492
rect 30837 10489 30849 10492
rect 30883 10489 30895 10523
rect 30837 10483 30895 10489
rect 26513 10455 26571 10461
rect 26513 10452 26525 10455
rect 25332 10424 26525 10452
rect 26513 10421 26525 10424
rect 26559 10421 26571 10455
rect 26513 10415 26571 10421
rect 28626 10412 28632 10464
rect 28684 10452 28690 10464
rect 29089 10455 29147 10461
rect 29089 10452 29101 10455
rect 28684 10424 29101 10452
rect 28684 10412 28690 10424
rect 29089 10421 29101 10424
rect 29135 10421 29147 10455
rect 29089 10415 29147 10421
rect 552 10362 31648 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 12096 10362
rect 12148 10310 12160 10362
rect 12212 10310 12224 10362
rect 12276 10310 12288 10362
rect 12340 10310 12352 10362
rect 12404 10310 19870 10362
rect 19922 10310 19934 10362
rect 19986 10310 19998 10362
rect 20050 10310 20062 10362
rect 20114 10310 20126 10362
rect 20178 10310 27644 10362
rect 27696 10310 27708 10362
rect 27760 10310 27772 10362
rect 27824 10310 27836 10362
rect 27888 10310 27900 10362
rect 27952 10310 31648 10362
rect 552 10288 31648 10310
rect 5902 10208 5908 10260
rect 5960 10208 5966 10260
rect 7190 10248 7196 10260
rect 6656 10220 7196 10248
rect 2038 10180 2044 10192
rect 1688 10152 2044 10180
rect 1688 10121 1716 10152
rect 2038 10140 2044 10152
rect 2096 10140 2102 10192
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 3927 10183 3985 10189
rect 3568 10152 3832 10180
rect 3568 10140 3574 10152
rect 3804 10124 3832 10152
rect 3927 10149 3939 10183
rect 3973 10180 3985 10183
rect 4430 10180 4436 10192
rect 3973 10152 4436 10180
rect 3973 10149 3985 10152
rect 3927 10143 3985 10149
rect 4430 10140 4436 10152
rect 4488 10140 4494 10192
rect 4706 10140 4712 10192
rect 4764 10180 4770 10192
rect 5350 10180 5356 10192
rect 4764 10152 5356 10180
rect 4764 10140 4770 10152
rect 5350 10140 5356 10152
rect 5408 10180 5414 10192
rect 6454 10180 6460 10192
rect 5408 10152 6460 10180
rect 5408 10140 5414 10152
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 6656 10189 6684 10220
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9306 10248 9312 10260
rect 8619 10220 9312 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 13538 10248 13544 10260
rect 12176 10220 13544 10248
rect 6641 10183 6699 10189
rect 6641 10149 6653 10183
rect 6687 10149 6699 10183
rect 6641 10143 6699 10149
rect 6822 10140 6828 10192
rect 6880 10189 6886 10192
rect 6880 10183 6909 10189
rect 6897 10149 6909 10183
rect 7742 10180 7748 10192
rect 6880 10143 6909 10149
rect 7208 10152 7748 10180
rect 6880 10140 6886 10143
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10081 1731 10115
rect 1673 10075 1731 10081
rect 1946 10072 1952 10124
rect 2004 10072 2010 10124
rect 2205 10115 2263 10121
rect 2205 10112 2217 10115
rect 2056 10084 2217 10112
rect 1578 10004 1584 10056
rect 1636 10044 1642 10056
rect 2056 10044 2084 10084
rect 2205 10081 2217 10084
rect 2251 10081 2263 10115
rect 2205 10075 2263 10081
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 3605 10115 3663 10121
rect 3605 10112 3617 10115
rect 3016 10084 3617 10112
rect 3016 10072 3022 10084
rect 3605 10081 3617 10084
rect 3651 10081 3663 10115
rect 3605 10075 3663 10081
rect 3694 10072 3700 10124
rect 3752 10072 3758 10124
rect 3786 10072 3792 10124
rect 3844 10072 3850 10124
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 4246 10112 4252 10124
rect 4111 10084 4252 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 6135 10084 6377 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6546 10072 6552 10124
rect 6604 10072 6610 10124
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 7208 10121 7236 10152
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 8662 10140 8668 10192
rect 8720 10180 8726 10192
rect 8720 10152 10548 10180
rect 8720 10140 8726 10152
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7282 10072 7288 10124
rect 7340 10072 7346 10124
rect 7460 10115 7518 10121
rect 7460 10081 7472 10115
rect 7506 10112 7518 10115
rect 8386 10112 8392 10124
rect 7506 10084 8392 10112
rect 7506 10081 7518 10084
rect 7460 10075 7518 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 9766 10072 9772 10124
rect 9824 10121 9830 10124
rect 9824 10112 9836 10121
rect 9824 10084 9869 10112
rect 9824 10075 9836 10084
rect 9824 10072 9830 10075
rect 10042 10072 10048 10124
rect 10100 10072 10106 10124
rect 1636 10016 2084 10044
rect 1636 10004 1642 10016
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 6270 10044 6276 10056
rect 4396 10016 6276 10044
rect 4396 10004 4402 10016
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 3786 9936 3792 9988
rect 3844 9976 3850 9988
rect 6748 9976 6776 10072
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 7300 10044 7328 10072
rect 7055 10016 7328 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 3844 9948 6776 9976
rect 10520 9976 10548 10152
rect 10962 10140 10968 10192
rect 11020 10180 11026 10192
rect 12066 10189 12072 10192
rect 12023 10183 12072 10189
rect 12023 10180 12035 10183
rect 11020 10152 12035 10180
rect 11020 10140 11026 10152
rect 12023 10149 12035 10152
rect 12069 10149 12072 10183
rect 12023 10143 12072 10149
rect 12066 10140 12072 10143
rect 12124 10140 12130 10192
rect 12176 10189 12204 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13998 10248 14004 10260
rect 13688 10220 14004 10248
rect 13688 10208 13694 10220
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 18414 10248 18420 10260
rect 18156 10220 18420 10248
rect 12161 10183 12219 10189
rect 12161 10149 12173 10183
rect 12207 10149 12219 10183
rect 12434 10180 12440 10192
rect 12161 10143 12219 10149
rect 12268 10152 12440 10180
rect 11146 10072 11152 10124
rect 11204 10072 11210 10124
rect 11238 10072 11244 10124
rect 11296 10112 11302 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11296 10084 11437 10112
rect 11296 10072 11302 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 11609 10115 11667 10121
rect 11609 10081 11621 10115
rect 11655 10112 11667 10115
rect 11698 10112 11704 10124
rect 11655 10084 11704 10112
rect 11655 10081 11667 10084
rect 11609 10075 11667 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 12268 10121 12296 10152
rect 12434 10140 12440 10152
rect 12492 10140 12498 10192
rect 12866 10183 12924 10189
rect 12866 10149 12878 10183
rect 12912 10180 12924 10183
rect 14820 10183 14878 10189
rect 12912 10149 12931 10180
rect 12866 10143 12931 10149
rect 14820 10149 14832 10183
rect 14866 10180 14878 10183
rect 15010 10180 15016 10192
rect 14866 10152 15016 10180
rect 14866 10149 14878 10152
rect 14820 10143 14878 10149
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 11992 10084 12265 10112
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 11388 10016 11897 10044
rect 11388 10004 11394 10016
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 10520 9948 11100 9976
rect 3844 9936 3850 9948
rect 1762 9868 1768 9920
rect 1820 9868 1826 9920
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 3329 9911 3387 9917
rect 3329 9908 3341 9911
rect 3292 9880 3341 9908
rect 3292 9868 3298 9880
rect 3329 9877 3341 9880
rect 3375 9877 3387 9911
rect 3329 9871 3387 9877
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 3694 9908 3700 9920
rect 3568 9880 3700 9908
rect 3568 9868 3574 9880
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6822 9908 6828 9920
rect 5776 9880 6828 9908
rect 5776 9868 5782 9880
rect 6822 9868 6828 9880
rect 6880 9908 6886 9920
rect 8478 9908 8484 9920
rect 6880 9880 8484 9908
rect 6880 9868 6886 9880
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 8665 9911 8723 9917
rect 8665 9877 8677 9911
rect 8711 9908 8723 9911
rect 8754 9908 8760 9920
rect 8711 9880 8760 9908
rect 8711 9877 8723 9880
rect 8665 9871 8723 9877
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 10965 9911 11023 9917
rect 10965 9908 10977 9911
rect 10836 9880 10977 9908
rect 10836 9868 10842 9880
rect 10965 9877 10977 9880
rect 11011 9877 11023 9911
rect 11072 9908 11100 9948
rect 11793 9911 11851 9917
rect 11793 9908 11805 9911
rect 11072 9880 11805 9908
rect 10965 9871 11023 9877
rect 11793 9877 11805 9880
rect 11839 9908 11851 9911
rect 11992 9908 12020 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 12342 10072 12348 10124
rect 12400 10072 12406 10124
rect 12618 10072 12624 10124
rect 12676 10072 12682 10124
rect 12903 10112 12931 10143
rect 15010 10140 15016 10152
rect 15068 10140 15074 10192
rect 18156 10189 18184 10220
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18748 10220 18889 10248
rect 18748 10208 18754 10220
rect 18877 10217 18889 10220
rect 18923 10217 18935 10251
rect 18877 10211 18935 10217
rect 21266 10208 21272 10260
rect 21324 10208 21330 10260
rect 25685 10251 25743 10257
rect 25685 10217 25697 10251
rect 25731 10217 25743 10251
rect 25685 10211 25743 10217
rect 18322 10189 18328 10192
rect 18141 10183 18199 10189
rect 18141 10149 18153 10183
rect 18187 10149 18199 10183
rect 18141 10143 18199 10149
rect 18279 10183 18328 10189
rect 18279 10149 18291 10183
rect 18325 10149 18328 10183
rect 18279 10143 18328 10149
rect 18322 10140 18328 10143
rect 18380 10140 18386 10192
rect 20438 10180 20444 10192
rect 18984 10152 20444 10180
rect 12719 10084 12931 10112
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 12719 10044 12747 10084
rect 14550 10072 14556 10124
rect 14608 10072 14614 10124
rect 16022 10072 16028 10124
rect 16080 10112 16086 10124
rect 17954 10112 17960 10124
rect 16080 10084 17960 10112
rect 16080 10072 16086 10084
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18046 10072 18052 10124
rect 18104 10072 18110 10124
rect 18874 10072 18880 10124
rect 18932 10112 18938 10124
rect 18984 10121 19012 10152
rect 20438 10140 20444 10152
rect 20496 10180 20502 10192
rect 20496 10152 22094 10180
rect 20496 10140 20502 10152
rect 18969 10115 19027 10121
rect 18969 10112 18981 10115
rect 18932 10084 18981 10112
rect 18932 10072 18938 10084
rect 18969 10081 18981 10084
rect 19015 10081 19027 10115
rect 18969 10075 19027 10081
rect 21542 10072 21548 10124
rect 21600 10072 21606 10124
rect 21637 10115 21695 10121
rect 21637 10081 21649 10115
rect 21683 10081 21695 10115
rect 21637 10075 21695 10081
rect 12575 10016 12747 10044
rect 18417 10047 18475 10053
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 18417 10013 18429 10047
rect 18463 10044 18475 10047
rect 21358 10044 21364 10056
rect 18463 10016 21364 10044
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 21652 10044 21680 10075
rect 21726 10072 21732 10124
rect 21784 10072 21790 10124
rect 21910 10072 21916 10124
rect 21968 10072 21974 10124
rect 22066 10112 22094 10152
rect 22370 10140 22376 10192
rect 22428 10180 22434 10192
rect 22465 10183 22523 10189
rect 22465 10180 22477 10183
rect 22428 10152 22477 10180
rect 22428 10140 22434 10152
rect 22465 10149 22477 10152
rect 22511 10180 22523 10183
rect 24210 10180 24216 10192
rect 22511 10152 24216 10180
rect 22511 10149 22523 10152
rect 22465 10143 22523 10149
rect 24210 10140 24216 10152
rect 24268 10140 24274 10192
rect 24854 10140 24860 10192
rect 24912 10180 24918 10192
rect 25409 10183 25467 10189
rect 25409 10180 25421 10183
rect 24912 10152 25421 10180
rect 24912 10140 24918 10152
rect 25409 10149 25421 10152
rect 25455 10149 25467 10183
rect 25700 10180 25728 10211
rect 25866 10208 25872 10260
rect 25924 10248 25930 10260
rect 26237 10251 26295 10257
rect 26237 10248 26249 10251
rect 25924 10220 26249 10248
rect 25924 10208 25930 10220
rect 26237 10217 26249 10220
rect 26283 10217 26295 10251
rect 26237 10211 26295 10217
rect 26326 10208 26332 10260
rect 26384 10248 26390 10260
rect 26881 10251 26939 10257
rect 26881 10248 26893 10251
rect 26384 10220 26893 10248
rect 26384 10208 26390 10220
rect 26881 10217 26893 10220
rect 26927 10217 26939 10251
rect 26881 10211 26939 10217
rect 29273 10251 29331 10257
rect 29273 10217 29285 10251
rect 29319 10248 29331 10251
rect 30098 10248 30104 10260
rect 29319 10220 30104 10248
rect 29319 10217 29331 10220
rect 29273 10211 29331 10217
rect 30098 10208 30104 10220
rect 30156 10248 30162 10260
rect 30282 10248 30288 10260
rect 30156 10220 30288 10248
rect 30156 10208 30162 10220
rect 30282 10208 30288 10220
rect 30340 10208 30346 10260
rect 25700 10152 26096 10180
rect 25409 10143 25467 10149
rect 22189 10115 22247 10121
rect 22189 10112 22201 10115
rect 22066 10084 22201 10112
rect 22189 10081 22201 10084
rect 22235 10081 22247 10115
rect 22189 10075 22247 10081
rect 22649 10115 22707 10121
rect 22649 10081 22661 10115
rect 22695 10112 22707 10115
rect 23474 10112 23480 10124
rect 22695 10084 23480 10112
rect 22695 10081 22707 10084
rect 22649 10075 22707 10081
rect 23474 10072 23480 10084
rect 23532 10112 23538 10124
rect 25038 10112 25044 10124
rect 23532 10084 25044 10112
rect 23532 10072 23538 10084
rect 25038 10072 25044 10084
rect 25096 10112 25102 10124
rect 25133 10115 25191 10121
rect 25133 10112 25145 10115
rect 25096 10084 25145 10112
rect 25096 10072 25102 10084
rect 25133 10081 25145 10084
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 25317 10115 25375 10121
rect 25317 10081 25329 10115
rect 25363 10112 25375 10115
rect 25501 10115 25559 10121
rect 25363 10084 25452 10112
rect 25363 10081 25375 10084
rect 25317 10075 25375 10081
rect 22002 10044 22008 10056
rect 21652 10016 22008 10044
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 11839 9880 12020 9908
rect 11839 9877 11851 9880
rect 11793 9871 11851 9877
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 15470 9908 15476 9920
rect 12492 9880 15476 9908
rect 12492 9868 12498 9880
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15933 9911 15991 9917
rect 15933 9877 15945 9911
rect 15979 9908 15991 9911
rect 16206 9908 16212 9920
rect 15979 9880 16212 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 16850 9868 16856 9920
rect 16908 9908 16914 9920
rect 17773 9911 17831 9917
rect 17773 9908 17785 9911
rect 16908 9880 17785 9908
rect 16908 9868 16914 9880
rect 17773 9877 17785 9880
rect 17819 9877 17831 9911
rect 17773 9871 17831 9877
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22281 9911 22339 9917
rect 22281 9908 22293 9911
rect 22152 9880 22293 9908
rect 22152 9868 22158 9880
rect 22281 9877 22293 9880
rect 22327 9877 22339 9911
rect 22281 9871 22339 9877
rect 22833 9911 22891 9917
rect 22833 9877 22845 9911
rect 22879 9908 22891 9911
rect 22922 9908 22928 9920
rect 22879 9880 22928 9908
rect 22879 9877 22891 9880
rect 22833 9871 22891 9877
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 25130 9868 25136 9920
rect 25188 9908 25194 9920
rect 25424 9908 25452 10084
rect 25501 10081 25513 10115
rect 25547 10081 25559 10115
rect 25501 10075 25559 10081
rect 25516 9976 25544 10075
rect 25774 10072 25780 10124
rect 25832 10072 25838 10124
rect 25866 10072 25872 10124
rect 25924 10072 25930 10124
rect 26068 10121 26096 10152
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10081 26111 10115
rect 26053 10075 26111 10081
rect 26605 10115 26663 10121
rect 26605 10081 26617 10115
rect 26651 10112 26663 10115
rect 26786 10112 26792 10124
rect 26651 10084 26792 10112
rect 26651 10081 26663 10084
rect 26605 10075 26663 10081
rect 26786 10072 26792 10084
rect 26844 10072 26850 10124
rect 26973 10115 27031 10121
rect 26973 10081 26985 10115
rect 27019 10081 27031 10115
rect 26973 10075 27031 10081
rect 26988 10044 27016 10075
rect 28626 10072 28632 10124
rect 28684 10072 28690 10124
rect 28810 10072 28816 10124
rect 28868 10112 28874 10124
rect 29089 10115 29147 10121
rect 29089 10112 29101 10115
rect 28868 10084 29101 10112
rect 28868 10072 28874 10084
rect 29089 10081 29101 10084
rect 29135 10081 29147 10115
rect 29089 10075 29147 10081
rect 30190 10072 30196 10124
rect 30248 10112 30254 10124
rect 30478 10115 30536 10121
rect 30478 10112 30490 10115
rect 30248 10084 30490 10112
rect 30248 10072 30254 10084
rect 30478 10081 30490 10084
rect 30524 10081 30536 10115
rect 30478 10075 30536 10081
rect 31018 10072 31024 10124
rect 31076 10072 31082 10124
rect 28902 10044 28908 10056
rect 26988 10016 28908 10044
rect 26326 9976 26332 9988
rect 25516 9948 26332 9976
rect 26326 9936 26332 9948
rect 26384 9936 26390 9988
rect 26513 9911 26571 9917
rect 26513 9908 26525 9911
rect 25188 9880 26525 9908
rect 25188 9868 25194 9880
rect 26513 9877 26525 9880
rect 26559 9877 26571 9911
rect 28736 9908 28764 10016
rect 28902 10004 28908 10016
rect 28960 10004 28966 10056
rect 30745 10047 30803 10053
rect 30745 10013 30757 10047
rect 30791 10044 30803 10047
rect 30929 10047 30987 10053
rect 30929 10044 30941 10047
rect 30791 10016 30941 10044
rect 30791 10013 30803 10016
rect 30745 10007 30803 10013
rect 30929 10013 30941 10016
rect 30975 10013 30987 10047
rect 30929 10007 30987 10013
rect 28813 9979 28871 9985
rect 28813 9945 28825 9979
rect 28859 9976 28871 9979
rect 28859 9948 29868 9976
rect 28859 9945 28871 9948
rect 28813 9939 28871 9945
rect 29365 9911 29423 9917
rect 29365 9908 29377 9911
rect 28736 9880 29377 9908
rect 26513 9871 26571 9877
rect 29365 9877 29377 9880
rect 29411 9877 29423 9911
rect 29840 9908 29868 9948
rect 30098 9908 30104 9920
rect 29840 9880 30104 9908
rect 29365 9871 29423 9877
rect 30098 9868 30104 9880
rect 30156 9868 30162 9920
rect 552 9818 31648 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 11436 9818
rect 11488 9766 11500 9818
rect 11552 9766 11564 9818
rect 11616 9766 11628 9818
rect 11680 9766 11692 9818
rect 11744 9766 19210 9818
rect 19262 9766 19274 9818
rect 19326 9766 19338 9818
rect 19390 9766 19402 9818
rect 19454 9766 19466 9818
rect 19518 9766 26984 9818
rect 27036 9766 27048 9818
rect 27100 9766 27112 9818
rect 27164 9766 27176 9818
rect 27228 9766 27240 9818
rect 27292 9766 31648 9818
rect 552 9744 31648 9766
rect 1578 9664 1584 9716
rect 1636 9664 1642 9716
rect 2038 9664 2044 9716
rect 2096 9704 2102 9716
rect 2096 9676 2774 9704
rect 2096 9664 2102 9676
rect 1213 9571 1271 9577
rect 1213 9537 1225 9571
rect 1259 9568 1271 9571
rect 2746 9568 2774 9676
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3740 9704 3746 9716
rect 3016 9676 3746 9704
rect 3016 9664 3022 9676
rect 3740 9664 3746 9676
rect 3798 9664 3804 9716
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 4430 9704 4436 9716
rect 4028 9676 4436 9704
rect 4028 9664 4034 9676
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 7190 9704 7196 9716
rect 4948 9676 7196 9704
rect 4948 9664 4954 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 9125 9707 9183 9713
rect 9125 9704 9137 9707
rect 8352 9676 9137 9704
rect 8352 9664 8358 9676
rect 9125 9673 9137 9676
rect 9171 9704 9183 9707
rect 10134 9704 10140 9716
rect 9171 9676 10140 9704
rect 9171 9673 9183 9676
rect 9125 9667 9183 9673
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 12342 9704 12348 9716
rect 11296 9676 12348 9704
rect 11296 9664 11302 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13541 9707 13599 9713
rect 13541 9704 13553 9707
rect 12768 9676 13553 9704
rect 12768 9664 12774 9676
rect 13541 9673 13553 9676
rect 13587 9673 13599 9707
rect 13541 9667 13599 9673
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15252 9676 15945 9704
rect 15252 9664 15258 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 21910 9704 21916 9716
rect 15933 9667 15991 9673
rect 20640 9676 21916 9704
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3510 9636 3516 9648
rect 3099 9608 3516 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3510 9596 3516 9608
rect 3568 9636 3574 9648
rect 5166 9636 5172 9648
rect 3568 9608 5172 9636
rect 3568 9596 3574 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 5534 9636 5540 9648
rect 5276 9608 5540 9636
rect 4890 9568 4896 9580
rect 1259 9540 1808 9568
rect 2746 9540 4896 9568
rect 1259 9537 1271 9540
rect 1213 9531 1271 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 1412 9432 1440 9463
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 1780 9500 1808 9540
rect 4890 9528 4896 9540
rect 4948 9568 4954 9580
rect 5276 9568 5304 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 9033 9639 9091 9645
rect 8904 9608 8984 9636
rect 8904 9596 8910 9608
rect 4948 9540 5304 9568
rect 4948 9528 4954 9540
rect 2866 9500 2872 9512
rect 1780 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3234 9460 3240 9512
rect 3292 9460 3298 9512
rect 3694 9460 3700 9512
rect 3752 9460 3758 9512
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3927 9472 4169 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4157 9463 4215 9469
rect 4338 9460 4344 9512
rect 4396 9460 4402 9512
rect 5276 9509 5304 9540
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7742 9568 7748 9580
rect 7064 9540 7748 9568
rect 7064 9528 7070 9540
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 8956 9568 8984 9608
rect 9033 9605 9045 9639
rect 9079 9636 9091 9639
rect 9674 9636 9680 9648
rect 9079 9608 9680 9636
rect 9079 9605 9091 9608
rect 9033 9599 9091 9605
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 16666 9636 16672 9648
rect 16592 9608 16672 9636
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 8628 9540 8892 9568
rect 8956 9540 9229 9568
rect 8628 9528 8634 9540
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5399 9472 5549 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 1940 9435 1998 9441
rect 1412 9404 1900 9432
rect 1872 9364 1900 9404
rect 1940 9401 1952 9435
rect 1986 9432 1998 9435
rect 2314 9432 2320 9444
rect 1986 9404 2320 9432
rect 1986 9401 1998 9404
rect 1940 9395 1998 9401
rect 2314 9392 2320 9404
rect 2372 9392 2378 9444
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 3375 9435 3433 9441
rect 3375 9432 3387 9435
rect 3200 9404 3387 9432
rect 3200 9392 3206 9404
rect 3375 9401 3387 9404
rect 3421 9401 3433 9435
rect 3375 9395 3433 9401
rect 3510 9392 3516 9444
rect 3568 9392 3574 9444
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 4246 9432 4252 9444
rect 3651 9404 4252 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 4246 9392 4252 9404
rect 4304 9392 4310 9444
rect 5804 9435 5862 9441
rect 5804 9401 5816 9435
rect 5850 9432 5862 9435
rect 7006 9432 7012 9444
rect 5850 9404 7012 9432
rect 5850 9401 5862 9404
rect 5804 9395 5862 9401
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 2958 9364 2964 9376
rect 1872 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 3973 9367 4031 9373
rect 3973 9364 3985 9367
rect 3292 9336 3985 9364
rect 3292 9324 3298 9336
rect 3973 9333 3985 9336
rect 4019 9333 4031 9367
rect 3973 9327 4031 9333
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6420 9336 6929 9364
rect 6420 9324 6426 9336
rect 6917 9333 6929 9336
rect 6963 9364 6975 9367
rect 7208 9364 7236 9463
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 8864 9509 8892 9540
rect 9217 9537 9229 9540
rect 9263 9537 9275 9571
rect 14274 9568 14280 9580
rect 9217 9531 9275 9537
rect 13464 9540 14280 9568
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9306 9500 9312 9512
rect 9180 9472 9312 9500
rect 9180 9460 9186 9472
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 9398 9460 9404 9512
rect 9456 9460 9462 9512
rect 10226 9460 10232 9512
rect 10284 9460 10290 9512
rect 10778 9509 10784 9512
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9500 10379 9503
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 10367 9472 10517 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10772 9500 10784 9509
rect 10739 9472 10784 9500
rect 10505 9463 10563 9469
rect 10772 9463 10784 9472
rect 10778 9460 10784 9463
rect 10836 9460 10842 9512
rect 11974 9460 11980 9512
rect 12032 9460 12038 9512
rect 12066 9460 12072 9512
rect 12124 9500 12130 9512
rect 12233 9503 12291 9509
rect 12233 9500 12245 9503
rect 12124 9472 12245 9500
rect 12124 9460 12130 9472
rect 12233 9469 12245 9472
rect 12279 9469 12291 9503
rect 13464 9500 13492 9540
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 16592 9577 16620 9608
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 20640 9636 20668 9676
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 25130 9664 25136 9716
rect 25188 9664 25194 9716
rect 25593 9707 25651 9713
rect 25593 9673 25605 9707
rect 25639 9704 25651 9707
rect 25774 9704 25780 9716
rect 25639 9676 25780 9704
rect 25639 9673 25651 9676
rect 25593 9667 25651 9673
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 26694 9704 26700 9716
rect 25884 9676 26700 9704
rect 19904 9608 20668 9636
rect 16577 9571 16635 9577
rect 16577 9537 16589 9571
rect 16623 9537 16635 9571
rect 16577 9531 16635 9537
rect 16776 9540 17264 9568
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 12233 9463 12291 9469
rect 12406 9472 13492 9500
rect 13556 9472 14105 9500
rect 8478 9392 8484 9444
rect 8536 9441 8542 9444
rect 8536 9435 8585 9441
rect 8536 9401 8539 9435
rect 8573 9401 8585 9435
rect 8536 9395 8585 9401
rect 8665 9435 8723 9441
rect 8665 9401 8677 9435
rect 8711 9432 8723 9435
rect 8938 9432 8944 9444
rect 8711 9404 8944 9432
rect 8711 9401 8723 9404
rect 8665 9395 8723 9401
rect 8536 9392 8542 9395
rect 8938 9392 8944 9404
rect 8996 9392 9002 9444
rect 11790 9432 11796 9444
rect 9508 9404 11796 9432
rect 6963 9336 7236 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 7834 9324 7840 9376
rect 7892 9324 7898 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 9508 9364 9536 9404
rect 11790 9392 11796 9404
rect 11848 9432 11854 9444
rect 12406 9432 12434 9472
rect 11848 9404 12434 9432
rect 11848 9392 11854 9404
rect 13556 9376 13584 9472
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 16114 9460 16120 9512
rect 16172 9460 16178 9512
rect 16206 9460 16212 9512
rect 16264 9460 16270 9512
rect 16776 9509 16804 9540
rect 16761 9503 16819 9509
rect 16761 9469 16773 9503
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17126 9460 17132 9512
rect 17184 9460 17190 9512
rect 17236 9500 17264 9540
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 19904 9568 19932 9608
rect 23474 9596 23480 9648
rect 23532 9596 23538 9648
rect 25685 9639 25743 9645
rect 25685 9636 25697 9639
rect 23584 9608 25697 9636
rect 18472 9540 19932 9568
rect 18472 9528 18478 9540
rect 18690 9500 18696 9512
rect 17236 9472 18696 9500
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 18874 9460 18880 9512
rect 18932 9460 18938 9512
rect 19904 9509 19932 9540
rect 20180 9540 20760 9568
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 20070 9460 20076 9512
rect 20128 9460 20134 9512
rect 20180 9509 20208 9540
rect 20165 9503 20223 9509
rect 20165 9469 20177 9503
rect 20211 9469 20223 9503
rect 20165 9463 20223 9469
rect 20257 9503 20315 9509
rect 20257 9469 20269 9503
rect 20303 9500 20315 9503
rect 20346 9500 20352 9512
rect 20303 9472 20352 9500
rect 20303 9469 20315 9472
rect 20257 9463 20315 9469
rect 14366 9392 14372 9444
rect 14424 9432 14430 9444
rect 14706 9435 14764 9441
rect 14706 9432 14718 9435
rect 14424 9404 14718 9432
rect 14424 9392 14430 9404
rect 14706 9401 14718 9404
rect 14752 9401 14764 9435
rect 14706 9395 14764 9401
rect 15930 9392 15936 9444
rect 15988 9432 15994 9444
rect 16301 9435 16359 9441
rect 16301 9432 16313 9435
rect 15988 9404 16313 9432
rect 15988 9392 15994 9404
rect 16301 9401 16313 9404
rect 16347 9401 16359 9435
rect 16301 9395 16359 9401
rect 16390 9392 16396 9444
rect 16448 9441 16454 9444
rect 16448 9435 16477 9441
rect 16465 9401 16477 9435
rect 16448 9395 16477 9401
rect 17037 9435 17095 9441
rect 17037 9401 17049 9435
rect 17083 9432 17095 9435
rect 17374 9435 17432 9441
rect 17374 9432 17386 9435
rect 17083 9404 17386 9432
rect 17083 9401 17095 9404
rect 17037 9395 17095 9401
rect 17374 9401 17386 9404
rect 17420 9401 17432 9435
rect 17374 9395 17432 9401
rect 16448 9392 16454 9395
rect 17494 9392 17500 9444
rect 17552 9432 17558 9444
rect 20272 9432 20300 9463
rect 20346 9460 20352 9472
rect 20404 9460 20410 9512
rect 20622 9460 20628 9512
rect 20680 9460 20686 9512
rect 20732 9500 20760 9540
rect 22094 9528 22100 9580
rect 22152 9528 22158 9580
rect 23106 9528 23112 9580
rect 23164 9568 23170 9580
rect 23584 9568 23612 9608
rect 25685 9605 25697 9608
rect 25731 9636 25743 9639
rect 25884 9636 25912 9676
rect 26694 9664 26700 9676
rect 26752 9664 26758 9716
rect 27433 9707 27491 9713
rect 27433 9673 27445 9707
rect 27479 9704 27491 9707
rect 28166 9704 28172 9716
rect 27479 9676 28172 9704
rect 27479 9673 27491 9676
rect 27433 9667 27491 9673
rect 28166 9664 28172 9676
rect 28224 9704 28230 9716
rect 28629 9707 28687 9713
rect 28629 9704 28641 9707
rect 28224 9676 28641 9704
rect 28224 9664 28230 9676
rect 28629 9673 28641 9676
rect 28675 9673 28687 9707
rect 28629 9667 28687 9673
rect 25731 9608 25912 9636
rect 25731 9605 25743 9608
rect 25685 9599 25743 9605
rect 25958 9596 25964 9648
rect 26016 9636 26022 9648
rect 26602 9636 26608 9648
rect 26016 9608 26608 9636
rect 26016 9596 26022 9608
rect 26602 9596 26608 9608
rect 26660 9596 26666 9648
rect 26878 9596 26884 9648
rect 26936 9636 26942 9648
rect 26973 9639 27031 9645
rect 26973 9636 26985 9639
rect 26936 9608 26985 9636
rect 26936 9596 26942 9608
rect 26973 9605 26985 9608
rect 27019 9605 27031 9639
rect 26973 9599 27031 9605
rect 27062 9596 27068 9648
rect 27120 9636 27126 9648
rect 28074 9636 28080 9648
rect 27120 9608 28080 9636
rect 27120 9596 27126 9608
rect 28074 9596 28080 9608
rect 28132 9596 28138 9648
rect 28353 9639 28411 9645
rect 28353 9605 28365 9639
rect 28399 9636 28411 9639
rect 28994 9636 29000 9648
rect 28399 9608 29000 9636
rect 28399 9605 28411 9608
rect 28353 9599 28411 9605
rect 28994 9596 29000 9608
rect 29052 9596 29058 9648
rect 23164 9540 23612 9568
rect 24136 9540 26255 9568
rect 23164 9528 23170 9540
rect 22002 9500 22008 9512
rect 20732 9472 22008 9500
rect 22002 9460 22008 9472
rect 22060 9460 22066 9512
rect 24136 9500 24164 9540
rect 22296 9472 24164 9500
rect 24213 9503 24271 9509
rect 17552 9404 20300 9432
rect 20533 9435 20591 9441
rect 17552 9392 17558 9404
rect 20533 9401 20545 9435
rect 20579 9432 20591 9435
rect 20870 9435 20928 9441
rect 20870 9432 20882 9435
rect 20579 9404 20882 9432
rect 20579 9401 20591 9404
rect 20533 9395 20591 9401
rect 20870 9401 20882 9404
rect 20916 9401 20928 9435
rect 20870 9395 20928 9401
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 22296 9432 22324 9472
rect 24213 9469 24225 9503
rect 24259 9469 24271 9503
rect 24213 9463 24271 9469
rect 24367 9503 24425 9509
rect 24367 9469 24379 9503
rect 24413 9500 24425 9503
rect 24854 9500 24860 9512
rect 24413 9472 24860 9500
rect 24413 9469 24425 9472
rect 24367 9463 24425 9469
rect 21140 9404 22324 9432
rect 22364 9435 22422 9441
rect 21140 9392 21146 9404
rect 22364 9401 22376 9435
rect 22410 9432 22422 9435
rect 22462 9432 22468 9444
rect 22410 9404 22468 9432
rect 22410 9401 22422 9404
rect 22364 9395 22422 9401
rect 22462 9392 22468 9404
rect 22520 9392 22526 9444
rect 24228 9432 24256 9463
rect 24854 9460 24860 9472
rect 24912 9500 24918 9512
rect 24912 9472 24992 9500
rect 24912 9460 24918 9472
rect 24486 9432 24492 9444
rect 24228 9404 24492 9432
rect 24486 9392 24492 9404
rect 24544 9392 24550 9444
rect 24964 9432 24992 9472
rect 25038 9460 25044 9512
rect 25096 9460 25102 9512
rect 25222 9460 25228 9512
rect 25280 9500 25286 9512
rect 25317 9503 25375 9509
rect 25317 9500 25329 9503
rect 25280 9472 25329 9500
rect 25280 9460 25286 9472
rect 25317 9469 25329 9472
rect 25363 9469 25375 9503
rect 25317 9463 25375 9469
rect 25406 9460 25412 9512
rect 25464 9460 25470 9512
rect 26068 9509 26096 9540
rect 26053 9503 26111 9509
rect 26053 9469 26065 9503
rect 26099 9469 26111 9503
rect 26227 9500 26255 9540
rect 26326 9528 26332 9580
rect 26384 9568 26390 9580
rect 26789 9571 26847 9577
rect 26789 9568 26801 9571
rect 26384 9540 26801 9568
rect 26384 9528 26390 9540
rect 26789 9537 26801 9540
rect 26835 9568 26847 9571
rect 27249 9571 27307 9577
rect 27249 9568 27261 9571
rect 26835 9540 27261 9568
rect 26835 9537 26847 9540
rect 26789 9531 26847 9537
rect 27249 9537 27261 9540
rect 27295 9537 27307 9571
rect 27249 9531 27307 9537
rect 27338 9528 27344 9580
rect 27396 9568 27402 9580
rect 27396 9540 29224 9568
rect 27396 9528 27402 9540
rect 26513 9503 26571 9509
rect 26513 9500 26525 9503
rect 26227 9472 26525 9500
rect 26053 9463 26111 9469
rect 26513 9469 26525 9472
rect 26559 9469 26571 9503
rect 26513 9463 26571 9469
rect 26602 9460 26608 9512
rect 26660 9460 26666 9512
rect 26694 9460 26700 9512
rect 26752 9460 26758 9512
rect 26878 9460 26884 9512
rect 26936 9500 26942 9512
rect 27157 9503 27215 9509
rect 27157 9500 27169 9503
rect 26936 9472 27169 9500
rect 26936 9460 26942 9472
rect 27157 9469 27169 9472
rect 27203 9500 27215 9503
rect 27203 9472 28028 9500
rect 27203 9469 27215 9472
rect 27157 9463 27215 9469
rect 25869 9435 25927 9441
rect 25869 9432 25881 9435
rect 24964 9404 25881 9432
rect 25869 9401 25881 9404
rect 25915 9432 25927 9435
rect 26142 9432 26148 9444
rect 25915 9404 26148 9432
rect 25915 9401 25927 9404
rect 25869 9395 25927 9401
rect 26142 9392 26148 9404
rect 26200 9392 26206 9444
rect 26234 9392 26240 9444
rect 26292 9432 26298 9444
rect 27062 9432 27068 9444
rect 26292 9404 27068 9432
rect 26292 9392 26298 9404
rect 27062 9392 27068 9404
rect 27120 9392 27126 9444
rect 27433 9435 27491 9441
rect 27433 9432 27445 9435
rect 27264 9404 27445 9432
rect 8444 9336 9536 9364
rect 9585 9367 9643 9373
rect 8444 9324 8450 9336
rect 9585 9333 9597 9367
rect 9631 9364 9643 9367
rect 10042 9364 10048 9376
rect 9631 9336 10048 9364
rect 9631 9333 9643 9336
rect 9585 9327 9643 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11664 9336 11897 9364
rect 11664 9324 11670 9336
rect 11885 9333 11897 9336
rect 11931 9333 11943 9367
rect 11885 9327 11943 9333
rect 13357 9367 13415 9373
rect 13357 9333 13369 9367
rect 13403 9364 13415 9367
rect 13538 9364 13544 9376
rect 13403 9336 13544 9364
rect 13403 9333 13415 9336
rect 13357 9327 13415 9333
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 15838 9364 15844 9376
rect 14884 9336 15844 9364
rect 14884 9324 14890 9336
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18012 9336 18521 9364
rect 18012 9324 18018 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 18782 9324 18788 9376
rect 18840 9324 18846 9376
rect 20070 9324 20076 9376
rect 20128 9364 20134 9376
rect 21266 9364 21272 9376
rect 20128 9336 21272 9364
rect 20128 9324 20134 9336
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 22005 9367 22063 9373
rect 22005 9333 22017 9367
rect 22051 9364 22063 9367
rect 22278 9364 22284 9376
rect 22051 9336 22284 9364
rect 22051 9333 22063 9336
rect 22005 9327 22063 9333
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 24581 9367 24639 9373
rect 24581 9333 24593 9367
rect 24627 9364 24639 9367
rect 24946 9364 24952 9376
rect 24627 9336 24952 9364
rect 24627 9333 24639 9336
rect 24581 9327 24639 9333
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 25958 9324 25964 9376
rect 26016 9324 26022 9376
rect 26329 9367 26387 9373
rect 26329 9333 26341 9367
rect 26375 9364 26387 9367
rect 26418 9364 26424 9376
rect 26375 9336 26424 9364
rect 26375 9333 26387 9336
rect 26329 9327 26387 9333
rect 26418 9324 26424 9336
rect 26476 9324 26482 9376
rect 26602 9324 26608 9376
rect 26660 9364 26666 9376
rect 27264 9364 27292 9404
rect 27433 9401 27445 9404
rect 27479 9401 27491 9435
rect 28000 9432 28028 9472
rect 28074 9460 28080 9512
rect 28132 9460 28138 9512
rect 28166 9460 28172 9512
rect 28224 9460 28230 9512
rect 29196 9509 29224 9540
rect 30190 9528 30196 9580
rect 30248 9528 30254 9580
rect 28353 9503 28411 9509
rect 28353 9469 28365 9503
rect 28399 9500 28411 9503
rect 29181 9503 29239 9509
rect 28399 9472 28856 9500
rect 28399 9469 28411 9472
rect 28353 9463 28411 9469
rect 28442 9432 28448 9444
rect 28000 9404 28448 9432
rect 27433 9395 27491 9401
rect 28442 9392 28448 9404
rect 28500 9392 28506 9444
rect 28828 9432 28856 9472
rect 29181 9469 29193 9503
rect 29227 9469 29239 9503
rect 29181 9463 29239 9469
rect 29914 9460 29920 9512
rect 29972 9460 29978 9512
rect 30098 9460 30104 9512
rect 30156 9460 30162 9512
rect 30282 9460 30288 9512
rect 30340 9460 30346 9512
rect 29365 9435 29423 9441
rect 29365 9432 29377 9435
rect 28828 9404 29377 9432
rect 29365 9401 29377 9404
rect 29411 9401 29423 9435
rect 29365 9395 29423 9401
rect 26660 9336 27292 9364
rect 26660 9324 26666 9336
rect 28074 9324 28080 9376
rect 28132 9364 28138 9376
rect 28645 9367 28703 9373
rect 28645 9364 28657 9367
rect 28132 9336 28657 9364
rect 28132 9324 28138 9336
rect 28645 9333 28657 9336
rect 28691 9333 28703 9367
rect 28645 9327 28703 9333
rect 28810 9324 28816 9376
rect 28868 9324 28874 9376
rect 29086 9324 29092 9376
rect 29144 9324 29150 9376
rect 552 9274 31648 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 12096 9274
rect 12148 9222 12160 9274
rect 12212 9222 12224 9274
rect 12276 9222 12288 9274
rect 12340 9222 12352 9274
rect 12404 9222 19870 9274
rect 19922 9222 19934 9274
rect 19986 9222 19998 9274
rect 20050 9222 20062 9274
rect 20114 9222 20126 9274
rect 20178 9222 27644 9274
rect 27696 9222 27708 9274
rect 27760 9222 27772 9274
rect 27824 9222 27836 9274
rect 27888 9222 27900 9274
rect 27952 9222 31648 9274
rect 552 9200 31648 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1857 9163 1915 9169
rect 1857 9160 1869 9163
rect 1728 9132 1869 9160
rect 1728 9120 1734 9132
rect 1857 9129 1869 9132
rect 1903 9129 1915 9163
rect 1857 9123 1915 9129
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3513 9163 3571 9169
rect 3513 9160 3525 9163
rect 3016 9132 3525 9160
rect 3016 9120 3022 9132
rect 3513 9129 3525 9132
rect 3559 9129 3571 9163
rect 6822 9160 6828 9172
rect 3513 9123 3571 9129
rect 4816 9132 6828 9160
rect 2038 9052 2044 9104
rect 2096 9052 2102 9104
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 3326 9092 3332 9104
rect 3108 9064 3332 9092
rect 3108 9052 3114 9064
rect 3326 9052 3332 9064
rect 3384 9092 3390 9104
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 3384 9064 3801 9092
rect 3384 9052 3390 9064
rect 3789 9061 3801 9064
rect 3835 9061 3847 9095
rect 3789 9055 3847 9061
rect 3970 9052 3976 9104
rect 4028 9101 4034 9104
rect 4028 9095 4077 9101
rect 4028 9061 4031 9095
rect 4065 9092 4077 9095
rect 4816 9092 4844 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7006 9120 7012 9172
rect 7064 9120 7070 9172
rect 7834 9160 7840 9172
rect 7300 9132 7840 9160
rect 4065 9064 4844 9092
rect 4065 9061 4077 9064
rect 4028 9055 4077 9061
rect 4028 9052 4034 9055
rect 4890 9052 4896 9104
rect 4948 9052 4954 9104
rect 7300 9092 7328 9132
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 10505 9163 10563 9169
rect 9539 9132 10180 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 7558 9101 7564 9104
rect 7377 9095 7435 9101
rect 7377 9092 7389 9095
rect 7300 9064 7389 9092
rect 7377 9061 7389 9064
rect 7423 9061 7435 9095
rect 7377 9055 7435 9061
rect 7515 9095 7564 9101
rect 7515 9061 7527 9095
rect 7561 9061 7564 9095
rect 7515 9055 7564 9061
rect 7558 9052 7564 9055
rect 7616 9052 7622 9104
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2056 9024 2084 9052
rect 1995 8996 2084 9024
rect 2308 9027 2366 9033
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2308 8993 2320 9027
rect 2354 9024 2366 9027
rect 3234 9024 3240 9036
rect 2354 8996 3240 9024
rect 2354 8993 2366 8996
rect 2308 8987 2366 8993
rect 3234 8984 3240 8996
rect 3292 8984 3298 9036
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 3694 9024 3700 9036
rect 3568 8996 3700 9024
rect 3568 8984 3574 8996
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1820 8928 2053 8956
rect 1820 8916 1826 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 3602 8956 3608 8968
rect 3384 8928 3608 8956
rect 3384 8916 3390 8928
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 3896 8888 3924 8987
rect 4154 8984 4160 9036
rect 4212 8984 4218 9036
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 5675 8996 6745 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5040 8928 5917 8956
rect 5040 8916 5046 8928
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 4614 8888 4620 8900
rect 3896 8860 4620 8888
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 4246 8820 4252 8832
rect 3467 8792 4252 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 4246 8780 4252 8792
rect 4304 8820 4310 8832
rect 4706 8820 4712 8832
rect 4304 8792 4712 8820
rect 4304 8780 4310 8792
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 6748 8820 6776 8987
rect 7208 8888 7236 8987
rect 7282 8984 7288 9036
rect 7340 8984 7346 9036
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 9024 7711 9027
rect 7742 9024 7748 9036
rect 7699 8996 7748 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 9306 8984 9312 9036
rect 9364 8984 9370 9036
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 9024 9551 9027
rect 9674 9024 9680 9036
rect 9539 8996 9680 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9769 9027 9827 9033
rect 9769 8993 9781 9027
rect 9815 9024 9827 9027
rect 9815 8996 9904 9024
rect 9815 8993 9827 8996
rect 9769 8987 9827 8993
rect 8662 8888 8668 8900
rect 7208 8860 8668 8888
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 9766 8820 9772 8832
rect 6748 8792 9772 8820
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 9876 8820 9904 8996
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10152 9033 10180 9132
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 11054 9160 11060 9172
rect 10551 9132 11060 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 12032 9132 12173 9160
rect 12032 9120 12038 9132
rect 12161 9129 12173 9132
rect 12207 9129 12219 9163
rect 13078 9160 13084 9172
rect 12161 9123 12219 9129
rect 12268 9132 13084 9160
rect 11606 9092 11612 9104
rect 11440 9064 11612 9092
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 9950 8916 9956 8968
rect 10008 8916 10014 8968
rect 10244 8888 10272 8987
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11440 9024 11468 9064
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 11882 9101 11888 9104
rect 11839 9095 11888 9101
rect 11839 9061 11851 9095
rect 11885 9061 11888 9095
rect 11839 9055 11888 9061
rect 11882 9052 11888 9055
rect 11940 9052 11946 9104
rect 12268 9092 12296 9132
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 13817 9163 13875 9169
rect 13817 9129 13829 9163
rect 13863 9160 13875 9163
rect 14458 9160 14464 9172
rect 13863 9132 14464 9160
rect 13863 9129 13875 9132
rect 13817 9123 13875 9129
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 15381 9163 15439 9169
rect 15381 9160 15393 9163
rect 14752 9132 15393 9160
rect 11992 9064 12296 9092
rect 11296 8996 11468 9024
rect 11517 9027 11575 9033
rect 11296 8984 11302 8996
rect 11517 8993 11529 9027
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 11204 8928 11345 8956
rect 11204 8916 11210 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11532 8956 11560 8987
rect 11698 8984 11704 9036
rect 11756 8984 11762 9036
rect 11992 9033 12020 9064
rect 14366 9052 14372 9104
rect 14424 9052 14430 9104
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 12253 9027 12311 9033
rect 12253 9024 12265 9027
rect 12124 8996 12265 9024
rect 12124 8984 12130 8996
rect 12253 8993 12265 8996
rect 12299 9024 12311 9027
rect 13722 9024 13728 9036
rect 12299 8996 13728 9024
rect 12299 8993 12311 8996
rect 12253 8987 12311 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 14185 9027 14243 9033
rect 13823 8996 14136 9024
rect 12526 8956 12532 8968
rect 11532 8928 12532 8956
rect 11333 8919 11391 8925
rect 12526 8916 12532 8928
rect 12584 8956 12590 8968
rect 13823 8956 13851 8996
rect 12584 8928 13851 8956
rect 14001 8959 14059 8965
rect 12584 8916 12590 8928
rect 14001 8925 14013 8959
rect 14047 8925 14059 8959
rect 14108 8956 14136 8996
rect 14185 8993 14197 9027
rect 14231 9024 14243 9027
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 14231 8996 14565 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 14553 8987 14611 8993
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 14752 9033 14780 9132
rect 15381 9129 15393 9132
rect 15427 9160 15439 9163
rect 16114 9160 16120 9172
rect 15427 9132 16120 9160
rect 15427 9129 15439 9132
rect 15381 9123 15439 9129
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17313 9163 17371 9169
rect 17313 9160 17325 9163
rect 17184 9132 17325 9160
rect 17184 9120 17190 9132
rect 17313 9129 17325 9132
rect 17359 9129 17371 9163
rect 18874 9160 18880 9172
rect 17313 9123 17371 9129
rect 17420 9132 18880 9160
rect 14826 9052 14832 9104
rect 14884 9052 14890 9104
rect 15059 9095 15117 9101
rect 15059 9061 15071 9095
rect 15105 9092 15117 9095
rect 16390 9092 16396 9104
rect 15105 9064 16396 9092
rect 15105 9061 15117 9064
rect 15059 9055 15117 9061
rect 15580 9036 15608 9064
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14700 8996 14749 9024
rect 14700 8984 14706 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 14660 8956 14688 8984
rect 14108 8928 14688 8956
rect 14936 8956 14964 8987
rect 15194 8984 15200 9036
rect 15252 8984 15258 9036
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 9024 15439 9027
rect 15470 9024 15476 9036
rect 15427 8996 15476 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 15562 8984 15568 9036
rect 15620 8984 15626 9036
rect 17420 9033 17448 9132
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 20622 9120 20628 9172
rect 20680 9160 20686 9172
rect 20809 9163 20867 9169
rect 20809 9160 20821 9163
rect 20680 9132 20821 9160
rect 20680 9120 20686 9132
rect 20809 9129 20821 9132
rect 20855 9129 20867 9163
rect 20809 9123 20867 9129
rect 21266 9120 21272 9172
rect 21324 9120 21330 9172
rect 22370 9160 22376 9172
rect 21836 9132 22376 9160
rect 18782 9092 18788 9104
rect 17972 9064 18788 9092
rect 17972 9033 18000 9064
rect 18782 9052 18788 9064
rect 18840 9052 18846 9104
rect 20346 9052 20352 9104
rect 20404 9092 20410 9104
rect 21082 9092 21088 9104
rect 20404 9064 21088 9092
rect 20404 9052 20410 9064
rect 21082 9052 21088 9064
rect 21140 9052 21146 9104
rect 21453 9095 21511 9101
rect 21453 9061 21465 9095
rect 21499 9092 21511 9095
rect 21729 9095 21787 9101
rect 21729 9092 21741 9095
rect 21499 9064 21741 9092
rect 21499 9061 21511 9064
rect 21453 9055 21511 9061
rect 21729 9061 21741 9064
rect 21775 9061 21787 9095
rect 21729 9055 21787 9061
rect 18230 9033 18236 9036
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 8993 17463 9027
rect 17405 8987 17463 8993
rect 17957 9027 18015 9033
rect 17957 8993 17969 9027
rect 18003 8993 18015 9027
rect 17957 8987 18015 8993
rect 18224 8987 18236 9033
rect 18230 8984 18236 8987
rect 18288 8984 18294 9036
rect 20438 8984 20444 9036
rect 20496 9024 20502 9036
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 20496 8996 20913 9024
rect 20496 8984 20502 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 21637 9027 21695 9033
rect 21637 8993 21649 9027
rect 21683 9024 21695 9027
rect 21836 9024 21864 9132
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 22462 9120 22468 9172
rect 22520 9120 22526 9172
rect 25317 9163 25375 9169
rect 23492 9132 25268 9160
rect 21910 9052 21916 9104
rect 21968 9092 21974 9104
rect 21968 9064 23152 9092
rect 21968 9052 21974 9064
rect 21683 8996 21864 9024
rect 21683 8993 21695 8996
rect 21637 8987 21695 8993
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 22741 9027 22799 9033
rect 22741 9024 22753 9027
rect 22152 8996 22753 9024
rect 22152 8984 22158 8996
rect 22741 8993 22753 8996
rect 22787 8993 22799 9027
rect 22741 8987 22799 8993
rect 22830 8984 22836 9036
rect 22888 8984 22894 9036
rect 22922 8984 22928 9036
rect 22980 8984 22986 9036
rect 23124 9033 23152 9064
rect 23109 9027 23167 9033
rect 23109 8993 23121 9027
rect 23155 8993 23167 9027
rect 23109 8987 23167 8993
rect 23201 9027 23259 9033
rect 23201 8993 23213 9027
rect 23247 8993 23259 9027
rect 23201 8987 23259 8993
rect 23294 9027 23352 9033
rect 23294 8993 23306 9027
rect 23340 9024 23352 9027
rect 23492 9024 23520 9132
rect 23569 9095 23627 9101
rect 23569 9061 23581 9095
rect 23615 9092 23627 9095
rect 23615 9064 24808 9092
rect 23615 9061 23627 9064
rect 23569 9055 23627 9061
rect 23340 8996 23520 9024
rect 23340 8993 23352 8996
rect 23294 8987 23352 8993
rect 15930 8956 15936 8968
rect 14936 8928 15936 8956
rect 14001 8919 14059 8925
rect 12710 8888 12716 8900
rect 10244 8860 12716 8888
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 14016 8888 14044 8919
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 22278 8916 22284 8968
rect 22336 8956 22342 8968
rect 22373 8959 22431 8965
rect 22373 8956 22385 8959
rect 22336 8928 22385 8956
rect 22336 8916 22342 8928
rect 22373 8925 22385 8928
rect 22419 8956 22431 8959
rect 23216 8956 23244 8987
rect 22419 8928 23244 8956
rect 22419 8925 22431 8928
rect 22373 8919 22431 8925
rect 15378 8888 15384 8900
rect 14016 8860 15384 8888
rect 15378 8848 15384 8860
rect 15436 8888 15442 8900
rect 16022 8888 16028 8900
rect 15436 8860 16028 8888
rect 15436 8848 15442 8860
rect 16022 8848 16028 8860
rect 16080 8848 16086 8900
rect 22002 8848 22008 8900
rect 22060 8888 22066 8900
rect 22830 8888 22836 8900
rect 22060 8860 22836 8888
rect 22060 8848 22066 8860
rect 22830 8848 22836 8860
rect 22888 8848 22894 8900
rect 10594 8820 10600 8832
rect 9876 8792 10600 8820
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11698 8820 11704 8832
rect 11204 8792 11704 8820
rect 11204 8780 11210 8792
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 18138 8820 18144 8832
rect 15528 8792 18144 8820
rect 15528 8780 15534 8792
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19337 8823 19395 8829
rect 19337 8820 19349 8823
rect 19024 8792 19349 8820
rect 19024 8780 19030 8792
rect 19337 8789 19349 8792
rect 19383 8789 19395 8823
rect 19337 8783 19395 8789
rect 20254 8780 20260 8832
rect 20312 8820 20318 8832
rect 23308 8820 23336 8987
rect 24486 8984 24492 9036
rect 24544 9024 24550 9036
rect 24780 9033 24808 9064
rect 24946 9052 24952 9104
rect 25004 9052 25010 9104
rect 25240 9092 25268 9132
rect 25317 9129 25329 9163
rect 25363 9160 25375 9163
rect 25866 9160 25872 9172
rect 25363 9132 25872 9160
rect 25363 9129 25375 9132
rect 25317 9123 25375 9129
rect 25866 9120 25872 9132
rect 25924 9120 25930 9172
rect 26694 9160 26700 9172
rect 26436 9132 26700 9160
rect 25958 9092 25964 9104
rect 25240 9064 25964 9092
rect 25958 9052 25964 9064
rect 26016 9052 26022 9104
rect 26234 9052 26240 9104
rect 26292 9052 26298 9104
rect 26436 9101 26464 9132
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 28442 9120 28448 9172
rect 28500 9160 28506 9172
rect 28905 9163 28963 9169
rect 28905 9160 28917 9163
rect 28500 9132 28917 9160
rect 28500 9120 28506 9132
rect 28905 9129 28917 9132
rect 28951 9160 28963 9163
rect 29914 9160 29920 9172
rect 28951 9132 29920 9160
rect 28951 9129 28963 9132
rect 28905 9123 28963 9129
rect 29914 9120 29920 9132
rect 29972 9120 29978 9172
rect 26421 9095 26479 9101
rect 26421 9061 26433 9095
rect 26467 9061 26479 9095
rect 26421 9055 26479 9061
rect 26510 9052 26516 9104
rect 26568 9092 26574 9104
rect 26605 9095 26663 9101
rect 26605 9092 26617 9095
rect 26568 9064 26617 9092
rect 26568 9052 26574 9064
rect 26605 9061 26617 9064
rect 26651 9061 26663 9095
rect 26605 9055 26663 9061
rect 29086 9052 29092 9104
rect 29144 9092 29150 9104
rect 29144 9064 30328 9092
rect 29144 9052 29150 9064
rect 24673 9027 24731 9033
rect 24673 9024 24685 9027
rect 24544 8996 24685 9024
rect 24544 8984 24550 8996
rect 24673 8993 24685 8996
rect 24719 8993 24731 9027
rect 24673 8987 24731 8993
rect 24766 9027 24824 9033
rect 24766 8993 24778 9027
rect 24812 8993 24824 9027
rect 24766 8987 24824 8993
rect 25041 9027 25099 9033
rect 25041 8993 25053 9027
rect 25087 8993 25099 9027
rect 25041 8987 25099 8993
rect 25179 9027 25237 9033
rect 25179 8993 25191 9027
rect 25225 9024 25237 9027
rect 25406 9024 25412 9036
rect 25225 8996 25412 9024
rect 25225 8993 25237 8996
rect 25179 8987 25237 8993
rect 24397 8959 24455 8965
rect 24397 8925 24409 8959
rect 24443 8956 24455 8959
rect 24578 8956 24584 8968
rect 24443 8928 24584 8956
rect 24443 8925 24455 8928
rect 24397 8919 24455 8925
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 25056 8956 25084 8987
rect 25406 8984 25412 8996
rect 25464 8984 25470 9036
rect 25501 9027 25559 9033
rect 25501 8993 25513 9027
rect 25547 9024 25559 9027
rect 26326 9024 26332 9036
rect 25547 8996 26332 9024
rect 25547 8993 25559 8996
rect 25501 8987 25559 8993
rect 26326 8984 26332 8996
rect 26384 8984 26390 9036
rect 26973 9027 27031 9033
rect 26973 8993 26985 9027
rect 27019 9024 27031 9027
rect 27893 9027 27951 9033
rect 27893 9024 27905 9027
rect 27019 8996 27905 9024
rect 27019 8993 27031 8996
rect 26973 8987 27031 8993
rect 27893 8993 27905 8996
rect 27939 8993 27951 9027
rect 27893 8987 27951 8993
rect 28166 8984 28172 9036
rect 28224 9024 28230 9036
rect 28445 9027 28503 9033
rect 28445 9024 28457 9027
rect 28224 8996 28457 9024
rect 28224 8984 28230 8996
rect 28445 8993 28457 8996
rect 28491 8993 28503 9027
rect 28445 8987 28503 8993
rect 30006 8984 30012 9036
rect 30064 9033 30070 9036
rect 30300 9033 30328 9064
rect 30064 8987 30076 9033
rect 30285 9027 30343 9033
rect 30285 8993 30297 9027
rect 30331 8993 30343 9027
rect 30285 8987 30343 8993
rect 30064 8984 30070 8987
rect 25424 8956 25452 8984
rect 25056 8928 25268 8956
rect 25424 8928 26832 8956
rect 25240 8900 25268 8928
rect 25222 8848 25228 8900
rect 25280 8848 25286 8900
rect 25961 8891 26019 8897
rect 25961 8857 25973 8891
rect 26007 8888 26019 8891
rect 26418 8888 26424 8900
rect 26007 8860 26424 8888
rect 26007 8857 26019 8860
rect 25961 8851 26019 8857
rect 26418 8848 26424 8860
rect 26476 8848 26482 8900
rect 26804 8832 26832 8928
rect 20312 8792 23336 8820
rect 23753 8823 23811 8829
rect 20312 8780 20318 8792
rect 23753 8789 23765 8823
rect 23799 8820 23811 8823
rect 24026 8820 24032 8832
rect 23799 8792 24032 8820
rect 23799 8789 23811 8792
rect 23753 8783 23811 8789
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 25590 8780 25596 8832
rect 25648 8780 25654 8832
rect 25774 8780 25780 8832
rect 25832 8780 25838 8832
rect 26786 8780 26792 8832
rect 26844 8820 26850 8832
rect 26881 8823 26939 8829
rect 26881 8820 26893 8823
rect 26844 8792 26893 8820
rect 26844 8780 26850 8792
rect 26881 8789 26893 8792
rect 26927 8789 26939 8823
rect 26881 8783 26939 8789
rect 552 8730 31648 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 11436 8730
rect 11488 8678 11500 8730
rect 11552 8678 11564 8730
rect 11616 8678 11628 8730
rect 11680 8678 11692 8730
rect 11744 8678 19210 8730
rect 19262 8678 19274 8730
rect 19326 8678 19338 8730
rect 19390 8678 19402 8730
rect 19454 8678 19466 8730
rect 19518 8678 26984 8730
rect 27036 8678 27048 8730
rect 27100 8678 27112 8730
rect 27164 8678 27176 8730
rect 27228 8678 27240 8730
rect 27292 8678 31648 8730
rect 552 8656 31648 8678
rect 2314 8576 2320 8628
rect 2372 8576 2378 8628
rect 4706 8576 4712 8628
rect 4764 8576 4770 8628
rect 6365 8619 6423 8625
rect 6365 8585 6377 8619
rect 6411 8616 6423 8619
rect 9306 8616 9312 8628
rect 6411 8588 9312 8616
rect 6411 8585 6423 8588
rect 6365 8579 6423 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 11606 8616 11612 8628
rect 9824 8588 11612 8616
rect 9824 8576 9830 8588
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 14001 8619 14059 8625
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 14550 8616 14556 8628
rect 14047 8588 14556 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18230 8616 18236 8628
rect 18187 8588 18236 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 23106 8616 23112 8628
rect 22296 8588 23112 8616
rect 4893 8551 4951 8557
rect 4893 8517 4905 8551
rect 4939 8548 4951 8551
rect 7101 8551 7159 8557
rect 4939 8520 6132 8548
rect 4939 8517 4951 8520
rect 4893 8511 4951 8517
rect 3418 8480 3424 8492
rect 2516 8452 3424 8480
rect 2516 8421 2544 8452
rect 3418 8440 3424 8452
rect 3476 8440 3482 8492
rect 6104 8489 6132 8520
rect 7101 8517 7113 8551
rect 7147 8548 7159 8551
rect 7282 8548 7288 8560
rect 7147 8520 7288 8548
rect 7147 8517 7159 8520
rect 7101 8511 7159 8517
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 14185 8551 14243 8557
rect 14185 8548 14197 8551
rect 12406 8520 14197 8548
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8449 6147 8483
rect 6914 8480 6920 8492
rect 6089 8443 6147 8449
rect 6380 8452 6920 8480
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 2866 8412 2872 8424
rect 2731 8384 2872 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 3050 8372 3056 8424
rect 3108 8412 3114 8424
rect 4246 8412 4252 8424
rect 3108 8384 4252 8412
rect 3108 8372 3114 8384
rect 4246 8372 4252 8384
rect 4304 8412 4310 8424
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 4304 8384 4537 8412
rect 4304 8372 4310 8384
rect 4525 8381 4537 8384
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 5166 8412 5172 8424
rect 4755 8384 5172 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 4982 8304 4988 8356
rect 5040 8344 5046 8356
rect 5276 8344 5304 8375
rect 6270 8372 6276 8424
rect 6328 8372 6334 8424
rect 6380 8421 6408 8452
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7466 8480 7472 8492
rect 7116 8452 7472 8480
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 6822 8372 6828 8424
rect 6880 8372 6886 8424
rect 7116 8421 7144 8452
rect 7466 8440 7472 8452
rect 7524 8480 7530 8492
rect 12406 8480 12434 8520
rect 14185 8517 14197 8520
rect 14231 8548 14243 8551
rect 15470 8548 15476 8560
rect 14231 8520 15476 8548
rect 14231 8517 14243 8520
rect 14185 8511 14243 8517
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 15930 8508 15936 8560
rect 15988 8548 15994 8560
rect 15988 8520 19012 8548
rect 15988 8508 15994 8520
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 7524 8452 12434 8480
rect 18340 8452 18705 8480
rect 7524 8440 7530 8452
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7650 8372 7656 8424
rect 7708 8372 7714 8424
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8812 8384 9321 8412
rect 8812 8372 8818 8384
rect 9309 8381 9321 8384
rect 9355 8412 9367 8415
rect 9950 8412 9956 8424
rect 9355 8384 9956 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 11974 8372 11980 8424
rect 12032 8372 12038 8424
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8412 15991 8415
rect 16206 8412 16212 8424
rect 15979 8384 16212 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 18340 8421 18368 8452
rect 18693 8449 18705 8452
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 18414 8372 18420 8424
rect 18472 8372 18478 8424
rect 18874 8372 18880 8424
rect 18932 8372 18938 8424
rect 18984 8412 19012 8520
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8480 19395 8483
rect 21542 8480 21548 8492
rect 19383 8452 21548 8480
rect 19383 8449 19395 8452
rect 19337 8443 19395 8449
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 18984 8384 19073 8412
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 19150 8372 19156 8424
rect 19208 8421 19214 8424
rect 19208 8415 19237 8421
rect 19225 8381 19237 8415
rect 19429 8415 19487 8421
rect 19429 8412 19441 8415
rect 19208 8375 19237 8381
rect 19352 8384 19441 8412
rect 19208 8372 19214 8375
rect 5040 8316 5304 8344
rect 7745 8347 7803 8353
rect 5040 8304 5046 8316
rect 7745 8313 7757 8347
rect 7791 8344 7803 8347
rect 9582 8344 9588 8356
rect 7791 8316 9588 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 10594 8304 10600 8356
rect 10652 8344 10658 8356
rect 13817 8347 13875 8353
rect 13817 8344 13829 8347
rect 10652 8316 13829 8344
rect 10652 8304 10658 8316
rect 13817 8313 13829 8316
rect 13863 8313 13875 8347
rect 13817 8307 13875 8313
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 18966 8344 18972 8356
rect 16724 8316 18972 8344
rect 16724 8304 16730 8316
rect 18966 8304 18972 8316
rect 19024 8304 19030 8356
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 8478 8276 8484 8288
rect 4948 8248 8484 8276
rect 4948 8236 4954 8248
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 9217 8279 9275 8285
rect 9217 8276 9229 8279
rect 8628 8248 9229 8276
rect 8628 8236 8634 8248
rect 9217 8245 9229 8248
rect 9263 8245 9275 8279
rect 9217 8239 9275 8245
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 14001 8279 14059 8285
rect 14001 8276 14013 8279
rect 11020 8248 14013 8276
rect 11020 8236 11026 8248
rect 14001 8245 14013 8248
rect 14047 8276 14059 8279
rect 14826 8276 14832 8288
rect 14047 8248 14832 8276
rect 14047 8245 14059 8248
rect 14001 8239 14059 8245
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15344 8248 15853 8276
rect 15344 8236 15350 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 15841 8239 15899 8245
rect 18782 8236 18788 8288
rect 18840 8276 18846 8288
rect 19352 8276 19380 8384
rect 19429 8381 19441 8384
rect 19475 8381 19487 8415
rect 19429 8375 19487 8381
rect 19610 8372 19616 8424
rect 19668 8372 19674 8424
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 22296 8421 22324 8588
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 23198 8576 23204 8628
rect 23256 8616 23262 8628
rect 23256 8588 24440 8616
rect 23256 8576 23262 8588
rect 23845 8551 23903 8557
rect 23845 8548 23857 8551
rect 22480 8520 23857 8548
rect 22480 8421 22508 8520
rect 23845 8517 23857 8520
rect 23891 8517 23903 8551
rect 23845 8511 23903 8517
rect 22830 8480 22836 8492
rect 22572 8452 22836 8480
rect 22572 8421 22600 8452
rect 22830 8440 22836 8452
rect 22888 8480 22894 8492
rect 23661 8483 23719 8489
rect 22888 8452 23336 8480
rect 22888 8440 22894 8452
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20496 8384 21005 8412
rect 20496 8372 20502 8384
rect 20993 8381 21005 8384
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 22189 8415 22247 8421
rect 22189 8381 22201 8415
rect 22235 8381 22247 8415
rect 22189 8375 22247 8381
rect 22281 8415 22339 8421
rect 22281 8381 22293 8415
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 22465 8415 22523 8421
rect 22465 8381 22477 8415
rect 22511 8381 22523 8415
rect 22465 8375 22523 8381
rect 22557 8415 22615 8421
rect 22557 8381 22569 8415
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 22204 8344 22232 8375
rect 22646 8372 22652 8424
rect 22704 8372 22710 8424
rect 23017 8415 23075 8421
rect 23017 8381 23029 8415
rect 23063 8412 23075 8415
rect 23106 8412 23112 8424
rect 23063 8384 23112 8412
rect 23063 8381 23075 8384
rect 23017 8375 23075 8381
rect 23106 8372 23112 8384
rect 23164 8372 23170 8424
rect 23198 8372 23204 8424
rect 23256 8372 23262 8424
rect 23308 8421 23336 8452
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 24302 8480 24308 8492
rect 23707 8452 24308 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 24302 8440 24308 8452
rect 24360 8440 24366 8492
rect 24412 8480 24440 8588
rect 24486 8576 24492 8628
rect 24544 8576 24550 8628
rect 26142 8576 26148 8628
rect 26200 8616 26206 8628
rect 27157 8619 27215 8625
rect 27157 8616 27169 8619
rect 26200 8588 27169 8616
rect 26200 8576 26206 8588
rect 27157 8585 27169 8588
rect 27203 8585 27215 8619
rect 27157 8579 27215 8585
rect 28166 8576 28172 8628
rect 28224 8616 28230 8628
rect 28813 8619 28871 8625
rect 28813 8616 28825 8619
rect 28224 8588 28825 8616
rect 28224 8576 28230 8588
rect 28813 8585 28825 8588
rect 28859 8585 28871 8619
rect 28813 8579 28871 8585
rect 29917 8619 29975 8625
rect 29917 8585 29929 8619
rect 29963 8616 29975 8619
rect 30006 8616 30012 8628
rect 29963 8588 30012 8616
rect 29963 8585 29975 8588
rect 29917 8579 29975 8585
rect 30006 8576 30012 8588
rect 30064 8576 30070 8628
rect 24578 8508 24584 8560
rect 24636 8508 24642 8560
rect 25409 8483 25467 8489
rect 25409 8480 25421 8483
rect 24412 8452 25421 8480
rect 25409 8449 25421 8452
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 25590 8440 25596 8492
rect 25648 8480 25654 8492
rect 25777 8483 25835 8489
rect 25777 8480 25789 8483
rect 25648 8452 25789 8480
rect 25648 8440 25654 8452
rect 25777 8449 25789 8452
rect 25823 8449 25835 8483
rect 25777 8443 25835 8449
rect 28994 8440 29000 8492
rect 29052 8440 29058 8492
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8381 23351 8415
rect 23293 8375 23351 8381
rect 23382 8372 23388 8424
rect 23440 8372 23446 8424
rect 25685 8415 25743 8421
rect 25685 8412 25697 8415
rect 23492 8384 25697 8412
rect 22738 8344 22744 8356
rect 22204 8316 22744 8344
rect 22738 8304 22744 8316
rect 22796 8344 22802 8356
rect 23492 8344 23520 8384
rect 25685 8381 25697 8384
rect 25731 8412 25743 8415
rect 26326 8412 26332 8424
rect 25731 8384 26332 8412
rect 25731 8381 25743 8384
rect 25685 8375 25743 8381
rect 26326 8372 26332 8384
rect 26384 8412 26390 8424
rect 27338 8412 27344 8424
rect 26384 8384 27344 8412
rect 26384 8372 26390 8384
rect 27338 8372 27344 8384
rect 27396 8372 27402 8424
rect 27433 8415 27491 8421
rect 27433 8381 27445 8415
rect 27479 8412 27491 8415
rect 27982 8412 27988 8424
rect 27479 8384 27988 8412
rect 27479 8381 27491 8384
rect 27433 8375 27491 8381
rect 27982 8372 27988 8384
rect 28040 8372 28046 8424
rect 28810 8372 28816 8424
rect 28868 8412 28874 8424
rect 29733 8415 29791 8421
rect 29733 8412 29745 8415
rect 28868 8384 29745 8412
rect 28868 8372 28874 8384
rect 29733 8381 29745 8384
rect 29779 8381 29791 8415
rect 29733 8375 29791 8381
rect 29917 8415 29975 8421
rect 29917 8381 29929 8415
rect 29963 8381 29975 8415
rect 29917 8375 29975 8381
rect 22796 8316 23520 8344
rect 22796 8304 22802 8316
rect 24026 8304 24032 8356
rect 24084 8304 24090 8356
rect 24210 8304 24216 8356
rect 24268 8304 24274 8356
rect 24854 8304 24860 8356
rect 24912 8344 24918 8356
rect 24949 8347 25007 8353
rect 24949 8344 24961 8347
rect 24912 8316 24961 8344
rect 24912 8304 24918 8316
rect 24949 8313 24961 8316
rect 24995 8313 25007 8347
rect 24949 8307 25007 8313
rect 25041 8347 25099 8353
rect 25041 8313 25053 8347
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 18840 8248 19380 8276
rect 18840 8236 18846 8248
rect 19794 8236 19800 8288
rect 19852 8236 19858 8288
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 22094 8236 22100 8288
rect 22152 8236 22158 8288
rect 22925 8279 22983 8285
rect 22925 8245 22937 8279
rect 22971 8276 22983 8279
rect 23014 8276 23020 8288
rect 22971 8248 23020 8276
rect 22971 8245 22983 8248
rect 22925 8239 22983 8245
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 24228 8276 24256 8304
rect 25056 8276 25084 8307
rect 25222 8304 25228 8356
rect 25280 8304 25286 8356
rect 25774 8304 25780 8356
rect 25832 8344 25838 8356
rect 26022 8347 26080 8353
rect 26022 8344 26034 8347
rect 25832 8316 26034 8344
rect 25832 8304 25838 8316
rect 26022 8313 26034 8316
rect 26068 8313 26080 8347
rect 26022 8307 26080 8313
rect 27522 8304 27528 8356
rect 27580 8344 27586 8356
rect 27678 8347 27736 8353
rect 27678 8344 27690 8347
rect 27580 8316 27690 8344
rect 27580 8304 27586 8316
rect 27678 8313 27690 8316
rect 27724 8313 27736 8347
rect 27678 8307 27736 8313
rect 29641 8347 29699 8353
rect 29641 8313 29653 8347
rect 29687 8344 29699 8347
rect 29932 8344 29960 8375
rect 29687 8316 29960 8344
rect 29687 8313 29699 8316
rect 29641 8307 29699 8313
rect 24228 8248 25084 8276
rect 25590 8236 25596 8288
rect 25648 8236 25654 8288
rect 552 8186 31648 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 12096 8186
rect 12148 8134 12160 8186
rect 12212 8134 12224 8186
rect 12276 8134 12288 8186
rect 12340 8134 12352 8186
rect 12404 8134 19870 8186
rect 19922 8134 19934 8186
rect 19986 8134 19998 8186
rect 20050 8134 20062 8186
rect 20114 8134 20126 8186
rect 20178 8134 27644 8186
rect 27696 8134 27708 8186
rect 27760 8134 27772 8186
rect 27824 8134 27836 8186
rect 27888 8134 27900 8186
rect 27952 8134 31648 8186
rect 552 8112 31648 8134
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 6822 8072 6828 8084
rect 5123 8044 6828 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 6914 8032 6920 8084
rect 6972 8032 6978 8084
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 7190 8072 7196 8084
rect 7064 8044 7196 8072
rect 7064 8032 7070 8044
rect 7190 8032 7196 8044
rect 7248 8072 7254 8084
rect 9766 8072 9772 8084
rect 7248 8044 9772 8072
rect 7248 8032 7254 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9916 8044 10149 8072
rect 9916 8032 9922 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 18598 8072 18604 8084
rect 14608 8044 18604 8072
rect 14608 8032 14614 8044
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 18874 8072 18880 8084
rect 18748 8044 18880 8072
rect 18748 8032 18754 8044
rect 18874 8032 18880 8044
rect 18932 8072 18938 8084
rect 19337 8075 19395 8081
rect 18932 8044 19196 8072
rect 18932 8032 18938 8044
rect 1394 7964 1400 8016
rect 1452 8004 1458 8016
rect 4982 8004 4988 8016
rect 1452 7976 4988 8004
rect 1452 7964 1458 7976
rect 2884 7945 2912 7976
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 5261 8007 5319 8013
rect 5261 7973 5273 8007
rect 5307 8004 5319 8007
rect 6086 8004 6092 8016
rect 5307 7976 6092 8004
rect 5307 7973 5319 7976
rect 5261 7967 5319 7973
rect 6086 7964 6092 7976
rect 6144 8004 6150 8016
rect 6457 8007 6515 8013
rect 6457 8004 6469 8007
rect 6144 7976 6469 8004
rect 6144 7964 6150 7976
rect 6457 7973 6469 7976
rect 6503 7973 6515 8007
rect 6457 7967 6515 7973
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 7377 8007 7435 8013
rect 7377 8004 7389 8007
rect 6788 7976 7389 8004
rect 6788 7964 6794 7976
rect 7377 7973 7389 7976
rect 7423 7973 7435 8007
rect 9490 8004 9496 8016
rect 7377 7967 7435 7973
rect 7944 7976 9496 8004
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 2869 7939 2927 7945
rect 2363 7934 2544 7936
rect 2363 7908 2636 7934
rect 2363 7905 2375 7908
rect 2516 7906 2636 7908
rect 2317 7899 2375 7905
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2608 7868 2636 7906
rect 2869 7905 2881 7939
rect 2915 7905 2927 7939
rect 2869 7899 2927 7905
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7936 4767 7939
rect 4890 7936 4896 7948
rect 4755 7908 4896 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5166 7896 5172 7948
rect 5224 7896 5230 7948
rect 6178 7896 6184 7948
rect 6236 7936 6242 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 6236 7908 6285 7936
rect 6236 7896 6242 7908
rect 6273 7905 6285 7908
rect 6319 7905 6331 7939
rect 6273 7899 6331 7905
rect 6546 7896 6552 7948
rect 6604 7896 6610 7948
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 3234 7868 3240 7880
rect 2608 7840 3240 7868
rect 2501 7831 2559 7837
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2516 7800 2544 7831
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4304 7840 4629 7868
rect 4304 7828 4310 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6656 7868 6684 7899
rect 7006 7896 7012 7948
rect 7064 7936 7070 7948
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 7064 7908 7113 7936
rect 7064 7896 7070 7908
rect 7101 7905 7113 7908
rect 7147 7905 7159 7939
rect 7101 7899 7159 7905
rect 7190 7896 7196 7948
rect 7248 7896 7254 7948
rect 7650 7896 7656 7948
rect 7708 7896 7714 7948
rect 7742 7896 7748 7948
rect 7800 7896 7806 7948
rect 7834 7896 7840 7948
rect 7892 7896 7898 7948
rect 7944 7868 7972 7976
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 11072 7976 11284 8004
rect 9953 7963 10011 7969
rect 8481 7939 8539 7945
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 8846 7936 8852 7948
rect 8527 7908 8852 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8846 7896 8852 7908
rect 8904 7936 8910 7948
rect 9122 7936 9128 7948
rect 8904 7908 9128 7936
rect 8904 7896 8910 7908
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 9768 7939 9826 7945
rect 9768 7936 9780 7939
rect 9732 7908 9780 7936
rect 9732 7896 9738 7908
rect 9768 7905 9780 7908
rect 9814 7905 9826 7939
rect 9768 7899 9826 7905
rect 9858 7896 9864 7948
rect 9916 7896 9922 7948
rect 9953 7929 9965 7963
rect 9999 7936 10011 7963
rect 10962 7936 10968 7948
rect 9999 7929 10968 7936
rect 9953 7923 10968 7929
rect 9968 7908 10968 7923
rect 9968 7880 9996 7908
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 6420 7840 6684 7868
rect 6748 7840 7972 7868
rect 8021 7871 8079 7877
rect 6420 7828 6426 7840
rect 6748 7800 6776 7840
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8294 7868 8300 7880
rect 8067 7840 8300 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 8662 7868 8668 7880
rect 8619 7840 8668 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 8772 7840 9904 7868
rect 2372 7772 6776 7800
rect 7469 7803 7527 7809
rect 2372 7760 2378 7772
rect 7469 7769 7481 7803
rect 7515 7800 7527 7803
rect 8772 7800 8800 7840
rect 7515 7772 8800 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 8846 7760 8852 7812
rect 8904 7760 8910 7812
rect 9033 7803 9091 7809
rect 9033 7769 9045 7803
rect 9079 7800 9091 7803
rect 9306 7800 9312 7812
rect 9079 7772 9312 7800
rect 9079 7769 9091 7772
rect 9033 7763 9091 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 9490 7760 9496 7812
rect 9548 7760 9554 7812
rect 9876 7800 9904 7840
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 11072 7800 11100 7976
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7905 11207 7939
rect 11256 7936 11284 7976
rect 11330 7964 11336 8016
rect 11388 8004 11394 8016
rect 11606 8004 11612 8016
rect 11388 7976 11612 8004
rect 11388 7964 11394 7976
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 12805 8007 12863 8013
rect 12805 7973 12817 8007
rect 12851 8004 12863 8007
rect 13262 8004 13268 8016
rect 12851 7976 13268 8004
rect 12851 7973 12863 7976
rect 12805 7967 12863 7973
rect 13262 7964 13268 7976
rect 13320 8004 13326 8016
rect 15838 8004 15844 8016
rect 13320 7976 14044 8004
rect 13320 7964 13326 7976
rect 11256 7908 11376 7936
rect 11149 7899 11207 7905
rect 9876 7772 11100 7800
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 2133 7735 2191 7741
rect 2133 7732 2145 7735
rect 2004 7704 2145 7732
rect 2004 7692 2010 7704
rect 2133 7701 2145 7704
rect 2179 7701 2191 7735
rect 2133 7695 2191 7701
rect 2774 7692 2780 7744
rect 2832 7692 2838 7744
rect 6825 7735 6883 7741
rect 6825 7701 6837 7735
rect 6871 7732 6883 7735
rect 7006 7732 7012 7744
rect 6871 7704 7012 7732
rect 6871 7701 6883 7704
rect 6825 7695 6883 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7377 7735 7435 7741
rect 7377 7701 7389 7735
rect 7423 7732 7435 7735
rect 7558 7732 7564 7744
rect 7423 7704 7564 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 8260 7704 8401 7732
rect 8260 7692 8266 7704
rect 8389 7701 8401 7704
rect 8435 7701 8447 7735
rect 8389 7695 8447 7701
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 11164 7732 11192 7899
rect 11238 7828 11244 7880
rect 11296 7828 11302 7880
rect 11348 7800 11376 7908
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 12032 7908 12357 7936
rect 12032 7896 12038 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12710 7896 12716 7948
rect 12768 7896 12774 7948
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12952 7908 13001 7936
rect 12952 7896 12958 7908
rect 12989 7905 13001 7908
rect 13035 7905 13047 7939
rect 12989 7899 13047 7905
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7905 13139 7939
rect 13081 7899 13139 7905
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 13096 7868 13124 7899
rect 13170 7896 13176 7948
rect 13228 7936 13234 7948
rect 13357 7939 13415 7945
rect 13228 7908 13273 7936
rect 13228 7896 13234 7908
rect 13357 7905 13369 7939
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 11563 7840 13124 7868
rect 13372 7868 13400 7899
rect 13446 7896 13452 7948
rect 13504 7896 13510 7948
rect 13538 7896 13544 7948
rect 13596 7945 13602 7948
rect 13596 7936 13604 7945
rect 13596 7908 13641 7936
rect 13596 7899 13604 7908
rect 13596 7896 13602 7899
rect 14016 7880 14044 7976
rect 14936 7976 15844 8004
rect 13372 7840 13492 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 13262 7800 13268 7812
rect 11348 7772 13268 7800
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 13464 7800 13492 7840
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 14056 7840 14381 7868
rect 14056 7828 14062 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 14516 7840 14749 7868
rect 14516 7828 14522 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14936 7868 14964 7976
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 16390 7964 16396 8016
rect 16448 8004 16454 8016
rect 19061 8007 19119 8013
rect 19061 8004 19073 8007
rect 16448 7976 19073 8004
rect 16448 7964 16454 7976
rect 19061 7973 19073 7976
rect 19107 7973 19119 8007
rect 19061 7967 19119 7973
rect 15013 7939 15071 7945
rect 15013 7905 15025 7939
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 14737 7831 14795 7837
rect 14844 7840 14964 7868
rect 15028 7868 15056 7899
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 15286 7896 15292 7948
rect 15344 7896 15350 7948
rect 15562 7896 15568 7948
rect 15620 7896 15626 7948
rect 18874 7945 18880 7948
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 18432 7908 18705 7936
rect 15378 7868 15384 7880
rect 15028 7840 15384 7868
rect 14844 7800 14872 7840
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7868 15715 7871
rect 16666 7868 16672 7880
rect 15703 7840 16672 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7868 16819 7871
rect 17034 7868 17040 7880
rect 16807 7840 17040 7868
rect 16807 7837 16819 7840
rect 16761 7831 16819 7837
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 13464 7772 14872 7800
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7800 14979 7803
rect 16485 7803 16543 7809
rect 14967 7772 15516 7800
rect 14967 7769 14979 7772
rect 14921 7763 14979 7769
rect 15488 7744 15516 7772
rect 16485 7769 16497 7803
rect 16531 7800 16543 7803
rect 17402 7800 17408 7812
rect 16531 7772 17408 7800
rect 16531 7769 16543 7772
rect 16485 7763 16543 7769
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 8536 7704 11192 7732
rect 8536 7692 8542 7704
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12584 7704 13001 7732
rect 12584 7692 12590 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 12989 7695 13047 7701
rect 13722 7692 13728 7744
rect 13780 7692 13786 7744
rect 13817 7735 13875 7741
rect 13817 7701 13829 7735
rect 13863 7732 13875 7735
rect 13906 7732 13912 7744
rect 13863 7704 13912 7732
rect 13863 7701 13875 7704
rect 13817 7695 13875 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14792 7704 14841 7732
rect 14792 7692 14798 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 14829 7695 14887 7701
rect 15102 7692 15108 7744
rect 15160 7732 15166 7744
rect 15289 7735 15347 7741
rect 15289 7732 15301 7735
rect 15160 7704 15301 7732
rect 15160 7692 15166 7704
rect 15289 7701 15301 7704
rect 15335 7701 15347 7735
rect 15289 7695 15347 7701
rect 15470 7692 15476 7744
rect 15528 7692 15534 7744
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15712 7704 15853 7732
rect 15712 7692 15718 7704
rect 15841 7701 15853 7704
rect 15887 7701 15899 7735
rect 15841 7695 15899 7701
rect 16298 7692 16304 7744
rect 16356 7692 16362 7744
rect 18432 7732 18460 7908
rect 18693 7905 18705 7908
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 18831 7939 18880 7945
rect 18831 7905 18843 7939
rect 18877 7905 18880 7939
rect 18831 7899 18880 7905
rect 18874 7896 18880 7899
rect 18932 7896 18938 7948
rect 18969 7939 19027 7945
rect 18969 7905 18981 7939
rect 19015 7905 19027 7939
rect 18969 7899 19027 7905
rect 18506 7828 18512 7880
rect 18564 7868 18570 7880
rect 18984 7868 19012 7899
rect 18564 7840 19012 7868
rect 18564 7828 18570 7840
rect 19076 7800 19104 7967
rect 19168 7945 19196 8044
rect 19337 8041 19349 8075
rect 19383 8072 19395 8075
rect 19610 8072 19616 8084
rect 19383 8044 19616 8072
rect 19383 8041 19395 8044
rect 19337 8035 19395 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 24121 8075 24179 8081
rect 24121 8041 24133 8075
rect 24167 8072 24179 8075
rect 24578 8072 24584 8084
rect 24167 8044 24584 8072
rect 24167 8041 24179 8044
rect 24121 8035 24179 8041
rect 24578 8032 24584 8044
rect 24636 8032 24642 8084
rect 27157 8075 27215 8081
rect 27157 8041 27169 8075
rect 27203 8072 27215 8075
rect 27522 8072 27528 8084
rect 27203 8044 27528 8072
rect 27203 8041 27215 8044
rect 27157 8035 27215 8041
rect 27522 8032 27528 8044
rect 27580 8032 27586 8084
rect 27617 8075 27675 8081
rect 27617 8041 27629 8075
rect 27663 8072 27675 8075
rect 27982 8072 27988 8084
rect 27663 8044 27988 8072
rect 27663 8041 27675 8044
rect 27617 8035 27675 8041
rect 27982 8032 27988 8044
rect 28040 8032 28046 8084
rect 19794 7964 19800 8016
rect 19852 8004 19858 8016
rect 20542 8007 20600 8013
rect 20542 8004 20554 8007
rect 19852 7976 20554 8004
rect 19852 7964 19858 7976
rect 20542 7973 20554 7976
rect 20588 7973 20600 8007
rect 25590 8004 25596 8016
rect 20542 7967 20600 7973
rect 24228 7976 25596 8004
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7936 19211 7939
rect 20714 7936 20720 7948
rect 19199 7908 20720 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 20809 7939 20867 7945
rect 20809 7905 20821 7939
rect 20855 7936 20867 7939
rect 20898 7936 20904 7948
rect 20855 7908 20904 7936
rect 20855 7905 20867 7908
rect 20809 7899 20867 7905
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 23014 7945 23020 7948
rect 22741 7939 22799 7945
rect 22741 7936 22753 7939
rect 22152 7908 22753 7936
rect 22152 7896 22158 7908
rect 22741 7905 22753 7908
rect 22787 7905 22799 7939
rect 23008 7936 23020 7945
rect 22975 7908 23020 7936
rect 22741 7899 22799 7905
rect 23008 7899 23020 7908
rect 23014 7896 23020 7899
rect 23072 7896 23078 7948
rect 24228 7945 24256 7976
rect 25590 7964 25596 7976
rect 25648 7964 25654 8016
rect 24213 7939 24271 7945
rect 24213 7905 24225 7939
rect 24259 7905 24271 7939
rect 24213 7899 24271 7905
rect 24302 7896 24308 7948
rect 24360 7936 24366 7948
rect 24469 7939 24527 7945
rect 24469 7936 24481 7939
rect 24360 7908 24481 7936
rect 24360 7896 24366 7908
rect 24469 7905 24481 7908
rect 24515 7905 24527 7939
rect 24469 7899 24527 7905
rect 26786 7896 26792 7948
rect 26844 7896 26850 7948
rect 27338 7896 27344 7948
rect 27396 7936 27402 7948
rect 27709 7939 27767 7945
rect 27709 7936 27721 7939
rect 27396 7908 27721 7936
rect 27396 7896 27402 7908
rect 27709 7905 27721 7908
rect 27755 7905 27767 7939
rect 27709 7899 27767 7905
rect 26234 7828 26240 7880
rect 26292 7868 26298 7880
rect 26697 7871 26755 7877
rect 26697 7868 26709 7871
rect 26292 7840 26709 7868
rect 26292 7828 26298 7840
rect 26697 7837 26709 7840
rect 26743 7837 26755 7871
rect 26697 7831 26755 7837
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 19076 7772 19441 7800
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 19429 7763 19487 7769
rect 25222 7760 25228 7812
rect 25280 7800 25286 7812
rect 25593 7803 25651 7809
rect 25593 7800 25605 7803
rect 25280 7772 25605 7800
rect 25280 7760 25286 7772
rect 25593 7769 25605 7772
rect 25639 7769 25651 7803
rect 25593 7763 25651 7769
rect 20990 7732 20996 7744
rect 18432 7704 20996 7732
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 552 7642 31648 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 11436 7642
rect 11488 7590 11500 7642
rect 11552 7590 11564 7642
rect 11616 7590 11628 7642
rect 11680 7590 11692 7642
rect 11744 7590 19210 7642
rect 19262 7590 19274 7642
rect 19326 7590 19338 7642
rect 19390 7590 19402 7642
rect 19454 7590 19466 7642
rect 19518 7590 26984 7642
rect 27036 7590 27048 7642
rect 27100 7590 27112 7642
rect 27164 7590 27176 7642
rect 27228 7590 27240 7642
rect 27292 7590 31648 7642
rect 552 7568 31648 7590
rect 3234 7488 3240 7540
rect 3292 7488 3298 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 7650 7528 7656 7540
rect 6687 7500 7656 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7800 7500 8033 7528
rect 7800 7488 7806 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8021 7491 8079 7497
rect 8938 7488 8944 7540
rect 8996 7488 9002 7540
rect 9048 7500 13676 7528
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7460 3111 7463
rect 3099 7432 6316 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 1305 7327 1363 7333
rect 1305 7293 1317 7327
rect 1351 7324 1363 7327
rect 1394 7324 1400 7336
rect 1351 7296 1400 7324
rect 1351 7293 1363 7296
rect 1305 7287 1363 7293
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 1946 7333 1952 7336
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7324 1547 7327
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1535 7296 1685 7324
rect 1535 7293 1547 7296
rect 1489 7287 1547 7293
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1940 7324 1952 7333
rect 1907 7296 1952 7324
rect 1673 7287 1731 7293
rect 1940 7287 1952 7296
rect 1946 7284 1952 7287
rect 2004 7284 2010 7336
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 3528 7333 3556 7432
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4706 7392 4712 7404
rect 4571 7364 4712 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6288 7401 6316 7432
rect 6546 7420 6552 7472
rect 6604 7460 6610 7472
rect 6604 7432 6868 7460
rect 6604 7420 6610 7432
rect 6273 7395 6331 7401
rect 6273 7361 6285 7395
rect 6319 7392 6331 7395
rect 6730 7392 6736 7404
rect 6319 7364 6736 7392
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7293 3571 7327
rect 3513 7287 3571 7293
rect 3878 7284 3884 7336
rect 3936 7284 3942 7336
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 4816 7296 5917 7324
rect 3326 7216 3332 7268
rect 3384 7256 3390 7268
rect 3605 7259 3663 7265
rect 3605 7256 3617 7259
rect 3384 7228 3617 7256
rect 3384 7216 3390 7228
rect 3605 7225 3617 7228
rect 3651 7225 3663 7259
rect 3605 7219 3663 7225
rect 3723 7259 3781 7265
rect 3723 7225 3735 7259
rect 3769 7225 3781 7259
rect 3723 7219 3781 7225
rect 1210 7148 1216 7200
rect 1268 7148 1274 7200
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 3738 7188 3766 7219
rect 4154 7188 4160 7200
rect 3200 7160 4160 7188
rect 3200 7148 3206 7160
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4816 7197 4844 7296
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 6086 7284 6092 7336
rect 6144 7284 6150 7336
rect 6196 7256 6224 7352
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7324 6515 7327
rect 6546 7324 6552 7336
rect 6503 7296 6552 7324
rect 6503 7293 6515 7296
rect 6457 7287 6515 7293
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 6638 7256 6644 7268
rect 6196 7228 6644 7256
rect 6638 7216 6644 7228
rect 6696 7216 6702 7268
rect 6840 7256 6868 7432
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 9048 7460 9076 7500
rect 6972 7432 7328 7460
rect 6972 7420 6978 7432
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7300 7333 7328 7432
rect 8772 7432 9076 7460
rect 9585 7463 9643 7469
rect 7558 7352 7564 7404
rect 7616 7352 7622 7404
rect 8772 7392 8800 7432
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 10318 7460 10324 7472
rect 9631 7432 10324 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 10318 7420 10324 7432
rect 10376 7460 10382 7472
rect 10686 7460 10692 7472
rect 10376 7432 10692 7460
rect 10376 7420 10382 7432
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 13262 7420 13268 7472
rect 13320 7420 13326 7472
rect 7852 7364 8800 7392
rect 7852 7333 7880 7364
rect 7009 7327 7067 7333
rect 7009 7324 7021 7327
rect 6972 7296 7021 7324
rect 6972 7284 6978 7296
rect 7009 7293 7021 7296
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7293 7711 7327
rect 7653 7287 7711 7293
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 6840 7228 6960 7256
rect 6932 7197 6960 7228
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 7484 7256 7512 7287
rect 7248 7228 7512 7256
rect 7668 7256 7696 7287
rect 8570 7284 8576 7336
rect 8628 7284 8634 7336
rect 8772 7333 8800 7364
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 8895 7364 9413 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9824 7364 9873 7392
rect 9824 7352 9830 7364
rect 9861 7361 9873 7364
rect 9907 7392 9919 7395
rect 13648 7392 13676 7500
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 13780 7500 13921 7528
rect 13780 7488 13786 7500
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 13909 7491 13967 7497
rect 13998 7488 14004 7540
rect 14056 7488 14062 7540
rect 14277 7531 14335 7537
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 14458 7528 14464 7540
rect 14323 7500 14464 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 14734 7488 14740 7540
rect 14792 7488 14798 7540
rect 15304 7500 16712 7528
rect 13817 7463 13875 7469
rect 13817 7429 13829 7463
rect 13863 7460 13875 7463
rect 15102 7460 15108 7472
rect 13863 7432 15108 7460
rect 13863 7429 13875 7432
rect 13817 7423 13875 7429
rect 15102 7420 15108 7432
rect 15160 7420 15166 7472
rect 9907 7364 10088 7392
rect 13648 7364 14780 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 10060 7324 10088 7364
rect 10167 7327 10225 7333
rect 10167 7324 10179 7327
rect 9140 7296 9996 7324
rect 10060 7296 10179 7324
rect 8588 7256 8616 7284
rect 7668 7228 8616 7256
rect 7248 7216 7254 7228
rect 4801 7191 4859 7197
rect 4801 7157 4813 7191
rect 4847 7157 4859 7191
rect 4801 7151 4859 7157
rect 6917 7191 6975 7197
rect 6917 7157 6929 7191
rect 6963 7188 6975 7191
rect 9140 7188 9168 7296
rect 9968 7256 9996 7296
rect 10167 7293 10179 7296
rect 10213 7293 10225 7327
rect 10167 7287 10225 7293
rect 10318 7284 10324 7336
rect 10376 7284 10382 7336
rect 10594 7284 10600 7336
rect 10652 7333 10658 7336
rect 10652 7327 10685 7333
rect 10673 7293 10685 7327
rect 10652 7287 10685 7293
rect 10652 7284 10658 7287
rect 10778 7284 10784 7336
rect 10836 7284 10842 7336
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 11790 7324 11796 7336
rect 11388 7296 11796 7324
rect 11388 7284 11394 7296
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 11882 7284 11888 7336
rect 11940 7284 11946 7336
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7324 13599 7327
rect 13630 7324 13636 7336
rect 13587 7296 13636 7324
rect 13587 7293 13599 7296
rect 13541 7287 13599 7293
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 14550 7284 14556 7336
rect 14608 7284 14614 7336
rect 9968 7228 10548 7256
rect 6963 7160 9168 7188
rect 6963 7157 6975 7160
rect 6917 7151 6975 7157
rect 9306 7148 9312 7200
rect 9364 7148 9370 7200
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9824 7160 9965 7188
rect 9824 7148 9830 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 10410 7148 10416 7200
rect 10468 7148 10474 7200
rect 10520 7188 10548 7228
rect 11054 7216 11060 7268
rect 11112 7216 11118 7268
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 12130 7259 12188 7265
rect 12130 7256 12142 7259
rect 11664 7228 12142 7256
rect 11664 7216 11670 7228
rect 12130 7225 12142 7228
rect 12176 7225 12188 7259
rect 13446 7256 13452 7268
rect 12130 7219 12188 7225
rect 13187 7228 13452 7256
rect 13187 7188 13215 7228
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 14369 7259 14427 7265
rect 14369 7256 14381 7259
rect 13780 7228 14381 7256
rect 13780 7216 13786 7228
rect 14369 7225 14381 7228
rect 14415 7225 14427 7259
rect 14752 7256 14780 7364
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 14918 7284 14924 7336
rect 14976 7284 14982 7336
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15068 7296 15113 7324
rect 15068 7284 15074 7296
rect 15194 7284 15200 7336
rect 15252 7284 15258 7336
rect 15304 7265 15332 7500
rect 15562 7420 15568 7472
rect 15620 7460 15626 7472
rect 15620 7432 16436 7460
rect 15620 7420 15626 7432
rect 15427 7327 15485 7333
rect 15427 7293 15439 7327
rect 15473 7324 15485 7327
rect 15562 7324 15568 7336
rect 15473 7296 15568 7324
rect 15473 7293 15485 7296
rect 15427 7287 15485 7293
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 15654 7284 15660 7336
rect 15712 7284 15718 7336
rect 15838 7284 15844 7336
rect 15896 7284 15902 7336
rect 15933 7327 15991 7333
rect 15933 7293 15945 7327
rect 15979 7293 15991 7327
rect 15933 7287 15991 7293
rect 16025 7327 16083 7333
rect 16025 7293 16037 7327
rect 16071 7324 16083 7327
rect 16114 7324 16120 7336
rect 16071 7296 16120 7324
rect 16071 7293 16083 7296
rect 16025 7287 16083 7293
rect 15289 7259 15347 7265
rect 15289 7256 15301 7259
rect 14752 7228 15301 7256
rect 14369 7219 14427 7225
rect 15289 7225 15301 7228
rect 15335 7225 15347 7259
rect 15948 7256 15976 7287
rect 16114 7284 16120 7296
rect 16172 7284 16178 7336
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7293 16267 7327
rect 16408 7324 16436 7432
rect 16684 7404 16712 7500
rect 18874 7488 18880 7540
rect 18932 7528 18938 7540
rect 21637 7531 21695 7537
rect 21637 7528 21649 7531
rect 18932 7500 21649 7528
rect 18932 7488 18938 7500
rect 21637 7497 21649 7500
rect 21683 7497 21695 7531
rect 21637 7491 21695 7497
rect 16666 7352 16672 7404
rect 16724 7352 16730 7404
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 19153 7395 19211 7401
rect 19153 7392 19165 7395
rect 18463 7364 19165 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 19153 7361 19165 7364
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 20438 7352 20444 7404
rect 20496 7392 20502 7404
rect 21361 7395 21419 7401
rect 21361 7392 21373 7395
rect 20496 7364 21373 7392
rect 20496 7352 20502 7364
rect 21361 7361 21373 7364
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 22281 7395 22339 7401
rect 21508 7364 22048 7392
rect 21508 7352 21514 7364
rect 16758 7324 16764 7336
rect 16408 7296 16764 7324
rect 16209 7287 16267 7293
rect 15289 7219 15347 7225
rect 15672 7228 15976 7256
rect 16224 7256 16252 7287
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 17402 7284 17408 7336
rect 17460 7284 17466 7336
rect 18325 7327 18383 7333
rect 18325 7293 18337 7327
rect 18371 7293 18383 7327
rect 18325 7287 18383 7293
rect 17129 7259 17187 7265
rect 16224 7228 16804 7256
rect 15672 7200 15700 7228
rect 16776 7200 16804 7228
rect 17129 7225 17141 7259
rect 17175 7256 17187 7259
rect 17313 7259 17371 7265
rect 17313 7256 17325 7259
rect 17175 7228 17325 7256
rect 17175 7225 17187 7228
rect 17129 7219 17187 7225
rect 17313 7225 17325 7228
rect 17359 7225 17371 7259
rect 17313 7219 17371 7225
rect 10520 7160 13215 7188
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 13814 7188 13820 7200
rect 13679 7160 13820 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 15562 7148 15568 7200
rect 15620 7148 15626 7200
rect 15654 7148 15660 7200
rect 15712 7148 15718 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 15804 7160 16405 7188
rect 15804 7148 15810 7160
rect 16393 7157 16405 7160
rect 16439 7157 16451 7191
rect 16393 7151 16451 7157
rect 16482 7148 16488 7200
rect 16540 7148 16546 7200
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 17420 7188 17448 7284
rect 18340 7256 18368 7287
rect 18782 7284 18788 7336
rect 18840 7284 18846 7336
rect 18874 7284 18880 7336
rect 18932 7284 18938 7336
rect 20456 7324 20484 7352
rect 18984 7296 20484 7324
rect 18984 7256 19012 7296
rect 20622 7284 20628 7336
rect 20680 7284 20686 7336
rect 20714 7284 20720 7336
rect 20772 7324 20778 7336
rect 22020 7333 22048 7364
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22370 7392 22376 7404
rect 22327 7364 22376 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22370 7352 22376 7364
rect 22428 7392 22434 7404
rect 23382 7392 23388 7404
rect 22428 7364 23388 7392
rect 22428 7352 22434 7364
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 20772 7296 21833 7324
rect 20772 7284 20778 7296
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 22005 7327 22063 7333
rect 22005 7293 22017 7327
rect 22051 7293 22063 7327
rect 22005 7287 22063 7293
rect 22557 7327 22615 7333
rect 22557 7293 22569 7327
rect 22603 7324 22615 7327
rect 22738 7324 22744 7336
rect 22603 7296 22744 7324
rect 22603 7293 22615 7296
rect 22557 7287 22615 7293
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 24854 7284 24860 7336
rect 24912 7324 24918 7336
rect 26053 7327 26111 7333
rect 26053 7324 26065 7327
rect 24912 7296 26065 7324
rect 24912 7284 24918 7296
rect 26053 7293 26065 7296
rect 26099 7293 26111 7327
rect 26053 7287 26111 7293
rect 26697 7327 26755 7333
rect 26697 7293 26709 7327
rect 26743 7324 26755 7327
rect 27338 7324 27344 7336
rect 26743 7296 27344 7324
rect 26743 7293 26755 7296
rect 26697 7287 26755 7293
rect 27338 7284 27344 7296
rect 27396 7324 27402 7336
rect 29181 7327 29239 7333
rect 29181 7324 29193 7327
rect 27396 7296 29193 7324
rect 27396 7284 27402 7296
rect 29181 7293 29193 7296
rect 29227 7324 29239 7327
rect 30374 7324 30380 7336
rect 29227 7296 30380 7324
rect 29227 7293 29239 7296
rect 29181 7287 29239 7293
rect 30374 7284 30380 7296
rect 30432 7284 30438 7336
rect 18340 7228 19012 7256
rect 19061 7259 19119 7265
rect 19061 7225 19073 7259
rect 19107 7256 19119 7259
rect 19398 7259 19456 7265
rect 19398 7256 19410 7259
rect 19107 7228 19410 7256
rect 19107 7225 19119 7228
rect 19061 7219 19119 7225
rect 19398 7225 19410 7228
rect 19444 7225 19456 7259
rect 19398 7219 19456 7225
rect 21913 7259 21971 7265
rect 21913 7225 21925 7259
rect 21959 7225 21971 7259
rect 21913 7219 21971 7225
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 17420 7160 20545 7188
rect 20533 7157 20545 7160
rect 20579 7188 20591 7191
rect 21928 7188 21956 7219
rect 22094 7216 22100 7268
rect 22152 7265 22158 7268
rect 22152 7259 22181 7265
rect 22169 7225 22181 7259
rect 27522 7256 27528 7268
rect 22152 7219 22181 7225
rect 26252 7228 27528 7256
rect 22152 7216 22158 7219
rect 26252 7200 26280 7228
rect 27522 7216 27528 7228
rect 27580 7216 27586 7268
rect 20579 7160 21956 7188
rect 20579 7157 20591 7160
rect 20533 7151 20591 7157
rect 22278 7148 22284 7200
rect 22336 7188 22342 7200
rect 22465 7191 22523 7197
rect 22465 7188 22477 7191
rect 22336 7160 22477 7188
rect 22336 7148 22342 7160
rect 22465 7157 22477 7160
rect 22511 7157 22523 7191
rect 22465 7151 22523 7157
rect 26234 7148 26240 7200
rect 26292 7148 26298 7200
rect 26418 7148 26424 7200
rect 26476 7188 26482 7200
rect 26605 7191 26663 7197
rect 26605 7188 26617 7191
rect 26476 7160 26617 7188
rect 26476 7148 26482 7160
rect 26605 7157 26617 7160
rect 26651 7157 26663 7191
rect 26605 7151 26663 7157
rect 29086 7148 29092 7200
rect 29144 7148 29150 7200
rect 552 7098 31648 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 12096 7098
rect 12148 7046 12160 7098
rect 12212 7046 12224 7098
rect 12276 7046 12288 7098
rect 12340 7046 12352 7098
rect 12404 7046 19870 7098
rect 19922 7046 19934 7098
rect 19986 7046 19998 7098
rect 20050 7046 20062 7098
rect 20114 7046 20126 7098
rect 20178 7046 27644 7098
rect 27696 7046 27708 7098
rect 27760 7046 27772 7098
rect 27824 7046 27836 7098
rect 27888 7046 27900 7098
rect 27952 7046 31648 7098
rect 552 7024 31648 7046
rect 2774 6984 2780 6996
rect 2746 6944 2780 6984
rect 2832 6944 2838 6996
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 6641 6987 6699 6993
rect 4212 6956 4594 6984
rect 4212 6944 4218 6956
rect 1121 6851 1179 6857
rect 1121 6817 1133 6851
rect 1167 6848 1179 6851
rect 1210 6848 1216 6860
rect 1167 6820 1216 6848
rect 1167 6817 1179 6820
rect 1121 6811 1179 6817
rect 1210 6808 1216 6820
rect 1268 6808 1274 6860
rect 1388 6851 1446 6857
rect 1388 6817 1400 6851
rect 1434 6848 1446 6851
rect 1946 6848 1952 6860
rect 1434 6820 1952 6848
rect 1434 6817 1446 6820
rect 1388 6811 1446 6817
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 2746 6848 2774 6944
rect 3326 6876 3332 6928
rect 3384 6916 3390 6928
rect 4566 6925 4594 6956
rect 6641 6953 6653 6987
rect 6687 6984 6699 6987
rect 7834 6984 7840 6996
rect 6687 6956 7840 6984
rect 6687 6953 6699 6956
rect 6641 6947 6699 6953
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10226 6984 10232 6996
rect 9732 6956 10232 6984
rect 9732 6944 9738 6956
rect 10226 6944 10232 6956
rect 10284 6984 10290 6996
rect 10778 6984 10784 6996
rect 10284 6956 10784 6984
rect 10284 6944 10290 6956
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 11882 6944 11888 6996
rect 11940 6984 11946 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11940 6956 12081 6984
rect 11940 6944 11946 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 13722 6984 13728 6996
rect 12069 6947 12127 6953
rect 13188 6956 13728 6984
rect 4433 6919 4491 6925
rect 4433 6916 4445 6919
rect 3384 6888 4445 6916
rect 3384 6876 3390 6888
rect 4433 6885 4445 6888
rect 4479 6885 4491 6919
rect 4433 6879 4491 6885
rect 4551 6919 4609 6925
rect 4551 6885 4563 6919
rect 4597 6885 4609 6919
rect 4551 6879 4609 6885
rect 6730 6876 6736 6928
rect 6788 6876 6794 6928
rect 7193 6919 7251 6925
rect 7193 6885 7205 6919
rect 7239 6916 7251 6919
rect 7374 6916 7380 6928
rect 7239 6888 7380 6916
rect 7239 6885 7251 6888
rect 7193 6879 7251 6885
rect 7374 6876 7380 6888
rect 7432 6916 7438 6928
rect 8570 6916 8576 6928
rect 7432 6888 7880 6916
rect 7432 6876 7438 6888
rect 2866 6857 2872 6860
rect 2639 6820 2774 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 2860 6811 2872 6857
rect 2866 6808 2872 6811
rect 2924 6808 2930 6860
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 4249 6851 4307 6857
rect 4249 6848 4261 6851
rect 3476 6820 4261 6848
rect 3476 6808 3482 6820
rect 4249 6817 4261 6820
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 4709 6851 4767 6857
rect 4709 6817 4721 6851
rect 4755 6848 4767 6851
rect 5074 6848 5080 6860
rect 4755 6820 5080 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 4356 6780 4384 6811
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 6089 6851 6147 6857
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6135 6820 6316 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6104 6780 6132 6811
rect 4356 6752 6132 6780
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 3528 6684 4077 6712
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3528 6644 3556 6684
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 3016 6616 3556 6644
rect 3973 6647 4031 6653
rect 3016 6604 3022 6616
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 4356 6644 4384 6752
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6288 6780 6316 6820
rect 6362 6808 6368 6860
rect 6420 6808 6426 6860
rect 6454 6808 6460 6860
rect 6512 6808 6518 6860
rect 6546 6808 6552 6860
rect 6604 6808 6610 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 6288 6752 6408 6780
rect 5905 6715 5963 6721
rect 5905 6681 5917 6715
rect 5951 6712 5963 6715
rect 6270 6712 6276 6724
rect 5951 6684 6276 6712
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 4019 6616 4384 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 6086 6604 6092 6656
rect 6144 6604 6150 6656
rect 6380 6644 6408 6752
rect 6840 6712 6868 6811
rect 6932 6780 6960 6811
rect 7006 6808 7012 6860
rect 7064 6848 7070 6860
rect 7852 6857 7880 6888
rect 8128 6888 8576 6916
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7064 6820 7757 6848
rect 7064 6808 7070 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 7838 6851 7896 6857
rect 7838 6817 7850 6851
rect 7884 6817 7896 6851
rect 7838 6811 7896 6817
rect 8018 6808 8024 6860
rect 8076 6808 8082 6860
rect 8128 6857 8156 6888
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 11606 6876 11612 6928
rect 11664 6916 11670 6928
rect 12345 6919 12403 6925
rect 12345 6916 12357 6919
rect 11664 6888 12357 6916
rect 11664 6876 11670 6888
rect 12345 6885 12357 6888
rect 12391 6885 12403 6919
rect 13188 6916 13216 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 15378 6944 15384 6996
rect 15436 6944 15442 6996
rect 15470 6944 15476 6996
rect 15528 6944 15534 6996
rect 18966 6944 18972 6996
rect 19024 6984 19030 6996
rect 22094 6984 22100 6996
rect 19024 6956 22100 6984
rect 19024 6944 19030 6956
rect 22094 6944 22100 6956
rect 22152 6944 22158 6996
rect 25777 6987 25835 6993
rect 25777 6953 25789 6987
rect 25823 6984 25835 6987
rect 25823 6956 25912 6984
rect 25823 6953 25835 6956
rect 25777 6947 25835 6953
rect 13538 6916 13544 6928
rect 12345 6879 12403 6885
rect 12728 6888 13216 6916
rect 12728 6860 12756 6888
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 8202 6808 8208 6860
rect 8260 6857 8266 6860
rect 8260 6848 8268 6857
rect 9217 6851 9275 6857
rect 8260 6820 8305 6848
rect 8260 6811 8268 6820
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9306 6848 9312 6860
rect 9263 6820 9312 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 8260 6808 8266 6811
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 7190 6780 7196 6792
rect 6932 6752 7196 6780
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7558 6780 7564 6792
rect 7392 6752 7564 6780
rect 7392 6712 7420 6752
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 9030 6780 9036 6792
rect 7699 6752 9036 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 9030 6740 9036 6752
rect 9088 6740 9094 6792
rect 9416 6780 9444 6811
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9640 6820 9965 6848
rect 9640 6808 9646 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 10962 6848 10968 6860
rect 9953 6811 10011 6817
rect 10152 6820 10968 6848
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9416 6752 9873 6780
rect 9861 6749 9873 6752
rect 9907 6780 9919 6783
rect 10152 6780 10180 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11054 6808 11060 6860
rect 11112 6808 11118 6860
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 12032 6820 12173 6848
rect 12032 6808 12038 6820
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 12526 6808 12532 6860
rect 12584 6808 12590 6860
rect 12710 6808 12716 6860
rect 12768 6808 12774 6860
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13188 6857 13216 6888
rect 13464 6888 13544 6916
rect 12989 6851 13047 6857
rect 12989 6848 13001 6851
rect 12952 6820 13001 6848
rect 12952 6808 12958 6820
rect 12989 6817 13001 6820
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 13173 6851 13231 6857
rect 13173 6817 13185 6851
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 13262 6808 13268 6860
rect 13320 6808 13326 6860
rect 13464 6857 13492 6888
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 15562 6876 15568 6928
rect 15620 6916 15626 6928
rect 15933 6919 15991 6925
rect 15933 6916 15945 6919
rect 15620 6888 15945 6916
rect 15620 6876 15626 6888
rect 15933 6885 15945 6888
rect 15979 6885 15991 6919
rect 15933 6879 15991 6885
rect 16114 6876 16120 6928
rect 16172 6916 16178 6928
rect 25884 6925 25912 6956
rect 25976 6956 26372 6984
rect 25869 6919 25927 6925
rect 16172 6888 16712 6916
rect 16172 6876 16178 6888
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 13630 6808 13636 6860
rect 13688 6808 13694 6860
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 13872 6820 14197 6848
rect 13872 6808 13878 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 14274 6808 14280 6860
rect 14332 6808 14338 6860
rect 15010 6808 15016 6860
rect 15068 6808 15074 6860
rect 15105 6851 15163 6857
rect 15105 6817 15117 6851
rect 15151 6817 15163 6851
rect 15105 6811 15163 6817
rect 15227 6851 15285 6857
rect 15227 6817 15239 6851
rect 15273 6848 15285 6851
rect 15470 6848 15476 6860
rect 15273 6820 15476 6848
rect 15273 6817 15285 6820
rect 15227 6811 15285 6817
rect 9907 6752 10180 6780
rect 10229 6783 10287 6789
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 6840 6684 7420 6712
rect 7466 6672 7472 6724
rect 7524 6672 7530 6724
rect 10244 6712 10272 6743
rect 10318 6740 10324 6792
rect 10376 6740 10382 6792
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 11238 6712 11244 6724
rect 7576 6684 9812 6712
rect 10244 6684 11244 6712
rect 7576 6644 7604 6684
rect 6380 6616 7604 6644
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 8849 6647 8907 6653
rect 8849 6644 8861 6647
rect 8720 6616 8861 6644
rect 8720 6604 8726 6616
rect 8849 6613 8861 6616
rect 8895 6613 8907 6647
rect 8849 6607 8907 6613
rect 9122 6604 9128 6656
rect 9180 6604 9186 6656
rect 9309 6647 9367 6653
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 9355 6616 9689 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 9784 6644 9812 6684
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 12820 6712 12848 6743
rect 13538 6740 13544 6792
rect 13596 6740 13602 6792
rect 14001 6783 14059 6789
rect 14001 6749 14013 6783
rect 14047 6780 14059 6783
rect 15120 6780 15148 6811
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15654 6808 15660 6860
rect 15712 6808 15718 6860
rect 16390 6808 16396 6860
rect 16448 6808 16454 6860
rect 16684 6857 16712 6888
rect 22112 6888 22416 6916
rect 16669 6851 16727 6857
rect 16669 6817 16681 6851
rect 16715 6848 16727 6851
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 16715 6820 17877 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 14047 6752 15148 6780
rect 15381 6783 15439 6789
rect 14047 6749 14059 6752
rect 14001 6743 14059 6749
rect 15381 6749 15393 6783
rect 15427 6780 15439 6783
rect 15746 6780 15752 6792
rect 15427 6752 15752 6780
rect 15427 6749 15439 6752
rect 15381 6743 15439 6749
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 13906 6712 13912 6724
rect 12820 6684 13912 6712
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 15856 6712 15884 6743
rect 16298 6740 16304 6792
rect 16356 6740 16362 6792
rect 16758 6740 16764 6792
rect 16816 6740 16822 6792
rect 16117 6715 16175 6721
rect 16117 6712 16129 6715
rect 15856 6684 16129 6712
rect 16117 6681 16129 6684
rect 16163 6681 16175 6715
rect 17972 6712 18000 6811
rect 18230 6808 18236 6860
rect 18288 6808 18294 6860
rect 18417 6851 18475 6857
rect 18417 6817 18429 6851
rect 18463 6848 18475 6851
rect 19622 6851 19680 6857
rect 19622 6848 19634 6851
rect 18463 6820 19634 6848
rect 18463 6817 18475 6820
rect 18417 6811 18475 6817
rect 19622 6817 19634 6820
rect 19668 6817 19680 6851
rect 19622 6811 19680 6817
rect 20349 6851 20407 6857
rect 20349 6817 20361 6851
rect 20395 6848 20407 6851
rect 20438 6848 20444 6860
rect 20395 6820 20444 6848
rect 20395 6817 20407 6820
rect 20349 6811 20407 6817
rect 20438 6808 20444 6820
rect 20496 6848 20502 6860
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 20496 6820 20637 6848
rect 20496 6808 20502 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 20714 6808 20720 6860
rect 20772 6808 20778 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20824 6820 20913 6848
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18782 6780 18788 6792
rect 18095 6752 18788 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 19889 6783 19947 6789
rect 19889 6749 19901 6783
rect 19935 6780 19947 6783
rect 20533 6783 20591 6789
rect 20533 6780 20545 6783
rect 19935 6752 20545 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 20533 6749 20545 6752
rect 20579 6749 20591 6783
rect 20533 6743 20591 6749
rect 17972 6684 18552 6712
rect 16117 6675 16175 6681
rect 10318 6644 10324 6656
rect 9784 6616 10324 6644
rect 9677 6607 9735 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 13170 6604 13176 6656
rect 13228 6604 13234 6656
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 16482 6644 16488 6656
rect 15979 6616 16488 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 18524 6653 18552 6684
rect 20438 6672 20444 6724
rect 20496 6712 20502 6724
rect 20824 6712 20852 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 21048 6820 21373 6848
rect 21048 6808 21054 6820
rect 21361 6817 21373 6820
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 21545 6851 21603 6857
rect 21545 6817 21557 6851
rect 21591 6848 21603 6851
rect 21818 6848 21824 6860
rect 21591 6820 21824 6848
rect 21591 6817 21603 6820
rect 21545 6811 21603 6817
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 21910 6808 21916 6860
rect 21968 6808 21974 6860
rect 22112 6857 22140 6888
rect 22097 6851 22155 6857
rect 22097 6817 22109 6851
rect 22143 6817 22155 6851
rect 22097 6811 22155 6817
rect 22189 6851 22247 6857
rect 22189 6817 22201 6851
rect 22235 6848 22247 6851
rect 22278 6848 22284 6860
rect 22235 6820 22284 6848
rect 22235 6817 22247 6820
rect 22189 6811 22247 6817
rect 22278 6808 22284 6820
rect 22336 6808 22342 6860
rect 22388 6848 22416 6888
rect 25869 6885 25881 6919
rect 25915 6885 25927 6919
rect 25869 6879 25927 6885
rect 22445 6851 22503 6857
rect 22445 6848 22457 6851
rect 22388 6820 22457 6848
rect 22445 6817 22457 6820
rect 22491 6817 22503 6851
rect 22445 6811 22503 6817
rect 25501 6851 25559 6857
rect 25501 6817 25513 6851
rect 25547 6817 25559 6851
rect 25501 6811 25559 6817
rect 25685 6851 25743 6857
rect 25685 6817 25697 6851
rect 25731 6817 25743 6851
rect 25685 6811 25743 6817
rect 25777 6851 25835 6857
rect 25777 6817 25789 6851
rect 25823 6848 25835 6851
rect 25976 6848 26004 6956
rect 26344 6916 26372 6956
rect 29086 6916 29092 6928
rect 25823 6820 26004 6848
rect 26099 6885 26157 6891
rect 26344 6888 26832 6916
rect 26099 6851 26111 6885
rect 26145 6882 26157 6885
rect 26145 6860 26280 6882
rect 26145 6854 26240 6860
rect 26145 6851 26157 6854
rect 26099 6845 26157 6851
rect 25823 6817 25835 6820
rect 25777 6811 25835 6817
rect 21729 6783 21787 6789
rect 21729 6749 21741 6783
rect 21775 6780 21787 6783
rect 21775 6752 21864 6780
rect 21775 6749 21787 6752
rect 21729 6743 21787 6749
rect 21836 6724 21864 6752
rect 20496 6684 20852 6712
rect 20496 6672 20502 6684
rect 21818 6672 21824 6724
rect 21876 6672 21882 6724
rect 25516 6712 25544 6811
rect 25700 6780 25728 6811
rect 26234 6808 26240 6854
rect 26292 6808 26298 6860
rect 26418 6808 26424 6860
rect 26476 6808 26482 6860
rect 26677 6851 26735 6857
rect 26677 6848 26689 6851
rect 26528 6820 26689 6848
rect 26142 6780 26148 6792
rect 25700 6752 26148 6780
rect 26142 6740 26148 6752
rect 26200 6740 26206 6792
rect 26528 6780 26556 6820
rect 26677 6817 26689 6820
rect 26723 6817 26735 6851
rect 26804 6848 26832 6888
rect 28828 6888 29092 6916
rect 26970 6848 26976 6860
rect 26804 6820 26976 6848
rect 26677 6811 26735 6817
rect 26970 6808 26976 6820
rect 27028 6848 27034 6860
rect 28074 6848 28080 6860
rect 27028 6820 28080 6848
rect 27028 6808 27034 6820
rect 28074 6808 28080 6820
rect 28132 6808 28138 6860
rect 28629 6851 28687 6857
rect 28629 6817 28641 6851
rect 28675 6848 28687 6851
rect 28828 6848 28856 6888
rect 29086 6876 29092 6888
rect 29144 6876 29150 6928
rect 28902 6857 28908 6860
rect 28675 6820 28856 6848
rect 28675 6817 28687 6820
rect 28629 6811 28687 6817
rect 28896 6811 28908 6857
rect 28960 6848 28966 6860
rect 28960 6820 28996 6848
rect 28902 6808 28908 6811
rect 28960 6808 28966 6820
rect 29270 6808 29276 6860
rect 29328 6848 29334 6860
rect 30101 6851 30159 6857
rect 30101 6848 30113 6851
rect 29328 6820 30113 6848
rect 29328 6808 29334 6820
rect 30101 6817 30113 6820
rect 30147 6817 30159 6851
rect 30101 6811 30159 6817
rect 30653 6783 30711 6789
rect 30653 6780 30665 6783
rect 26252 6752 26556 6780
rect 30024 6752 30665 6780
rect 26252 6721 26280 6752
rect 26237 6715 26295 6721
rect 25516 6684 26188 6712
rect 18509 6647 18567 6653
rect 18509 6613 18521 6647
rect 18555 6644 18567 6647
rect 18966 6644 18972 6656
rect 18555 6616 18972 6644
rect 18555 6613 18567 6616
rect 18509 6607 18567 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 20901 6647 20959 6653
rect 20901 6613 20913 6647
rect 20947 6644 20959 6647
rect 20990 6644 20996 6656
rect 20947 6616 20996 6644
rect 20947 6613 20959 6616
rect 20901 6607 20959 6613
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 22002 6644 22008 6656
rect 21600 6616 22008 6644
rect 21600 6604 21606 6616
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 23569 6647 23627 6653
rect 23569 6644 23581 6647
rect 23440 6616 23581 6644
rect 23440 6604 23446 6616
rect 23569 6613 23581 6616
rect 23615 6613 23627 6647
rect 23569 6607 23627 6613
rect 26050 6604 26056 6656
rect 26108 6604 26114 6656
rect 26160 6644 26188 6684
rect 26237 6681 26249 6715
rect 26283 6681 26295 6715
rect 26237 6675 26295 6681
rect 27522 6672 27528 6724
rect 27580 6712 27586 6724
rect 28350 6712 28356 6724
rect 27580 6684 28356 6712
rect 27580 6672 27586 6684
rect 28350 6672 28356 6684
rect 28408 6672 28414 6724
rect 30024 6656 30052 6752
rect 30653 6749 30665 6752
rect 30699 6749 30711 6783
rect 30653 6743 30711 6749
rect 26326 6644 26332 6656
rect 26160 6616 26332 6644
rect 26326 6604 26332 6616
rect 26384 6644 26390 6656
rect 27430 6644 27436 6656
rect 26384 6616 27436 6644
rect 26384 6604 26390 6616
rect 27430 6604 27436 6616
rect 27488 6644 27494 6656
rect 27801 6647 27859 6653
rect 27801 6644 27813 6647
rect 27488 6616 27813 6644
rect 27488 6604 27494 6616
rect 27801 6613 27813 6616
rect 27847 6613 27859 6647
rect 27801 6607 27859 6613
rect 28537 6647 28595 6653
rect 28537 6613 28549 6647
rect 28583 6644 28595 6647
rect 28902 6644 28908 6656
rect 28583 6616 28908 6644
rect 28583 6613 28595 6616
rect 28537 6607 28595 6613
rect 28902 6604 28908 6616
rect 28960 6604 28966 6656
rect 30006 6604 30012 6656
rect 30064 6604 30070 6656
rect 552 6554 31648 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 11436 6554
rect 11488 6502 11500 6554
rect 11552 6502 11564 6554
rect 11616 6502 11628 6554
rect 11680 6502 11692 6554
rect 11744 6502 19210 6554
rect 19262 6502 19274 6554
rect 19326 6502 19338 6554
rect 19390 6502 19402 6554
rect 19454 6502 19466 6554
rect 19518 6502 26984 6554
rect 27036 6502 27048 6554
rect 27100 6502 27112 6554
rect 27164 6502 27176 6554
rect 27228 6502 27240 6554
rect 27292 6502 31648 6554
rect 552 6480 31648 6502
rect 1946 6400 1952 6452
rect 2004 6400 2010 6452
rect 7653 6443 7711 6449
rect 7653 6409 7665 6443
rect 7699 6440 7711 6443
rect 8018 6440 8024 6452
rect 7699 6412 8024 6440
rect 7699 6409 7711 6412
rect 7653 6403 7711 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 9033 6443 9091 6449
rect 8312 6412 8984 6440
rect 3142 6372 3148 6384
rect 2976 6344 3148 6372
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2976 6304 3004 6344
rect 3142 6332 3148 6344
rect 3200 6332 3206 6384
rect 3234 6332 3240 6384
rect 3292 6332 3298 6384
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 6457 6375 6515 6381
rect 6457 6372 6469 6375
rect 6328 6344 6469 6372
rect 6328 6332 6334 6344
rect 6457 6341 6469 6344
rect 6503 6341 6515 6375
rect 6457 6335 6515 6341
rect 7558 6332 7564 6384
rect 7616 6372 7622 6384
rect 8312 6372 8340 6412
rect 7616 6344 8340 6372
rect 7616 6332 7622 6344
rect 8386 6332 8392 6384
rect 8444 6372 8450 6384
rect 8956 6372 8984 6412
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9858 6440 9864 6452
rect 9079 6412 9864 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6440 10011 6443
rect 10318 6440 10324 6452
rect 9999 6412 10324 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 15470 6400 15476 6452
rect 15528 6440 15534 6452
rect 17126 6440 17132 6452
rect 15528 6412 17132 6440
rect 15528 6400 15534 6412
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 18230 6400 18236 6452
rect 18288 6440 18294 6452
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 18288 6412 18705 6440
rect 18288 6400 18294 6412
rect 18693 6409 18705 6412
rect 18739 6409 18751 6443
rect 18693 6403 18751 6409
rect 18782 6400 18788 6452
rect 18840 6440 18846 6452
rect 21818 6440 21824 6452
rect 18840 6412 21824 6440
rect 18840 6400 18846 6412
rect 21818 6400 21824 6412
rect 21876 6400 21882 6452
rect 21910 6400 21916 6452
rect 21968 6440 21974 6452
rect 22189 6443 22247 6449
rect 22189 6440 22201 6443
rect 21968 6412 22201 6440
rect 21968 6400 21974 6412
rect 22189 6409 22201 6412
rect 22235 6409 22247 6443
rect 22189 6403 22247 6409
rect 26142 6400 26148 6452
rect 26200 6400 26206 6452
rect 26234 6400 26240 6452
rect 26292 6440 26298 6452
rect 28353 6443 28411 6449
rect 28353 6440 28365 6443
rect 26292 6412 28365 6440
rect 26292 6400 26298 6412
rect 28353 6409 28365 6412
rect 28399 6409 28411 6443
rect 28353 6403 28411 6409
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 8444 6344 8892 6372
rect 8956 6344 12173 6372
rect 8444 6332 8450 6344
rect 2910 6276 3004 6304
rect 2130 6196 2136 6248
rect 2188 6196 2194 6248
rect 2590 6196 2596 6248
rect 2648 6196 2654 6248
rect 2774 6196 2780 6248
rect 2832 6196 2838 6248
rect 2910 6245 2938 6276
rect 3050 6264 3056 6316
rect 3108 6264 3114 6316
rect 6086 6304 6092 6316
rect 3528 6276 6092 6304
rect 3528 6248 3556 6276
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6564 6276 6653 6304
rect 2910 6239 2973 6245
rect 2910 6208 2927 6239
rect 2915 6205 2927 6208
rect 2961 6205 2973 6239
rect 2915 6199 2973 6205
rect 3418 6196 3424 6248
rect 3476 6196 3482 6248
rect 3510 6196 3516 6248
rect 3568 6196 3574 6248
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4062 6236 4068 6248
rect 3927 6208 4068 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6362 6236 6368 6248
rect 6227 6208 6368 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6362 6196 6368 6208
rect 6420 6196 6426 6248
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 6564 6236 6592 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8352 6276 8585 6304
rect 8352 6264 8358 6276
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 8864 6313 8892 6344
rect 12161 6341 12173 6344
rect 12207 6372 12219 6375
rect 12207 6344 12434 6372
rect 12207 6341 12219 6344
rect 12161 6335 12219 6341
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9548 6276 9597 6304
rect 9548 6264 9554 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6304 10103 6307
rect 11238 6304 11244 6316
rect 10091 6276 11244 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 12406 6304 12434 6344
rect 12894 6332 12900 6384
rect 12952 6372 12958 6384
rect 20438 6372 20444 6384
rect 12952 6344 20444 6372
rect 12952 6332 12958 6344
rect 20438 6332 20444 6344
rect 20496 6332 20502 6384
rect 20990 6332 20996 6384
rect 21048 6372 21054 6384
rect 24854 6372 24860 6384
rect 21048 6344 24860 6372
rect 21048 6332 21054 6344
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 26160 6372 26188 6400
rect 27246 6372 27252 6384
rect 26160 6344 27252 6372
rect 27246 6332 27252 6344
rect 27304 6372 27310 6384
rect 27982 6372 27988 6384
rect 27304 6344 27988 6372
rect 27304 6332 27310 6344
rect 27982 6332 27988 6344
rect 28040 6372 28046 6384
rect 29089 6375 29147 6381
rect 29089 6372 29101 6375
rect 28040 6344 29101 6372
rect 28040 6332 28046 6344
rect 16298 6304 16304 6316
rect 12406 6276 16304 6304
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 18414 6264 18420 6316
rect 18472 6304 18478 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 18472 6276 19349 6304
rect 18472 6264 18478 6276
rect 19337 6273 19349 6276
rect 19383 6304 19395 6307
rect 19702 6304 19708 6316
rect 19383 6276 19708 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 20640 6276 25360 6304
rect 20640 6248 20668 6276
rect 6512 6208 6592 6236
rect 6512 6196 6518 6208
rect 6730 6196 6736 6248
rect 6788 6196 6794 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7561 6239 7619 6245
rect 7561 6236 7573 6239
rect 7524 6208 7573 6236
rect 7524 6196 7530 6208
rect 7561 6205 7573 6208
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 11698 6236 11704 6248
rect 10367 6208 11704 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 2682 6128 2688 6180
rect 2740 6128 2746 6180
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 3605 6171 3663 6177
rect 3605 6168 3617 6171
rect 3384 6140 3617 6168
rect 3384 6128 3390 6140
rect 3605 6137 3617 6140
rect 3651 6137 3663 6171
rect 3605 6131 3663 6137
rect 3743 6171 3801 6177
rect 3743 6137 3755 6171
rect 3789 6168 3801 6171
rect 4154 6168 4160 6180
rect 3789 6140 4160 6168
rect 3789 6137 3801 6140
rect 3743 6131 3801 6137
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 6822 6128 6828 6180
rect 6880 6128 6886 6180
rect 8772 6168 8800 6199
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12253 6239 12311 6245
rect 12253 6236 12265 6239
rect 12032 6208 12265 6236
rect 12032 6196 12038 6208
rect 12253 6205 12265 6208
rect 12299 6236 12311 6239
rect 14826 6236 14832 6248
rect 12299 6208 14832 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 18322 6196 18328 6248
rect 18380 6236 18386 6248
rect 18690 6236 18696 6248
rect 18380 6208 18696 6236
rect 18380 6196 18386 6208
rect 18690 6196 18696 6208
rect 18748 6236 18754 6248
rect 18877 6239 18935 6245
rect 18877 6236 18889 6239
rect 18748 6208 18889 6236
rect 18748 6196 18754 6208
rect 18877 6205 18889 6208
rect 18923 6205 18935 6239
rect 18877 6199 18935 6205
rect 18966 6196 18972 6248
rect 19024 6196 19030 6248
rect 20349 6239 20407 6245
rect 19076 6208 20300 6236
rect 19076 6180 19104 6208
rect 8938 6168 8944 6180
rect 8772 6140 8944 6168
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 9493 6171 9551 6177
rect 9493 6168 9505 6171
rect 9180 6140 9505 6168
rect 9180 6128 9186 6140
rect 9493 6137 9505 6140
rect 9539 6137 9551 6171
rect 9493 6131 9551 6137
rect 9677 6171 9735 6177
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 10410 6168 10416 6180
rect 9723 6140 10416 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 18506 6128 18512 6180
rect 18564 6168 18570 6180
rect 19058 6168 19064 6180
rect 18564 6140 19064 6168
rect 18564 6128 18570 6140
rect 19058 6128 19064 6140
rect 19116 6128 19122 6180
rect 19179 6171 19237 6177
rect 19179 6137 19191 6171
rect 19225 6137 19237 6171
rect 19179 6131 19237 6137
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2409 6103 2467 6109
rect 2409 6100 2421 6103
rect 2280 6072 2421 6100
rect 2280 6060 2286 6072
rect 2409 6069 2421 6072
rect 2455 6069 2467 6103
rect 2409 6063 2467 6069
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 3344 6100 3372 6128
rect 2832 6072 3372 6100
rect 2832 6060 2838 6072
rect 6546 6060 6552 6112
rect 6604 6100 6610 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 6604 6072 10241 6100
rect 6604 6060 6610 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10229 6063 10287 6069
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12802 6100 12808 6112
rect 11940 6072 12808 6100
rect 11940 6060 11946 6072
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 13078 6060 13084 6112
rect 13136 6100 13142 6112
rect 13722 6100 13728 6112
rect 13136 6072 13728 6100
rect 13136 6060 13142 6072
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 18874 6060 18880 6112
rect 18932 6100 18938 6112
rect 19194 6100 19222 6131
rect 19610 6128 19616 6180
rect 19668 6128 19674 6180
rect 20272 6168 20300 6208
rect 20349 6205 20361 6239
rect 20395 6236 20407 6239
rect 20622 6236 20628 6248
rect 20395 6208 20628 6236
rect 20395 6205 20407 6208
rect 20349 6199 20407 6205
rect 20622 6196 20628 6208
rect 20680 6196 20686 6248
rect 21082 6196 21088 6248
rect 21140 6236 21146 6248
rect 21726 6245 21732 6248
rect 21545 6239 21603 6245
rect 21545 6236 21557 6239
rect 21140 6208 21557 6236
rect 21140 6196 21146 6208
rect 21545 6205 21557 6208
rect 21591 6205 21603 6239
rect 21545 6199 21603 6205
rect 21703 6239 21732 6245
rect 21703 6205 21715 6239
rect 21703 6199 21732 6205
rect 21726 6196 21732 6199
rect 21784 6196 21790 6248
rect 22002 6196 22008 6248
rect 22060 6236 22066 6248
rect 22462 6236 22468 6248
rect 22060 6208 22468 6236
rect 22060 6196 22066 6208
rect 22462 6196 22468 6208
rect 22520 6196 22526 6248
rect 23658 6196 23664 6248
rect 23716 6236 23722 6248
rect 24673 6239 24731 6245
rect 24673 6236 24685 6239
rect 23716 6208 24685 6236
rect 23716 6196 23722 6208
rect 24673 6205 24685 6208
rect 24719 6205 24731 6239
rect 24673 6199 24731 6205
rect 21450 6168 21456 6180
rect 20272 6140 21456 6168
rect 21450 6128 21456 6140
rect 21508 6168 21514 6180
rect 21821 6171 21879 6177
rect 21821 6168 21833 6171
rect 21508 6140 21833 6168
rect 21508 6128 21514 6140
rect 21821 6137 21833 6140
rect 21867 6137 21879 6171
rect 21821 6131 21879 6137
rect 21913 6171 21971 6177
rect 21913 6137 21925 6171
rect 21959 6168 21971 6171
rect 22278 6168 22284 6180
rect 21959 6140 22284 6168
rect 21959 6137 21971 6140
rect 21913 6131 21971 6137
rect 22278 6128 22284 6140
rect 22336 6168 22342 6180
rect 23382 6168 23388 6180
rect 22336 6140 23388 6168
rect 22336 6128 22342 6140
rect 23382 6128 23388 6140
rect 23440 6128 23446 6180
rect 18932 6072 19222 6100
rect 24688 6100 24716 6199
rect 24946 6196 24952 6248
rect 25004 6196 25010 6248
rect 25041 6239 25099 6245
rect 25041 6205 25053 6239
rect 25087 6236 25099 6239
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25087 6208 25237 6236
rect 25087 6205 25099 6208
rect 25041 6199 25099 6205
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25332 6236 25360 6276
rect 27430 6264 27436 6316
rect 27488 6264 27494 6316
rect 27522 6264 27528 6316
rect 27580 6304 27586 6316
rect 28169 6307 28227 6313
rect 28169 6304 28181 6307
rect 27580 6276 28181 6304
rect 27580 6264 27586 6276
rect 28169 6273 28181 6276
rect 28215 6273 28227 6307
rect 28169 6267 28227 6273
rect 26418 6236 26424 6248
rect 25332 6208 26424 6236
rect 25225 6199 25283 6205
rect 26418 6196 26424 6208
rect 26476 6236 26482 6248
rect 26697 6239 26755 6245
rect 26697 6236 26709 6239
rect 26476 6208 26709 6236
rect 26476 6196 26482 6208
rect 26697 6205 26709 6208
rect 26743 6205 26755 6239
rect 27448 6236 27476 6264
rect 27893 6239 27951 6245
rect 27893 6236 27905 6239
rect 27448 6208 27905 6236
rect 26697 6199 26755 6205
rect 27893 6205 27905 6208
rect 27939 6205 27951 6239
rect 27893 6199 27951 6205
rect 25492 6171 25550 6177
rect 25492 6137 25504 6171
rect 25538 6168 25550 6171
rect 25590 6168 25596 6180
rect 25538 6140 25596 6168
rect 25538 6137 25550 6140
rect 25492 6131 25550 6137
rect 25590 6128 25596 6140
rect 25648 6128 25654 6180
rect 27430 6168 27436 6180
rect 26252 6140 27436 6168
rect 26252 6100 26280 6140
rect 27430 6128 27436 6140
rect 27488 6128 27494 6180
rect 27908 6168 27936 6199
rect 27982 6196 27988 6248
rect 28040 6196 28046 6248
rect 28074 6196 28080 6248
rect 28132 6196 28138 6248
rect 28828 6245 28856 6344
rect 29089 6341 29101 6344
rect 29135 6341 29147 6375
rect 29089 6335 29147 6341
rect 28537 6239 28595 6245
rect 28537 6205 28549 6239
rect 28583 6205 28595 6239
rect 28537 6199 28595 6205
rect 28813 6239 28871 6245
rect 28813 6205 28825 6239
rect 28859 6205 28871 6239
rect 28813 6199 28871 6205
rect 28552 6168 28580 6199
rect 30466 6196 30472 6248
rect 30524 6196 30530 6248
rect 27908 6140 28580 6168
rect 29914 6128 29920 6180
rect 29972 6168 29978 6180
rect 30202 6171 30260 6177
rect 30202 6168 30214 6171
rect 29972 6140 30214 6168
rect 29972 6128 29978 6140
rect 30202 6137 30214 6140
rect 30248 6137 30260 6171
rect 30202 6131 30260 6137
rect 24688 6072 26280 6100
rect 18932 6060 18938 6072
rect 26326 6060 26332 6112
rect 26384 6100 26390 6112
rect 26605 6103 26663 6109
rect 26605 6100 26617 6103
rect 26384 6072 26617 6100
rect 26384 6060 26390 6072
rect 26605 6069 26617 6072
rect 26651 6069 26663 6103
rect 26605 6063 26663 6069
rect 26694 6060 26700 6112
rect 26752 6100 26758 6112
rect 27709 6103 27767 6109
rect 27709 6100 27721 6103
rect 26752 6072 27721 6100
rect 26752 6060 26758 6072
rect 27709 6069 27721 6072
rect 27755 6069 27767 6103
rect 27709 6063 27767 6069
rect 28074 6060 28080 6112
rect 28132 6100 28138 6112
rect 28721 6103 28779 6109
rect 28721 6100 28733 6103
rect 28132 6072 28733 6100
rect 28132 6060 28138 6072
rect 28721 6069 28733 6072
rect 28767 6100 28779 6103
rect 30006 6100 30012 6112
rect 28767 6072 30012 6100
rect 28767 6069 28779 6072
rect 28721 6063 28779 6069
rect 30006 6060 30012 6072
rect 30064 6060 30070 6112
rect 552 6010 31648 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 12096 6010
rect 12148 5958 12160 6010
rect 12212 5958 12224 6010
rect 12276 5958 12288 6010
rect 12340 5958 12352 6010
rect 12404 5958 19870 6010
rect 19922 5958 19934 6010
rect 19986 5958 19998 6010
rect 20050 5958 20062 6010
rect 20114 5958 20126 6010
rect 20178 5958 27644 6010
rect 27696 5958 27708 6010
rect 27760 5958 27772 6010
rect 27824 5958 27836 6010
rect 27888 5958 27900 6010
rect 27952 5958 31648 6010
rect 552 5936 31648 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 2866 5896 2872 5908
rect 2823 5868 2872 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8996 5868 9045 5896
rect 8996 5856 9002 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 12437 5899 12495 5905
rect 11756 5868 12112 5896
rect 11756 5856 11762 5868
rect 1964 5800 3464 5828
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1964 5769 1992 5800
rect 1949 5763 2007 5769
rect 1949 5760 1961 5763
rect 1452 5732 1961 5760
rect 1452 5720 1458 5732
rect 1949 5729 1961 5732
rect 1995 5729 2007 5763
rect 1949 5723 2007 5729
rect 2222 5720 2228 5772
rect 2280 5720 2286 5772
rect 2314 5720 2320 5772
rect 2372 5760 2378 5772
rect 2372 5732 2774 5760
rect 2372 5720 2378 5732
rect 2746 5692 2774 5732
rect 2958 5720 2964 5772
rect 3016 5720 3022 5772
rect 3436 5769 3464 5800
rect 8294 5788 8300 5840
rect 8352 5828 8358 5840
rect 8665 5831 8723 5837
rect 8665 5828 8677 5831
rect 8352 5800 8677 5828
rect 8352 5788 8358 5800
rect 8665 5797 8677 5800
rect 8711 5797 8723 5831
rect 8665 5791 8723 5797
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 9125 5831 9183 5837
rect 9125 5828 9137 5831
rect 8803 5800 9137 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 9125 5797 9137 5800
rect 9171 5797 9183 5831
rect 9125 5791 9183 5797
rect 9398 5788 9404 5840
rect 9456 5828 9462 5840
rect 9493 5831 9551 5837
rect 9493 5828 9505 5831
rect 9456 5800 9505 5828
rect 9456 5788 9462 5800
rect 9493 5797 9505 5800
rect 9539 5828 9551 5831
rect 11425 5831 11483 5837
rect 9539 5800 9812 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 4154 5760 4160 5772
rect 3467 5732 4160 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 8386 5720 8392 5772
rect 8444 5720 8450 5772
rect 8478 5720 8484 5772
rect 8536 5720 8542 5772
rect 8895 5763 8953 5769
rect 8895 5729 8907 5763
rect 8941 5760 8953 5763
rect 9309 5763 9367 5769
rect 8941 5732 9260 5760
rect 8941 5729 8953 5732
rect 8895 5723 8953 5729
rect 3145 5695 3203 5701
rect 3145 5692 3157 5695
rect 2746 5664 3157 5692
rect 3145 5661 3157 5664
rect 3191 5661 3203 5695
rect 9232 5692 9260 5732
rect 9309 5729 9321 5763
rect 9355 5760 9367 5763
rect 9582 5760 9588 5772
rect 9355 5732 9588 5760
rect 9355 5729 9367 5732
rect 9309 5723 9367 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9784 5769 9812 5800
rect 11425 5797 11437 5831
rect 11471 5828 11483 5831
rect 11790 5828 11796 5840
rect 11471 5800 11796 5828
rect 11471 5797 11483 5800
rect 11425 5791 11483 5797
rect 11790 5788 11796 5800
rect 11848 5828 11854 5840
rect 11848 5800 12020 5828
rect 11848 5788 11854 5800
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5760 11391 5763
rect 11379 5732 11468 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9232 5664 9689 5692
rect 3145 5655 3203 5661
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 6178 5624 6184 5636
rect 2832 5596 6184 5624
rect 2832 5584 2838 5596
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 9950 5624 9956 5636
rect 8628 5596 9956 5624
rect 8628 5584 8634 5596
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 1670 5516 1676 5568
rect 1728 5556 1734 5568
rect 1857 5559 1915 5565
rect 1857 5556 1869 5559
rect 1728 5528 1869 5556
rect 1728 5516 1734 5528
rect 1857 5525 1869 5528
rect 1903 5525 1915 5559
rect 1857 5519 1915 5525
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 2004 5528 2053 5556
rect 2004 5516 2010 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3329 5559 3387 5565
rect 3329 5556 3341 5559
rect 3200 5528 3341 5556
rect 3200 5516 3206 5528
rect 3329 5525 3341 5528
rect 3375 5525 3387 5559
rect 3329 5519 3387 5525
rect 11146 5516 11152 5568
rect 11204 5516 11210 5568
rect 11440 5556 11468 5732
rect 11514 5720 11520 5772
rect 11572 5720 11578 5772
rect 11655 5763 11713 5769
rect 11655 5729 11667 5763
rect 11701 5760 11713 5763
rect 11882 5760 11888 5772
rect 11701 5732 11888 5760
rect 11701 5729 11713 5732
rect 11655 5723 11713 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 11992 5701 12020 5800
rect 12084 5769 12112 5868
rect 12437 5865 12449 5899
rect 12483 5896 12495 5899
rect 13262 5896 13268 5908
rect 12483 5868 13268 5896
rect 12483 5865 12495 5868
rect 12437 5859 12495 5865
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 14737 5899 14795 5905
rect 13556 5868 14688 5896
rect 13556 5828 13584 5868
rect 13843 5831 13901 5837
rect 13843 5828 13855 5831
rect 13004 5800 13584 5828
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11624 5664 11805 5692
rect 11624 5636 11652 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 11606 5584 11612 5636
rect 11664 5584 11670 5636
rect 11882 5584 11888 5636
rect 11940 5624 11946 5636
rect 12084 5624 12112 5723
rect 12158 5720 12164 5772
rect 12216 5760 12222 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12216 5732 12909 5760
rect 12216 5720 12222 5732
rect 12897 5729 12909 5732
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 13004 5701 13032 5800
rect 13832 5797 13855 5828
rect 13889 5797 13901 5831
rect 14660 5828 14688 5868
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 15654 5896 15660 5908
rect 14783 5868 15660 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 22370 5896 22376 5908
rect 15804 5868 22376 5896
rect 15804 5856 15810 5868
rect 22370 5856 22376 5868
rect 22428 5896 22434 5908
rect 23382 5896 23388 5908
rect 22428 5868 23388 5896
rect 22428 5856 22434 5868
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 25590 5856 25596 5908
rect 25648 5856 25654 5908
rect 25777 5899 25835 5905
rect 25777 5865 25789 5899
rect 25823 5896 25835 5899
rect 26694 5896 26700 5908
rect 25823 5868 26700 5896
rect 25823 5865 25835 5868
rect 25777 5859 25835 5865
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 27801 5899 27859 5905
rect 27801 5865 27813 5899
rect 27847 5896 27859 5899
rect 27982 5896 27988 5908
rect 27847 5868 27988 5896
rect 27847 5865 27859 5868
rect 27801 5859 27859 5865
rect 27982 5856 27988 5868
rect 28040 5856 28046 5908
rect 29003 5899 29061 5905
rect 29003 5865 29015 5899
rect 29049 5896 29061 5899
rect 29049 5868 29408 5896
rect 29049 5865 29061 5868
rect 29003 5859 29061 5865
rect 17954 5828 17960 5840
rect 14660 5800 17960 5828
rect 13832 5791 13901 5797
rect 13538 5720 13544 5772
rect 13596 5720 13602 5772
rect 13630 5720 13636 5772
rect 13688 5720 13694 5772
rect 13722 5720 13728 5772
rect 13780 5720 13786 5772
rect 13832 5704 13860 5791
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 18690 5788 18696 5840
rect 18748 5788 18754 5840
rect 18785 5831 18843 5837
rect 18785 5797 18797 5831
rect 18831 5828 18843 5831
rect 19058 5828 19064 5840
rect 18831 5800 19064 5828
rect 18831 5797 18843 5800
rect 18785 5791 18843 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 26418 5788 26424 5840
rect 26476 5788 26482 5840
rect 27249 5831 27307 5837
rect 27249 5797 27261 5831
rect 27295 5828 27307 5831
rect 27338 5828 27344 5840
rect 27295 5800 27344 5828
rect 27295 5797 27307 5800
rect 27249 5791 27307 5797
rect 13998 5720 14004 5772
rect 14056 5720 14062 5772
rect 14090 5720 14096 5772
rect 14148 5720 14154 5772
rect 14231 5763 14289 5769
rect 14231 5729 14243 5763
rect 14277 5729 14289 5763
rect 14231 5723 14289 5729
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5661 13047 5695
rect 13814 5692 13820 5704
rect 12989 5655 13047 5661
rect 13189 5664 13820 5692
rect 11940 5596 12112 5624
rect 11940 5584 11946 5596
rect 12802 5584 12808 5636
rect 12860 5624 12866 5636
rect 13189 5624 13217 5664
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14256 5692 14284 5723
rect 14366 5720 14372 5772
rect 14424 5720 14430 5772
rect 14458 5720 14464 5772
rect 14516 5720 14522 5772
rect 14550 5720 14556 5772
rect 14608 5769 14614 5772
rect 14608 5760 14616 5769
rect 14608 5732 14653 5760
rect 14608 5723 14616 5732
rect 14608 5720 14614 5723
rect 14826 5720 14832 5772
rect 14884 5720 14890 5772
rect 14983 5763 15041 5769
rect 14983 5729 14995 5763
rect 15029 5760 15041 5763
rect 16390 5760 16396 5772
rect 15029 5732 16396 5760
rect 15029 5729 15041 5732
rect 14983 5723 15041 5729
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18601 5766 18659 5769
rect 18524 5763 18659 5766
rect 18524 5760 18613 5763
rect 18380 5738 18613 5760
rect 18380 5732 18552 5738
rect 18380 5720 18386 5732
rect 18601 5729 18613 5738
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18874 5720 18880 5772
rect 18932 5769 18938 5772
rect 18932 5763 18961 5769
rect 18949 5729 18961 5763
rect 18932 5723 18961 5729
rect 18932 5720 18938 5723
rect 19610 5720 19616 5772
rect 19668 5760 19674 5772
rect 21545 5763 21603 5769
rect 21545 5760 21557 5763
rect 19668 5732 21557 5760
rect 19668 5720 19674 5732
rect 21545 5729 21557 5732
rect 21591 5729 21603 5763
rect 21910 5760 21916 5772
rect 21545 5723 21603 5729
rect 21652 5732 21916 5760
rect 14642 5692 14648 5704
rect 14256 5664 14648 5692
rect 14642 5652 14648 5664
rect 14700 5652 14706 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5692 19119 5695
rect 21652 5692 21680 5732
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 22646 5720 22652 5772
rect 22704 5720 22710 5772
rect 22738 5720 22744 5772
rect 22796 5760 22802 5772
rect 23109 5763 23167 5769
rect 23109 5760 23121 5763
rect 22796 5732 23121 5760
rect 22796 5720 22802 5732
rect 23109 5729 23121 5732
rect 23155 5729 23167 5763
rect 23109 5723 23167 5729
rect 24946 5720 24952 5772
rect 25004 5760 25010 5772
rect 25317 5763 25375 5769
rect 25317 5760 25329 5763
rect 25004 5732 25329 5760
rect 25004 5720 25010 5732
rect 25317 5729 25329 5732
rect 25363 5760 25375 5763
rect 27264 5760 27292 5791
rect 27338 5788 27344 5800
rect 27396 5788 27402 5840
rect 28000 5828 28028 5856
rect 28813 5831 28871 5837
rect 28000 5800 28672 5828
rect 25363 5732 27292 5760
rect 27617 5763 27675 5769
rect 25363 5729 25375 5732
rect 25317 5723 25375 5729
rect 27617 5729 27629 5763
rect 27663 5729 27675 5763
rect 27617 5723 27675 5729
rect 27709 5763 27767 5769
rect 27709 5729 27721 5763
rect 27755 5729 27767 5763
rect 27709 5723 27767 5729
rect 27985 5763 28043 5769
rect 27985 5729 27997 5763
rect 28031 5760 28043 5763
rect 28074 5760 28080 5772
rect 28031 5732 28080 5760
rect 28031 5729 28043 5732
rect 27985 5723 28043 5729
rect 19107 5664 21680 5692
rect 19107 5661 19119 5664
rect 19061 5655 19119 5661
rect 12860 5596 13217 5624
rect 13265 5627 13323 5633
rect 12860 5584 12866 5596
rect 13265 5593 13277 5627
rect 13311 5624 13323 5627
rect 14090 5624 14096 5636
rect 13311 5596 14096 5624
rect 13311 5593 13323 5596
rect 13265 5587 13323 5593
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 19076 5624 19104 5655
rect 21818 5652 21824 5704
rect 21876 5692 21882 5704
rect 22465 5695 22523 5701
rect 22465 5692 22477 5695
rect 21876 5664 22477 5692
rect 21876 5652 21882 5664
rect 22465 5661 22477 5664
rect 22511 5692 22523 5695
rect 22925 5695 22983 5701
rect 22925 5692 22937 5695
rect 22511 5664 22937 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 22925 5661 22937 5664
rect 22971 5661 22983 5695
rect 22925 5655 22983 5661
rect 26326 5652 26332 5704
rect 26384 5692 26390 5704
rect 27522 5692 27528 5704
rect 26384 5664 27528 5692
rect 26384 5652 26390 5664
rect 27522 5652 27528 5664
rect 27580 5692 27586 5704
rect 27632 5692 27660 5723
rect 27580 5664 27660 5692
rect 27580 5652 27586 5664
rect 14844 5596 19104 5624
rect 12894 5556 12900 5568
rect 11440 5528 12900 5556
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13354 5516 13360 5568
rect 13412 5516 13418 5568
rect 13446 5516 13452 5568
rect 13504 5556 13510 5568
rect 14844 5556 14872 5596
rect 19702 5584 19708 5636
rect 19760 5624 19766 5636
rect 26145 5627 26203 5633
rect 19760 5596 21680 5624
rect 19760 5584 19766 5596
rect 13504 5528 14872 5556
rect 13504 5516 13510 5528
rect 14918 5516 14924 5568
rect 14976 5556 14982 5568
rect 15013 5559 15071 5565
rect 15013 5556 15025 5559
rect 14976 5528 15025 5556
rect 14976 5516 14982 5528
rect 15013 5525 15025 5528
rect 15059 5525 15071 5559
rect 15013 5519 15071 5525
rect 18322 5516 18328 5568
rect 18380 5556 18386 5568
rect 18417 5559 18475 5565
rect 18417 5556 18429 5559
rect 18380 5528 18429 5556
rect 18380 5516 18386 5528
rect 18417 5525 18429 5528
rect 18463 5525 18475 5559
rect 18417 5519 18475 5525
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 18690 5556 18696 5568
rect 18564 5528 18696 5556
rect 18564 5516 18570 5528
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 21266 5516 21272 5568
rect 21324 5556 21330 5568
rect 21453 5559 21511 5565
rect 21453 5556 21465 5559
rect 21324 5528 21465 5556
rect 21324 5516 21330 5528
rect 21453 5525 21465 5528
rect 21499 5525 21511 5559
rect 21652 5556 21680 5596
rect 26145 5593 26157 5627
rect 26191 5593 26203 5627
rect 26145 5587 26203 5593
rect 22002 5556 22008 5568
rect 21652 5528 22008 5556
rect 21453 5519 21511 5525
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 22833 5559 22891 5565
rect 22833 5525 22845 5559
rect 22879 5556 22891 5559
rect 23106 5556 23112 5568
rect 22879 5528 23112 5556
rect 22879 5525 22891 5528
rect 22833 5519 22891 5525
rect 23106 5516 23112 5528
rect 23164 5516 23170 5568
rect 23293 5559 23351 5565
rect 23293 5525 23305 5559
rect 23339 5556 23351 5559
rect 23934 5556 23940 5568
rect 23339 5528 23940 5556
rect 23339 5525 23351 5528
rect 23293 5519 23351 5525
rect 23934 5516 23940 5528
rect 23992 5516 23998 5568
rect 25777 5559 25835 5565
rect 25777 5525 25789 5559
rect 25823 5556 25835 5559
rect 26050 5556 26056 5568
rect 25823 5528 26056 5556
rect 25823 5525 25835 5528
rect 25777 5519 25835 5525
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 26160 5556 26188 5587
rect 26234 5584 26240 5636
rect 26292 5624 26298 5636
rect 27724 5624 27752 5723
rect 28074 5720 28080 5732
rect 28132 5760 28138 5772
rect 28644 5769 28672 5800
rect 28813 5797 28825 5831
rect 28859 5828 28871 5831
rect 28905 5831 28963 5837
rect 28905 5828 28917 5831
rect 28859 5800 28917 5828
rect 28859 5797 28871 5800
rect 28813 5791 28871 5797
rect 28905 5797 28917 5800
rect 28951 5797 28963 5831
rect 28905 5791 28963 5797
rect 29089 5831 29147 5837
rect 29089 5797 29101 5831
rect 29135 5828 29147 5831
rect 29270 5828 29276 5840
rect 29135 5800 29276 5828
rect 29135 5797 29147 5800
rect 29089 5791 29147 5797
rect 29270 5788 29276 5800
rect 29328 5788 29334 5840
rect 29380 5769 29408 5868
rect 29914 5856 29920 5908
rect 29972 5856 29978 5908
rect 30466 5856 30472 5908
rect 30524 5856 30530 5908
rect 28537 5763 28595 5769
rect 28537 5760 28549 5763
rect 28132 5732 28549 5760
rect 28132 5720 28138 5732
rect 28537 5729 28549 5732
rect 28583 5729 28595 5763
rect 28537 5723 28595 5729
rect 28629 5763 28687 5769
rect 28629 5729 28641 5763
rect 28675 5760 28687 5763
rect 29181 5763 29239 5769
rect 29181 5760 29193 5763
rect 28675 5732 29193 5760
rect 28675 5729 28687 5732
rect 28629 5723 28687 5729
rect 29181 5729 29193 5732
rect 29227 5729 29239 5763
rect 29181 5723 29239 5729
rect 29365 5763 29423 5769
rect 29365 5729 29377 5763
rect 29411 5729 29423 5763
rect 29365 5723 29423 5729
rect 30285 5763 30343 5769
rect 30285 5729 30297 5763
rect 30331 5729 30343 5763
rect 30285 5723 30343 5729
rect 28350 5652 28356 5704
rect 28408 5692 28414 5704
rect 28813 5695 28871 5701
rect 28813 5692 28825 5695
rect 28408 5664 28825 5692
rect 28408 5652 28414 5664
rect 28813 5661 28825 5664
rect 28859 5692 28871 5695
rect 29086 5692 29092 5704
rect 28859 5664 29092 5692
rect 28859 5661 28871 5664
rect 28813 5655 28871 5661
rect 29086 5652 29092 5664
rect 29144 5692 29150 5704
rect 30009 5695 30067 5701
rect 30009 5692 30021 5695
rect 29144 5664 30021 5692
rect 29144 5652 29150 5664
rect 30009 5661 30021 5664
rect 30055 5661 30067 5695
rect 30300 5692 30328 5723
rect 30374 5720 30380 5772
rect 30432 5720 30438 5772
rect 30466 5692 30472 5704
rect 30300 5664 30472 5692
rect 30009 5655 30067 5661
rect 30466 5652 30472 5664
rect 30524 5652 30530 5704
rect 26292 5596 27752 5624
rect 30101 5627 30159 5633
rect 26292 5584 26298 5596
rect 30101 5593 30113 5627
rect 30147 5624 30159 5627
rect 30650 5624 30656 5636
rect 30147 5596 30656 5624
rect 30147 5593 30159 5596
rect 30101 5587 30159 5593
rect 30650 5584 30656 5596
rect 30708 5584 30714 5636
rect 27433 5559 27491 5565
rect 27433 5556 27445 5559
rect 26160 5528 27445 5556
rect 27433 5525 27445 5528
rect 27479 5556 27491 5559
rect 28074 5556 28080 5568
rect 27479 5528 28080 5556
rect 27479 5525 27491 5528
rect 27433 5519 27491 5525
rect 28074 5516 28080 5528
rect 28132 5556 28138 5568
rect 29638 5556 29644 5568
rect 28132 5528 29644 5556
rect 28132 5516 28138 5528
rect 29638 5516 29644 5528
rect 29696 5556 29702 5568
rect 30193 5559 30251 5565
rect 30193 5556 30205 5559
rect 29696 5528 30205 5556
rect 29696 5516 29702 5528
rect 30193 5525 30205 5528
rect 30239 5525 30251 5559
rect 30193 5519 30251 5525
rect 552 5466 31648 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 11436 5466
rect 11488 5414 11500 5466
rect 11552 5414 11564 5466
rect 11616 5414 11628 5466
rect 11680 5414 11692 5466
rect 11744 5414 19210 5466
rect 19262 5414 19274 5466
rect 19326 5414 19338 5466
rect 19390 5414 19402 5466
rect 19454 5414 19466 5466
rect 19518 5414 26984 5466
rect 27036 5414 27048 5466
rect 27100 5414 27112 5466
rect 27164 5414 27176 5466
rect 27228 5414 27240 5466
rect 27292 5414 31648 5466
rect 552 5392 31648 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 2832 5324 3065 5352
rect 2832 5312 2838 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 4062 5352 4068 5364
rect 3559 5324 4068 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 5166 5352 5172 5364
rect 4203 5324 5172 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 8113 5355 8171 5361
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 8294 5352 8300 5364
rect 8159 5324 8300 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 8386 5312 8392 5364
rect 8444 5312 8450 5364
rect 11146 5352 11152 5364
rect 10336 5324 11152 5352
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 3881 5287 3939 5293
rect 3881 5284 3893 5287
rect 3660 5256 3893 5284
rect 3660 5244 3666 5256
rect 3881 5253 3893 5256
rect 3927 5284 3939 5287
rect 3973 5287 4031 5293
rect 3973 5284 3985 5287
rect 3927 5256 3985 5284
rect 3927 5253 3939 5256
rect 3881 5247 3939 5253
rect 3973 5253 3985 5256
rect 4019 5253 4031 5287
rect 3973 5247 4031 5253
rect 7561 5287 7619 5293
rect 7561 5253 7573 5287
rect 7607 5284 7619 5287
rect 8478 5284 8484 5296
rect 7607 5256 8484 5284
rect 7607 5253 7619 5256
rect 7561 5247 7619 5253
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 8588 5256 9352 5284
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 8588 5216 8616 5256
rect 7432 5188 8616 5216
rect 7432 5176 7438 5188
rect 8846 5176 8852 5228
rect 8904 5176 8910 5228
rect 1394 5108 1400 5160
rect 1452 5108 1458 5160
rect 1946 5157 1952 5160
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 1673 5151 1731 5157
rect 1673 5148 1685 5151
rect 1535 5120 1685 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 1673 5117 1685 5120
rect 1719 5117 1731 5151
rect 1940 5148 1952 5157
rect 1907 5120 1952 5148
rect 1673 5111 1731 5117
rect 1940 5111 1952 5120
rect 1946 5108 1952 5111
rect 2004 5108 2010 5160
rect 6178 5108 6184 5160
rect 6236 5148 6242 5160
rect 9324 5157 9352 5256
rect 7469 5151 7527 5157
rect 7469 5148 7481 5151
rect 6236 5120 7481 5148
rect 6236 5108 6242 5120
rect 7469 5117 7481 5120
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 8757 5151 8815 5157
rect 7699 5120 7880 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 4246 5040 4252 5092
rect 4304 5080 4310 5092
rect 4341 5083 4399 5089
rect 4341 5080 4353 5083
rect 4304 5052 4353 5080
rect 4304 5040 4310 5052
rect 4341 5049 4353 5052
rect 4387 5049 4399 5083
rect 7484 5080 7512 5111
rect 7852 5092 7880 5120
rect 8757 5117 8769 5151
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 7484 5052 7757 5080
rect 4341 5043 4399 5049
rect 7745 5049 7757 5052
rect 7791 5049 7803 5083
rect 7745 5043 7803 5049
rect 7834 5040 7840 5092
rect 7892 5080 7898 5092
rect 7929 5083 7987 5089
rect 7929 5080 7941 5083
rect 7892 5052 7941 5080
rect 7892 5040 7898 5052
rect 7929 5049 7941 5052
rect 7975 5049 7987 5083
rect 8772 5080 8800 5111
rect 10042 5108 10048 5160
rect 10100 5108 10106 5160
rect 10137 5151 10195 5157
rect 10137 5117 10149 5151
rect 10183 5148 10195 5151
rect 10336 5148 10364 5324
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11790 5312 11796 5364
rect 11848 5312 11854 5364
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 13630 5352 13636 5364
rect 12759 5324 13636 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 14185 5355 14243 5361
rect 14185 5321 14197 5355
rect 14231 5352 14243 5355
rect 15010 5352 15016 5364
rect 14231 5324 15016 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 17126 5312 17132 5364
rect 17184 5312 17190 5364
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 18506 5352 18512 5364
rect 18104 5324 18512 5352
rect 18104 5312 18110 5324
rect 18506 5312 18512 5324
rect 18564 5352 18570 5364
rect 20073 5355 20131 5361
rect 20073 5352 20085 5355
rect 18564 5324 20085 5352
rect 18564 5312 18570 5324
rect 20073 5321 20085 5324
rect 20119 5321 20131 5355
rect 20073 5315 20131 5321
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 21508 5324 22324 5352
rect 21508 5312 21514 5324
rect 14366 5284 14372 5296
rect 13096 5256 14372 5284
rect 13096 5216 13124 5256
rect 14366 5244 14372 5256
rect 14424 5284 14430 5296
rect 18690 5284 18696 5296
rect 14424 5256 14780 5284
rect 14424 5244 14430 5256
rect 13004 5188 13124 5216
rect 10183 5120 10364 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 10410 5108 10416 5160
rect 10468 5108 10474 5160
rect 12894 5108 12900 5160
rect 12952 5108 12958 5160
rect 13004 5157 13032 5188
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 13357 5219 13415 5225
rect 13357 5216 13369 5219
rect 13320 5188 13369 5216
rect 13320 5176 13326 5188
rect 13357 5185 13369 5188
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 14550 5216 14556 5228
rect 13832 5188 14556 5216
rect 12989 5151 13047 5157
rect 12989 5117 13001 5151
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13078 5108 13084 5160
rect 13136 5108 13142 5160
rect 13538 5108 13544 5160
rect 13596 5108 13602 5160
rect 13648 5148 13676 5176
rect 13832 5160 13860 5188
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 14752 5160 14780 5256
rect 18156 5256 18696 5284
rect 18156 5225 18184 5256
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 21818 5284 21824 5296
rect 20824 5256 21824 5284
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 18141 5219 18199 5225
rect 16347 5188 18092 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 13725 5151 13783 5157
rect 13725 5148 13737 5151
rect 13648 5120 13737 5148
rect 13725 5117 13737 5120
rect 13771 5117 13783 5151
rect 13725 5111 13783 5117
rect 13814 5108 13820 5160
rect 13872 5108 13878 5160
rect 14369 5151 14427 5157
rect 14369 5117 14381 5151
rect 14415 5148 14427 5151
rect 14458 5148 14464 5160
rect 14415 5120 14464 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 9858 5080 9864 5092
rect 8772 5052 9864 5080
rect 7929 5043 7987 5049
rect 9858 5040 9864 5052
rect 9916 5040 9922 5092
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5080 10379 5083
rect 10658 5083 10716 5089
rect 10658 5080 10670 5083
rect 10367 5052 10670 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 10658 5049 10670 5052
rect 10704 5049 10716 5083
rect 10658 5043 10716 5049
rect 11716 5052 12434 5080
rect 3329 5015 3387 5021
rect 3329 4981 3341 5015
rect 3375 5012 3387 5015
rect 3418 5012 3424 5024
rect 3375 4984 3424 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 3510 4972 3516 5024
rect 3568 4972 3574 5024
rect 4141 5015 4199 5021
rect 4141 4981 4153 5015
rect 4187 5012 4199 5015
rect 5074 5012 5080 5024
rect 4187 4984 5080 5012
rect 4187 4981 4199 4984
rect 4141 4975 4199 4981
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 5012 9459 5015
rect 11716 5012 11744 5052
rect 9447 4984 11744 5012
rect 12406 5012 12434 5052
rect 12802 5040 12808 5092
rect 12860 5080 12866 5092
rect 13219 5083 13277 5089
rect 13219 5080 13231 5083
rect 12860 5052 13231 5080
rect 12860 5040 12866 5052
rect 13219 5049 13231 5052
rect 13265 5049 13277 5083
rect 14384 5080 14412 5111
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 14642 5108 14648 5160
rect 14700 5108 14706 5160
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 14918 5108 14924 5160
rect 14976 5108 14982 5160
rect 15010 5108 15016 5160
rect 15068 5108 15074 5160
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15252 5120 15853 5148
rect 15252 5108 15258 5120
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 15841 5111 15899 5117
rect 16114 5108 16120 5160
rect 16172 5157 16178 5160
rect 16172 5151 16201 5157
rect 16189 5117 16201 5151
rect 16172 5111 16201 5117
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5117 16635 5151
rect 16577 5111 16635 5117
rect 16172 5108 16178 5111
rect 13219 5043 13277 5049
rect 13740 5052 14412 5080
rect 13740 5012 13768 5052
rect 15930 5040 15936 5092
rect 15988 5040 15994 5092
rect 16025 5083 16083 5089
rect 16025 5049 16037 5083
rect 16071 5049 16083 5083
rect 16025 5043 16083 5049
rect 12406 4984 13768 5012
rect 9447 4981 9459 4984
rect 9401 4975 9459 4981
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 13872 4984 13921 5012
rect 13872 4972 13878 4984
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 13909 4975 13967 4981
rect 14918 4972 14924 5024
rect 14976 5012 14982 5024
rect 15105 5015 15163 5021
rect 15105 5012 15117 5015
rect 14976 4984 15117 5012
rect 14976 4972 14982 4984
rect 15105 4981 15117 4984
rect 15151 4981 15163 5015
rect 15105 4975 15163 4981
rect 15657 5015 15715 5021
rect 15657 4981 15669 5015
rect 15703 5012 15715 5015
rect 15746 5012 15752 5024
rect 15703 4984 15752 5012
rect 15703 4981 15715 4984
rect 15657 4975 15715 4981
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 15838 4972 15844 5024
rect 15896 5012 15902 5024
rect 16040 5012 16068 5043
rect 15896 4984 16068 5012
rect 15896 4972 15902 4984
rect 16482 4972 16488 5024
rect 16540 4972 16546 5024
rect 16592 5012 16620 5111
rect 17126 5108 17132 5160
rect 17184 5108 17190 5160
rect 17313 5151 17371 5157
rect 17313 5117 17325 5151
rect 17359 5148 17371 5151
rect 17586 5148 17592 5160
rect 17359 5120 17592 5148
rect 17359 5117 17371 5120
rect 17313 5111 17371 5117
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 18064 5148 18092 5188
rect 18141 5185 18153 5219
rect 18187 5185 18199 5219
rect 18414 5216 18420 5228
rect 18141 5179 18199 5185
rect 18248 5188 18420 5216
rect 18248 5148 18276 5188
rect 18414 5176 18420 5188
rect 18472 5176 18478 5228
rect 20824 5225 20852 5256
rect 21818 5244 21824 5256
rect 21876 5244 21882 5296
rect 22002 5244 22008 5296
rect 22060 5284 22066 5296
rect 22094 5284 22100 5296
rect 22060 5256 22100 5284
rect 22060 5244 22066 5256
rect 22094 5244 22100 5256
rect 22152 5244 22158 5296
rect 22296 5284 22324 5324
rect 22646 5312 22652 5364
rect 22704 5352 22710 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 22704 5324 22753 5352
rect 22704 5312 22710 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 22741 5315 22799 5321
rect 22296 5256 23152 5284
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5216 18567 5219
rect 20809 5219 20867 5225
rect 18555 5188 18828 5216
rect 18555 5185 18567 5188
rect 18509 5179 18567 5185
rect 18064 5120 18276 5148
rect 18322 5108 18328 5160
rect 18380 5108 18386 5160
rect 18700 5151 18758 5157
rect 18700 5117 18712 5151
rect 18746 5117 18758 5151
rect 18800 5148 18828 5188
rect 20809 5185 20821 5219
rect 20855 5185 20867 5219
rect 21542 5216 21548 5228
rect 20809 5179 20867 5185
rect 21468 5188 21548 5216
rect 21468 5157 21496 5188
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 21910 5176 21916 5228
rect 21968 5176 21974 5228
rect 18949 5151 19007 5157
rect 18949 5148 18961 5151
rect 18800 5120 18961 5148
rect 18700 5111 18758 5117
rect 18949 5117 18961 5120
rect 18995 5117 19007 5151
rect 18949 5111 19007 5117
rect 20993 5151 21051 5157
rect 20993 5117 21005 5151
rect 21039 5148 21051 5151
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 21039 5120 21281 5148
rect 21039 5117 21051 5120
rect 20993 5111 21051 5117
rect 21269 5117 21281 5120
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 21453 5151 21511 5157
rect 21453 5117 21465 5151
rect 21499 5117 21511 5151
rect 21453 5111 21511 5117
rect 18506 5040 18512 5092
rect 18564 5080 18570 5092
rect 18708 5080 18736 5111
rect 21634 5108 21640 5160
rect 21692 5108 21698 5160
rect 22002 5108 22008 5160
rect 22060 5108 22066 5160
rect 22296 5157 22324 5256
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5216 22707 5219
rect 22738 5216 22744 5228
rect 22695 5188 22744 5216
rect 22695 5185 22707 5188
rect 22649 5179 22707 5185
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 22281 5151 22339 5157
rect 22281 5117 22293 5151
rect 22327 5117 22339 5151
rect 22281 5111 22339 5117
rect 22462 5108 22468 5160
rect 22520 5148 22526 5160
rect 23124 5157 23152 5256
rect 30558 5244 30564 5296
rect 30616 5284 30622 5296
rect 30653 5287 30711 5293
rect 30653 5284 30665 5287
rect 30616 5256 30665 5284
rect 30616 5244 30622 5256
rect 30653 5253 30665 5256
rect 30699 5253 30711 5287
rect 30653 5247 30711 5253
rect 23382 5176 23388 5228
rect 23440 5176 23446 5228
rect 25038 5176 25044 5228
rect 25096 5216 25102 5228
rect 26234 5225 26240 5228
rect 26053 5219 26111 5225
rect 26053 5216 26065 5219
rect 25096 5188 26065 5216
rect 25096 5176 25102 5188
rect 26053 5185 26065 5188
rect 26099 5185 26111 5219
rect 26053 5179 26111 5185
rect 26212 5219 26240 5225
rect 26212 5185 26224 5219
rect 26212 5179 26240 5185
rect 26234 5176 26240 5179
rect 26292 5176 26298 5228
rect 26326 5176 26332 5228
rect 26384 5176 26390 5228
rect 26602 5176 26608 5228
rect 26660 5176 26666 5228
rect 26878 5176 26884 5228
rect 26936 5216 26942 5228
rect 27065 5219 27123 5225
rect 27065 5216 27077 5219
rect 26936 5188 27077 5216
rect 26936 5176 26942 5188
rect 27065 5185 27077 5188
rect 27111 5185 27123 5219
rect 27065 5179 27123 5185
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5216 27307 5219
rect 27338 5216 27344 5228
rect 27295 5188 27344 5216
rect 27295 5185 27307 5188
rect 27249 5179 27307 5185
rect 27338 5176 27344 5188
rect 27396 5176 27402 5228
rect 29917 5219 29975 5225
rect 29917 5216 29929 5219
rect 29564 5188 29929 5216
rect 22925 5151 22983 5157
rect 22925 5148 22937 5151
rect 22520 5120 22937 5148
rect 22520 5108 22526 5120
rect 22925 5117 22937 5120
rect 22971 5117 22983 5151
rect 22925 5111 22983 5117
rect 23109 5151 23167 5157
rect 23109 5117 23121 5151
rect 23155 5117 23167 5151
rect 23109 5111 23167 5117
rect 23658 5108 23664 5160
rect 23716 5108 23722 5160
rect 27430 5108 27436 5160
rect 27488 5148 27494 5160
rect 28077 5151 28135 5157
rect 28077 5148 28089 5151
rect 27488 5120 28089 5148
rect 27488 5108 27494 5120
rect 28077 5117 28089 5120
rect 28123 5148 28135 5151
rect 28629 5151 28687 5157
rect 28629 5148 28641 5151
rect 28123 5120 28641 5148
rect 28123 5117 28135 5120
rect 28077 5111 28135 5117
rect 28629 5117 28641 5120
rect 28675 5117 28687 5151
rect 28629 5111 28687 5117
rect 29362 5108 29368 5160
rect 29420 5108 29426 5160
rect 29454 5108 29460 5160
rect 29512 5148 29518 5160
rect 29564 5157 29592 5188
rect 29917 5185 29929 5188
rect 29963 5185 29975 5219
rect 29917 5179 29975 5185
rect 30392 5188 30972 5216
rect 29549 5151 29607 5157
rect 29549 5148 29561 5151
rect 29512 5120 29561 5148
rect 29512 5108 29518 5120
rect 29549 5117 29561 5120
rect 29595 5117 29607 5151
rect 29549 5111 29607 5117
rect 29638 5108 29644 5160
rect 29696 5148 29702 5160
rect 30392 5148 30420 5188
rect 29696 5120 30420 5148
rect 29696 5108 29702 5120
rect 30466 5108 30472 5160
rect 30524 5148 30530 5160
rect 30561 5151 30619 5157
rect 30561 5148 30573 5151
rect 30524 5120 30573 5148
rect 30524 5108 30530 5120
rect 30561 5117 30573 5120
rect 30607 5117 30619 5151
rect 30561 5111 30619 5117
rect 18564 5052 18736 5080
rect 21545 5083 21603 5089
rect 18564 5040 18570 5052
rect 21545 5049 21557 5083
rect 21591 5080 21603 5083
rect 21591 5052 21680 5080
rect 21591 5049 21603 5052
rect 21545 5043 21603 5049
rect 21652 5024 21680 5052
rect 21726 5040 21732 5092
rect 21784 5089 21790 5092
rect 21784 5083 21813 5089
rect 21801 5080 21813 5083
rect 22143 5083 22201 5089
rect 22143 5080 22155 5083
rect 21801 5052 22155 5080
rect 21801 5049 21813 5052
rect 21784 5043 21813 5049
rect 22143 5049 22155 5052
rect 22189 5080 22201 5083
rect 22189 5052 22324 5080
rect 22189 5049 22201 5052
rect 22143 5043 22201 5049
rect 21784 5040 21790 5043
rect 19610 5012 19616 5024
rect 16592 4984 19616 5012
rect 19610 4972 19616 4984
rect 19668 4972 19674 5024
rect 21174 4972 21180 5024
rect 21232 4972 21238 5024
rect 21634 4972 21640 5024
rect 21692 4972 21698 5024
rect 22296 5012 22324 5052
rect 22370 5040 22376 5092
rect 22428 5040 22434 5092
rect 23014 5040 23020 5092
rect 23072 5040 23078 5092
rect 23227 5083 23285 5089
rect 23227 5049 23239 5083
rect 23273 5049 23285 5083
rect 23227 5043 23285 5049
rect 28169 5083 28227 5089
rect 28169 5049 28181 5083
rect 28215 5080 28227 5083
rect 28902 5080 28908 5092
rect 28215 5052 28908 5080
rect 28215 5049 28227 5052
rect 28169 5043 28227 5049
rect 23242 5012 23270 5043
rect 28902 5040 28908 5052
rect 28960 5040 28966 5092
rect 30576 5080 30604 5111
rect 30650 5108 30656 5160
rect 30708 5108 30714 5160
rect 30944 5157 30972 5188
rect 30929 5151 30987 5157
rect 30929 5117 30941 5151
rect 30975 5117 30987 5151
rect 30929 5111 30987 5117
rect 30837 5083 30895 5089
rect 30837 5080 30849 5083
rect 30576 5052 30849 5080
rect 30837 5049 30849 5052
rect 30883 5049 30895 5083
rect 30837 5043 30895 5049
rect 22296 4984 23270 5012
rect 23566 4972 23572 5024
rect 23624 4972 23630 5024
rect 25406 4972 25412 5024
rect 25464 4972 25470 5024
rect 28718 4972 28724 5024
rect 28776 4972 28782 5024
rect 28994 4972 29000 5024
rect 29052 5012 29058 5024
rect 29181 5015 29239 5021
rect 29181 5012 29193 5015
rect 29052 4984 29193 5012
rect 29052 4972 29058 4984
rect 29181 4981 29193 4984
rect 29227 4981 29239 5015
rect 29181 4975 29239 4981
rect 552 4922 31648 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 12096 4922
rect 12148 4870 12160 4922
rect 12212 4870 12224 4922
rect 12276 4870 12288 4922
rect 12340 4870 12352 4922
rect 12404 4870 19870 4922
rect 19922 4870 19934 4922
rect 19986 4870 19998 4922
rect 20050 4870 20062 4922
rect 20114 4870 20126 4922
rect 20178 4870 27644 4922
rect 27696 4870 27708 4922
rect 27760 4870 27772 4922
rect 27824 4870 27836 4922
rect 27888 4870 27900 4922
rect 27952 4870 31648 4922
rect 552 4848 31648 4870
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4777 3111 4811
rect 3053 4771 3111 4777
rect 3068 4740 3096 4771
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 3568 4780 4629 4808
rect 3568 4768 3574 4780
rect 4617 4777 4629 4780
rect 4663 4777 4675 4811
rect 4617 4771 4675 4777
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4808 5043 4811
rect 5166 4808 5172 4820
rect 5031 4780 5172 4808
rect 5031 4777 5043 4780
rect 4985 4771 5043 4777
rect 5166 4768 5172 4780
rect 5224 4808 5230 4820
rect 6638 4808 6644 4820
rect 5224 4780 6644 4808
rect 5224 4768 5230 4780
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 7374 4768 7380 4820
rect 7432 4768 7438 4820
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10468 4780 10609 4808
rect 10468 4768 10474 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 11057 4811 11115 4817
rect 11057 4777 11069 4811
rect 11103 4808 11115 4811
rect 11238 4808 11244 4820
rect 11103 4780 11244 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13722 4808 13728 4820
rect 13587 4780 13728 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14642 4768 14648 4820
rect 14700 4768 14706 4820
rect 18506 4768 18512 4820
rect 18564 4808 18570 4820
rect 18877 4811 18935 4817
rect 18877 4808 18889 4811
rect 18564 4780 18889 4808
rect 18564 4768 18570 4780
rect 18877 4777 18889 4780
rect 18923 4777 18935 4811
rect 21634 4808 21640 4820
rect 18877 4771 18935 4777
rect 20824 4780 21640 4808
rect 3326 4740 3332 4752
rect 3068 4712 3332 4740
rect 3326 4700 3332 4712
rect 3384 4740 3390 4752
rect 4890 4740 4896 4752
rect 3384 4712 4896 4740
rect 3384 4700 3390 4712
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 7653 4743 7711 4749
rect 7653 4740 7665 4743
rect 6972 4712 7665 4740
rect 6972 4700 6978 4712
rect 7653 4709 7665 4712
rect 7699 4709 7711 4743
rect 7653 4703 7711 4709
rect 7929 4743 7987 4749
rect 7929 4709 7941 4743
rect 7975 4740 7987 4743
rect 8202 4740 8208 4752
rect 7975 4712 8208 4740
rect 7975 4709 7987 4712
rect 7929 4703 7987 4709
rect 8202 4700 8208 4712
rect 8260 4740 8266 4752
rect 14660 4740 14688 4768
rect 16022 4740 16028 4752
rect 8260 4712 14688 4740
rect 15580 4712 16028 4740
rect 8260 4700 8266 4712
rect 1670 4632 1676 4684
rect 1728 4632 1734 4684
rect 1940 4675 1998 4681
rect 1940 4641 1952 4675
rect 1986 4672 1998 4675
rect 2498 4672 2504 4684
rect 1986 4644 2504 4672
rect 1986 4641 1998 4644
rect 1940 4635 1998 4641
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 3142 4632 3148 4684
rect 3200 4632 3206 4684
rect 3418 4681 3424 4684
rect 3412 4672 3424 4681
rect 3379 4644 3424 4672
rect 3412 4635 3424 4644
rect 3418 4632 3424 4635
rect 3476 4632 3482 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4540 4644 4813 4672
rect 4246 4496 4252 4548
rect 4304 4536 4310 4548
rect 4540 4545 4568 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 5132 4644 6193 4672
rect 5132 4632 5138 4644
rect 6181 4641 6193 4644
rect 6227 4672 6239 4675
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6227 4644 7113 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4641 7343 4675
rect 7285 4635 7343 4641
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 7834 4672 7840 4684
rect 7515 4644 7840 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 7300 4604 7328 4635
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 11054 4672 11060 4684
rect 10735 4644 11060 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11146 4632 11152 4684
rect 11204 4632 11210 4684
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 13354 4672 13360 4684
rect 13311 4644 13360 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 13449 4675 13507 4681
rect 13449 4641 13461 4675
rect 13495 4672 13507 4675
rect 14654 4675 14712 4681
rect 14654 4672 14666 4675
rect 13495 4644 14666 4672
rect 13495 4641 13507 4644
rect 13449 4635 13507 4641
rect 14654 4641 14666 4644
rect 14700 4641 14712 4675
rect 14654 4635 14712 4641
rect 14918 4632 14924 4684
rect 14976 4632 14982 4684
rect 15580 4681 15608 4712
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 16482 4740 16488 4752
rect 16132 4712 16488 4740
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 7650 4604 7656 4616
rect 7300 4576 7656 4604
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13127 4576 13215 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 4525 4539 4583 4545
rect 4525 4536 4537 4539
rect 4304 4508 4537 4536
rect 4304 4496 4310 4508
rect 4525 4505 4537 4508
rect 4571 4505 4583 4539
rect 4525 4499 4583 4505
rect 10042 4496 10048 4548
rect 10100 4536 10106 4548
rect 13187 4536 13215 4576
rect 10100 4508 13215 4536
rect 10100 4496 10106 4508
rect 6270 4428 6276 4480
rect 6328 4428 6334 4480
rect 13187 4468 13215 4508
rect 13538 4468 13544 4480
rect 13187 4440 13544 4468
rect 13538 4428 13544 4440
rect 13596 4468 13602 4480
rect 15580 4468 15608 4635
rect 15746 4632 15752 4684
rect 15804 4632 15810 4684
rect 16132 4681 16160 4712
rect 16482 4700 16488 4712
rect 16540 4700 16546 4752
rect 16666 4700 16672 4752
rect 16724 4740 16730 4752
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 16724 4712 18429 4740
rect 16724 4700 16730 4712
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 18417 4703 18475 4709
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16373 4675 16431 4681
rect 16373 4672 16385 4675
rect 16117 4635 16175 4641
rect 16224 4644 16385 4672
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16224 4604 16252 4644
rect 16373 4641 16385 4644
rect 16419 4641 16431 4675
rect 16373 4635 16431 4641
rect 17957 4675 18015 4681
rect 17957 4641 17969 4675
rect 18003 4672 18015 4675
rect 18230 4672 18236 4684
rect 18003 4644 18236 4672
rect 18003 4641 18015 4644
rect 17957 4635 18015 4641
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 15979 4576 16252 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 17586 4564 17592 4616
rect 17644 4564 17650 4616
rect 18046 4564 18052 4616
rect 18104 4564 18110 4616
rect 18432 4604 18460 4703
rect 18598 4700 18604 4752
rect 18656 4740 18662 4752
rect 20533 4743 20591 4749
rect 20533 4740 20545 4743
rect 18656 4712 20545 4740
rect 18656 4700 18662 4712
rect 20533 4709 20545 4712
rect 20579 4740 20591 4743
rect 20622 4740 20628 4752
rect 20579 4712 20628 4740
rect 20579 4709 20591 4712
rect 20533 4703 20591 4709
rect 20622 4700 20628 4712
rect 20680 4700 20686 4752
rect 18969 4675 19027 4681
rect 18969 4641 18981 4675
rect 19015 4672 19027 4675
rect 19610 4672 19616 4684
rect 19015 4644 19616 4672
rect 19015 4641 19027 4644
rect 18969 4635 19027 4641
rect 19610 4632 19616 4644
rect 19668 4632 19674 4684
rect 20714 4632 20720 4684
rect 20772 4632 20778 4684
rect 20824 4681 20852 4780
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 25406 4768 25412 4820
rect 25464 4808 25470 4820
rect 25685 4811 25743 4817
rect 25685 4808 25697 4811
rect 25464 4780 25697 4808
rect 25464 4768 25470 4780
rect 25685 4777 25697 4780
rect 25731 4777 25743 4811
rect 25685 4771 25743 4777
rect 27893 4811 27951 4817
rect 27893 4777 27905 4811
rect 27939 4808 27951 4811
rect 28074 4808 28080 4820
rect 27939 4780 28080 4808
rect 27939 4777 27951 4780
rect 27893 4771 27951 4777
rect 28074 4768 28080 4780
rect 28132 4768 28138 4820
rect 28994 4768 29000 4820
rect 29052 4768 29058 4820
rect 29181 4811 29239 4817
rect 29181 4777 29193 4811
rect 29227 4777 29239 4811
rect 29181 4771 29239 4777
rect 21174 4700 21180 4752
rect 21232 4740 21238 4752
rect 21514 4743 21572 4749
rect 21514 4740 21526 4743
rect 21232 4712 21526 4740
rect 21232 4700 21238 4712
rect 21514 4709 21526 4712
rect 21560 4709 21572 4743
rect 23566 4740 23572 4752
rect 21514 4703 21572 4709
rect 23032 4712 23572 4740
rect 20809 4675 20867 4681
rect 20809 4641 20821 4675
rect 20855 4641 20867 4675
rect 20809 4635 20867 4641
rect 21082 4632 21088 4684
rect 21140 4632 21146 4684
rect 21266 4632 21272 4684
rect 21324 4632 21330 4684
rect 23032 4681 23060 4712
rect 23566 4700 23572 4712
rect 23624 4700 23630 4752
rect 27985 4743 28043 4749
rect 27985 4709 27997 4743
rect 28031 4740 28043 4743
rect 28166 4740 28172 4752
rect 28031 4712 28172 4740
rect 28031 4709 28043 4712
rect 27985 4703 28043 4709
rect 28166 4700 28172 4712
rect 28224 4700 28230 4752
rect 29196 4740 29224 4771
rect 29362 4768 29368 4820
rect 29420 4808 29426 4820
rect 30653 4811 30711 4817
rect 30653 4808 30665 4811
rect 29420 4780 30665 4808
rect 29420 4768 29426 4780
rect 30653 4777 30665 4780
rect 30699 4777 30711 4811
rect 30653 4771 30711 4777
rect 29518 4743 29576 4749
rect 29518 4740 29530 4743
rect 29196 4712 29530 4740
rect 29518 4709 29530 4712
rect 29564 4709 29576 4743
rect 29518 4703 29576 4709
rect 23017 4675 23075 4681
rect 23017 4641 23029 4675
rect 23063 4641 23075 4675
rect 23017 4635 23075 4641
rect 23106 4632 23112 4684
rect 23164 4672 23170 4684
rect 23273 4675 23331 4681
rect 23273 4672 23285 4675
rect 23164 4644 23285 4672
rect 23164 4632 23170 4644
rect 23273 4641 23285 4644
rect 23319 4641 23331 4675
rect 23273 4635 23331 4641
rect 28074 4632 28080 4684
rect 28132 4632 28138 4684
rect 28353 4675 28411 4681
rect 28353 4641 28365 4675
rect 28399 4641 28411 4675
rect 28353 4635 28411 4641
rect 28537 4675 28595 4681
rect 28537 4641 28549 4675
rect 28583 4641 28595 4675
rect 28537 4635 28595 4641
rect 20070 4604 20076 4616
rect 18432 4576 20076 4604
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 25774 4564 25780 4616
rect 25832 4564 25838 4616
rect 25869 4607 25927 4613
rect 25869 4573 25881 4607
rect 25915 4573 25927 4607
rect 25869 4567 25927 4573
rect 27709 4607 27767 4613
rect 27709 4573 27721 4607
rect 27755 4604 27767 4607
rect 27982 4604 27988 4616
rect 27755 4576 27988 4604
rect 27755 4573 27767 4576
rect 27709 4567 27767 4573
rect 25682 4536 25688 4548
rect 24412 4508 25688 4536
rect 13596 4440 15608 4468
rect 13596 4428 13602 4440
rect 15930 4428 15936 4480
rect 15988 4468 15994 4480
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 15988 4440 17509 4468
rect 15988 4428 15994 4440
rect 17497 4437 17509 4440
rect 17543 4437 17555 4471
rect 17497 4431 17555 4437
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 18012 4440 18245 4468
rect 18012 4428 18018 4440
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 20993 4471 21051 4477
rect 20993 4437 21005 4471
rect 21039 4468 21051 4471
rect 21542 4468 21548 4480
rect 21039 4440 21548 4468
rect 21039 4437 21051 4440
rect 20993 4431 21051 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 22646 4428 22652 4480
rect 22704 4428 22710 4480
rect 23014 4428 23020 4480
rect 23072 4468 23078 4480
rect 24412 4477 24440 4508
rect 25682 4496 25688 4508
rect 25740 4536 25746 4548
rect 25884 4536 25912 4567
rect 27982 4564 27988 4576
rect 28040 4604 28046 4616
rect 28368 4604 28396 4635
rect 28040 4576 28396 4604
rect 28552 4604 28580 4635
rect 28718 4632 28724 4684
rect 28776 4672 28782 4684
rect 29273 4675 29331 4681
rect 29273 4672 29285 4675
rect 28776 4644 29285 4672
rect 28776 4632 28782 4644
rect 29273 4641 29285 4644
rect 29319 4641 29331 4675
rect 29273 4635 29331 4641
rect 28994 4604 29000 4616
rect 28552 4576 29000 4604
rect 28040 4564 28046 4576
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 25740 4508 25912 4536
rect 25740 4496 25746 4508
rect 28258 4496 28264 4548
rect 28316 4496 28322 4548
rect 28629 4539 28687 4545
rect 28629 4505 28641 4539
rect 28675 4536 28687 4539
rect 29086 4536 29092 4548
rect 28675 4508 29092 4536
rect 28675 4505 28687 4508
rect 28629 4499 28687 4505
rect 29086 4496 29092 4508
rect 29144 4496 29150 4548
rect 24397 4471 24455 4477
rect 24397 4468 24409 4471
rect 23072 4440 24409 4468
rect 23072 4428 23078 4440
rect 24397 4437 24409 4440
rect 24443 4437 24455 4471
rect 24397 4431 24455 4437
rect 25314 4428 25320 4480
rect 25372 4428 25378 4480
rect 28534 4428 28540 4480
rect 28592 4428 28598 4480
rect 28997 4471 29055 4477
rect 28997 4437 29009 4471
rect 29043 4468 29055 4471
rect 29178 4468 29184 4480
rect 29043 4440 29184 4468
rect 29043 4437 29055 4440
rect 28997 4431 29055 4437
rect 29178 4428 29184 4440
rect 29236 4428 29242 4480
rect 552 4378 31648 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 11436 4378
rect 11488 4326 11500 4378
rect 11552 4326 11564 4378
rect 11616 4326 11628 4378
rect 11680 4326 11692 4378
rect 11744 4326 19210 4378
rect 19262 4326 19274 4378
rect 19326 4326 19338 4378
rect 19390 4326 19402 4378
rect 19454 4326 19466 4378
rect 19518 4326 26984 4378
rect 27036 4326 27048 4378
rect 27100 4326 27112 4378
rect 27164 4326 27176 4378
rect 27228 4326 27240 4378
rect 27292 4326 31648 4378
rect 552 4304 31648 4326
rect 2498 4224 2504 4276
rect 2556 4264 2562 4276
rect 2685 4267 2743 4273
rect 2685 4264 2697 4267
rect 2556 4236 2697 4264
rect 2556 4224 2562 4236
rect 2685 4233 2697 4236
rect 2731 4233 2743 4267
rect 2685 4227 2743 4233
rect 2869 4267 2927 4273
rect 2869 4233 2881 4267
rect 2915 4264 2927 4267
rect 4062 4264 4068 4276
rect 2915 4236 4068 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 4764 4236 5089 4264
rect 4764 4224 4770 4236
rect 5077 4233 5089 4236
rect 5123 4264 5135 4267
rect 5166 4264 5172 4276
rect 5123 4236 5172 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 6733 4267 6791 4273
rect 6733 4233 6745 4267
rect 6779 4264 6791 4267
rect 6822 4264 6828 4276
rect 6779 4236 6828 4264
rect 6779 4233 6791 4236
rect 6733 4227 6791 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7834 4224 7840 4276
rect 7892 4264 7898 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 7892 4236 8217 4264
rect 7892 4224 7898 4236
rect 8205 4233 8217 4236
rect 8251 4233 8263 4267
rect 8205 4227 8263 4233
rect 8573 4267 8631 4273
rect 8573 4233 8585 4267
rect 8619 4264 8631 4267
rect 8754 4264 8760 4276
rect 8619 4236 8760 4264
rect 8619 4233 8631 4236
rect 8573 4227 8631 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13136 4236 14688 4264
rect 13136 4224 13142 4236
rect 14660 4196 14688 4236
rect 14734 4224 14740 4276
rect 14792 4264 14798 4276
rect 14921 4267 14979 4273
rect 14921 4264 14933 4267
rect 14792 4236 14933 4264
rect 14792 4224 14798 4236
rect 14921 4233 14933 4236
rect 14967 4233 14979 4267
rect 14921 4227 14979 4233
rect 16853 4267 16911 4273
rect 16853 4233 16865 4267
rect 16899 4264 16911 4267
rect 17126 4264 17132 4276
rect 16899 4236 17132 4264
rect 16899 4233 16911 4236
rect 16853 4227 16911 4233
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17770 4224 17776 4276
rect 17828 4224 17834 4276
rect 18322 4224 18328 4276
rect 18380 4264 18386 4276
rect 19610 4264 19616 4276
rect 18380 4236 19616 4264
rect 18380 4224 18386 4236
rect 19610 4224 19616 4236
rect 19668 4224 19674 4276
rect 20070 4224 20076 4276
rect 20128 4224 20134 4276
rect 21542 4224 21548 4276
rect 21600 4264 21606 4276
rect 22005 4267 22063 4273
rect 22005 4264 22017 4267
rect 21600 4236 22017 4264
rect 21600 4224 21606 4236
rect 22005 4233 22017 4236
rect 22051 4233 22063 4267
rect 25314 4264 25320 4276
rect 22005 4227 22063 4233
rect 22112 4236 25320 4264
rect 15838 4196 15844 4208
rect 14660 4168 15844 4196
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 17405 4199 17463 4205
rect 17405 4165 17417 4199
rect 17451 4165 17463 4199
rect 17405 4159 17463 4165
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16393 4131 16451 4137
rect 16393 4128 16405 4131
rect 15988 4100 16405 4128
rect 15988 4088 15994 4100
rect 16393 4097 16405 4100
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 17310 4088 17316 4140
rect 17368 4128 17374 4140
rect 17420 4128 17448 4159
rect 20714 4156 20720 4208
rect 20772 4196 20778 4208
rect 22112 4196 22140 4236
rect 25314 4224 25320 4236
rect 25372 4224 25378 4276
rect 25774 4224 25780 4276
rect 25832 4264 25838 4276
rect 26145 4267 26203 4273
rect 26145 4264 26157 4267
rect 25832 4236 26157 4264
rect 25832 4224 25838 4236
rect 26145 4233 26157 4236
rect 26191 4233 26203 4267
rect 26145 4227 26203 4233
rect 26602 4224 26608 4276
rect 26660 4264 26666 4276
rect 28997 4267 29055 4273
rect 26660 4236 27384 4264
rect 26660 4224 26666 4236
rect 20772 4168 22140 4196
rect 20772 4156 20778 4168
rect 17368 4100 18828 4128
rect 17368 4088 17374 4100
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 3384 4032 3433 4060
rect 3384 4020 3390 4032
rect 3421 4029 3433 4032
rect 3467 4029 3479 4063
rect 3421 4023 3479 4029
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 3568 4032 3617 4060
rect 3568 4020 3574 4032
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 3786 4060 3792 4072
rect 3743 4032 3792 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 5350 4020 5356 4072
rect 5408 4020 5414 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 8941 4063 8999 4069
rect 8941 4060 8953 4063
rect 8720 4032 8953 4060
rect 8720 4020 8726 4032
rect 8941 4029 8953 4032
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11238 4060 11244 4072
rect 11112 4032 11244 4060
rect 11112 4020 11118 4032
rect 11238 4020 11244 4032
rect 11296 4060 11302 4072
rect 13814 4069 13820 4072
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 11296 4032 13185 4060
rect 11296 4020 11302 4032
rect 13173 4029 13185 4032
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13311 4032 13553 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13808 4060 13820 4069
rect 13775 4032 13820 4060
rect 13541 4023 13599 4029
rect 13808 4023 13820 4032
rect 13814 4020 13820 4023
rect 13872 4020 13878 4072
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 16485 4063 16543 4069
rect 16485 4060 16497 4063
rect 14424 4032 16497 4060
rect 14424 4020 14430 4032
rect 16485 4029 16497 4032
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 18322 4060 18328 4072
rect 16632 4032 18328 4060
rect 16632 4020 16638 4032
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 18693 4063 18751 4069
rect 18693 4060 18705 4063
rect 18463 4032 18705 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18693 4029 18705 4032
rect 18739 4029 18751 4063
rect 18800 4060 18828 4100
rect 18800 4032 19334 4060
rect 18693 4023 18751 4029
rect 3970 4001 3976 4004
rect 3053 3995 3111 4001
rect 3053 3961 3065 3995
rect 3099 3992 3111 3995
rect 3237 3995 3295 4001
rect 3237 3992 3249 3995
rect 3099 3964 3249 3992
rect 3099 3961 3111 3964
rect 3053 3955 3111 3961
rect 3237 3961 3249 3964
rect 3283 3961 3295 3995
rect 3237 3955 3295 3961
rect 3964 3955 3976 4001
rect 3970 3952 3976 3955
rect 4028 3952 4034 4004
rect 5620 3995 5678 4001
rect 5620 3961 5632 3995
rect 5666 3992 5678 3995
rect 5810 3992 5816 4004
rect 5666 3964 5816 3992
rect 5666 3961 5678 3964
rect 5620 3955 5678 3961
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 7092 3995 7150 4001
rect 7092 3961 7104 3995
rect 7138 3992 7150 3995
rect 7138 3964 8432 3992
rect 7138 3961 7150 3964
rect 7092 3955 7150 3961
rect 2853 3927 2911 3933
rect 2853 3893 2865 3927
rect 2899 3924 2911 3927
rect 3326 3924 3332 3936
rect 2899 3896 3332 3924
rect 2899 3893 2911 3896
rect 2853 3887 2911 3893
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 8404 3933 8432 3964
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 13998 3992 14004 4004
rect 10100 3964 14004 3992
rect 10100 3952 10106 3964
rect 13998 3952 14004 3964
rect 14056 3952 14062 4004
rect 18938 3995 18996 4001
rect 18938 3992 18950 3995
rect 18432 3964 18950 3992
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 8570 3884 8576 3936
rect 8628 3884 8634 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 11020 3896 11161 3924
rect 11020 3884 11026 3896
rect 11149 3893 11161 3896
rect 11195 3893 11207 3927
rect 11149 3887 11207 3893
rect 17773 3927 17831 3933
rect 17773 3893 17785 3927
rect 17819 3924 17831 3927
rect 17862 3924 17868 3936
rect 17819 3896 17868 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 17957 3927 18015 3933
rect 17957 3893 17969 3927
rect 18003 3924 18015 3927
rect 18432 3924 18460 3964
rect 18938 3961 18950 3964
rect 18984 3961 18996 3995
rect 18938 3955 18996 3961
rect 18003 3896 18460 3924
rect 19306 3924 19334 4032
rect 20070 4020 20076 4072
rect 20128 4060 20134 4072
rect 21376 4069 21404 4168
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 27356 4205 27384 4236
rect 28997 4233 29009 4267
rect 29043 4264 29055 4267
rect 29086 4264 29092 4276
rect 29043 4236 29092 4264
rect 29043 4233 29055 4236
rect 28997 4227 29055 4233
rect 29086 4224 29092 4236
rect 29144 4224 29150 4276
rect 29181 4267 29239 4273
rect 29181 4233 29193 4267
rect 29227 4264 29239 4267
rect 29362 4264 29368 4276
rect 29227 4236 29368 4264
rect 29227 4233 29239 4236
rect 29181 4227 29239 4233
rect 25409 4199 25467 4205
rect 25409 4196 25421 4199
rect 24912 4168 25421 4196
rect 24912 4156 24918 4168
rect 25409 4165 25421 4168
rect 25455 4165 25467 4199
rect 25409 4159 25467 4165
rect 27341 4199 27399 4205
rect 27341 4165 27353 4199
rect 27387 4165 27399 4199
rect 28074 4196 28080 4208
rect 27341 4159 27399 4165
rect 28000 4168 28080 4196
rect 21453 4131 21511 4137
rect 21453 4097 21465 4131
rect 21499 4128 21511 4131
rect 21634 4128 21640 4140
rect 21499 4100 21640 4128
rect 21499 4097 21511 4100
rect 21453 4091 21511 4097
rect 21634 4088 21640 4100
rect 21692 4128 21698 4140
rect 22646 4128 22652 4140
rect 21692 4100 22652 4128
rect 21692 4088 21698 4100
rect 22646 4088 22652 4100
rect 22704 4088 22710 4140
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 25740 4100 25789 4128
rect 25740 4088 25746 4100
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 26789 4131 26847 4137
rect 26789 4128 26801 4131
rect 25777 4091 25835 4097
rect 25884 4100 26801 4128
rect 21177 4063 21235 4069
rect 21177 4060 21189 4063
rect 20128 4032 21189 4060
rect 20128 4020 20134 4032
rect 21177 4029 21189 4032
rect 21223 4029 21235 4063
rect 21177 4023 21235 4029
rect 21360 4063 21418 4069
rect 21360 4029 21372 4063
rect 21406 4029 21418 4063
rect 21360 4023 21418 4029
rect 21542 4020 21548 4072
rect 21600 4020 21606 4072
rect 21729 4063 21787 4069
rect 21729 4029 21741 4063
rect 21775 4029 21787 4063
rect 21729 4023 21787 4029
rect 21082 3952 21088 4004
rect 21140 3992 21146 4004
rect 21744 3992 21772 4023
rect 22186 4020 22192 4072
rect 22244 4020 22250 4072
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4060 22339 4063
rect 23014 4060 23020 4072
rect 22327 4032 23020 4060
rect 22327 4029 22339 4032
rect 22281 4023 22339 4029
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4029 23535 4063
rect 23477 4023 23535 4029
rect 23569 4063 23627 4069
rect 23569 4029 23581 4063
rect 23615 4060 23627 4063
rect 23845 4063 23903 4069
rect 23845 4060 23857 4063
rect 23615 4032 23857 4060
rect 23615 4029 23627 4032
rect 23569 4023 23627 4029
rect 23845 4029 23857 4032
rect 23891 4029 23903 4063
rect 23845 4023 23903 4029
rect 23492 3992 23520 4023
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 24101 4063 24159 4069
rect 24101 4060 24113 4063
rect 23992 4032 24113 4060
rect 23992 4020 23998 4032
rect 24101 4029 24113 4032
rect 24147 4029 24159 4063
rect 24101 4023 24159 4029
rect 25038 4020 25044 4072
rect 25096 4060 25102 4072
rect 25884 4060 25912 4100
rect 26789 4097 26801 4100
rect 26835 4097 26847 4131
rect 26789 4091 26847 4097
rect 27065 4131 27123 4137
rect 27065 4097 27077 4131
rect 27111 4128 27123 4131
rect 27246 4128 27252 4140
rect 27111 4100 27252 4128
rect 27111 4097 27123 4100
rect 27065 4091 27123 4097
rect 27246 4088 27252 4100
rect 27304 4088 27310 4140
rect 28000 4137 28028 4168
rect 28074 4156 28080 4168
rect 28132 4196 28138 4208
rect 29196 4196 29224 4227
rect 29362 4224 29368 4236
rect 29420 4224 29426 4276
rect 29454 4224 29460 4276
rect 29512 4224 29518 4276
rect 28132 4168 29224 4196
rect 28132 4156 28138 4168
rect 27985 4131 28043 4137
rect 27985 4097 27997 4131
rect 28031 4097 28043 4131
rect 27985 4091 28043 4097
rect 28166 4088 28172 4140
rect 28224 4088 28230 4140
rect 28258 4088 28264 4140
rect 28316 4128 28322 4140
rect 29472 4128 29500 4224
rect 28316 4100 29500 4128
rect 28316 4088 28322 4100
rect 26970 4069 26976 4072
rect 25096 4032 25912 4060
rect 26948 4063 26976 4069
rect 25096 4020 25102 4032
rect 26948 4029 26960 4063
rect 26948 4023 26976 4029
rect 26970 4020 26976 4023
rect 27028 4020 27034 4072
rect 27801 4063 27859 4069
rect 27801 4029 27813 4063
rect 27847 4060 27859 4063
rect 28276 4060 28304 4088
rect 27847 4032 28304 4060
rect 27847 4029 27859 4032
rect 27801 4023 27859 4029
rect 23658 3992 23664 4004
rect 21140 3964 23428 3992
rect 23492 3964 23664 3992
rect 21140 3952 21146 3964
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 19306 3896 21833 3924
rect 18003 3893 18015 3896
rect 17957 3887 18015 3893
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 23400 3924 23428 3964
rect 23658 3952 23664 3964
rect 23716 3952 23722 4004
rect 29365 3995 29423 4001
rect 24228 3964 25360 3992
rect 24228 3924 24256 3964
rect 23400 3896 24256 3924
rect 21821 3887 21879 3893
rect 25038 3884 25044 3936
rect 25096 3924 25102 3936
rect 25332 3933 25360 3964
rect 29365 3961 29377 3995
rect 29411 3992 29423 3995
rect 29472 3992 29500 4100
rect 30837 4131 30895 4137
rect 30837 4097 30849 4131
rect 30883 4128 30895 4131
rect 31021 4131 31079 4137
rect 31021 4128 31033 4131
rect 30883 4100 31033 4128
rect 30883 4097 30895 4100
rect 30837 4091 30895 4097
rect 31021 4097 31033 4100
rect 31067 4097 31079 4131
rect 31021 4091 31079 4097
rect 30558 4020 30564 4072
rect 30616 4069 30622 4072
rect 30616 4060 30628 4069
rect 30616 4032 30661 4060
rect 30616 4023 30628 4032
rect 30616 4020 30622 4023
rect 30926 4020 30932 4072
rect 30984 4020 30990 4072
rect 29411 3964 29500 3992
rect 29411 3961 29423 3964
rect 29365 3955 29423 3961
rect 25225 3927 25283 3933
rect 25225 3924 25237 3927
rect 25096 3896 25237 3924
rect 25096 3884 25102 3896
rect 25225 3893 25237 3896
rect 25271 3893 25283 3927
rect 25225 3887 25283 3893
rect 25317 3927 25375 3933
rect 25317 3893 25329 3927
rect 25363 3893 25375 3927
rect 25317 3887 25375 3893
rect 28810 3884 28816 3936
rect 28868 3884 28874 3936
rect 29165 3927 29223 3933
rect 29165 3893 29177 3927
rect 29211 3924 29223 3927
rect 29638 3924 29644 3936
rect 29211 3896 29644 3924
rect 29211 3893 29223 3896
rect 29165 3887 29223 3893
rect 29638 3884 29644 3896
rect 29696 3884 29702 3936
rect 552 3834 31648 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 12096 3834
rect 12148 3782 12160 3834
rect 12212 3782 12224 3834
rect 12276 3782 12288 3834
rect 12340 3782 12352 3834
rect 12404 3782 19870 3834
rect 19922 3782 19934 3834
rect 19986 3782 19998 3834
rect 20050 3782 20062 3834
rect 20114 3782 20126 3834
rect 20178 3782 27644 3834
rect 27696 3782 27708 3834
rect 27760 3782 27772 3834
rect 27824 3782 27836 3834
rect 27888 3782 27900 3834
rect 27952 3782 31648 3834
rect 552 3760 31648 3782
rect 3326 3680 3332 3732
rect 3384 3680 3390 3732
rect 3786 3680 3792 3732
rect 3844 3680 3850 3732
rect 3970 3680 3976 3732
rect 4028 3680 4034 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4614 3720 4620 3732
rect 4120 3692 4620 3720
rect 4120 3680 4126 3692
rect 4614 3680 4620 3692
rect 4672 3720 4678 3732
rect 4672 3692 5304 3720
rect 4672 3680 4678 3692
rect 4154 3652 4160 3664
rect 3896 3624 4160 3652
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 3292 3556 3341 3584
rect 3292 3544 3298 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3329 3547 3387 3553
rect 3510 3544 3516 3596
rect 3568 3544 3574 3596
rect 3896 3593 3924 3624
rect 4154 3612 4160 3624
rect 4212 3652 4218 3664
rect 5276 3652 5304 3692
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5408 3692 5549 3720
rect 5408 3680 5414 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 5537 3683 5595 3689
rect 5810 3680 5816 3732
rect 5868 3680 5874 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 8205 3723 8263 3729
rect 7432 3692 7604 3720
rect 7432 3680 7438 3692
rect 4212 3624 5212 3652
rect 5276 3624 6500 3652
rect 4212 3612 4218 3624
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3553 3939 3587
rect 3881 3547 3939 3553
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3553 4399 3587
rect 4341 3547 4399 3553
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 4264 3380 4292 3547
rect 4356 3448 4384 3547
rect 4448 3516 4476 3547
rect 4614 3544 4620 3596
rect 4672 3544 4678 3596
rect 4706 3544 4712 3596
rect 4764 3544 4770 3596
rect 4893 3587 4951 3593
rect 4893 3553 4905 3587
rect 4939 3584 4951 3587
rect 5074 3584 5080 3596
rect 4939 3556 5080 3584
rect 4939 3553 4951 3556
rect 4893 3547 4951 3553
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4448 3488 4813 3516
rect 4801 3485 4813 3488
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4908 3448 4936 3547
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5184 3584 5212 3624
rect 5626 3584 5632 3596
rect 5184 3556 5632 3584
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 6089 3587 6147 3593
rect 6089 3553 6101 3587
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 6104 3516 6132 3547
rect 6178 3544 6184 3596
rect 6236 3544 6242 3596
rect 6270 3544 6276 3596
rect 6328 3544 6334 3596
rect 6472 3593 6500 3624
rect 7576 3596 7604 3692
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 8570 3720 8576 3732
rect 8251 3692 8576 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 11054 3720 11060 3732
rect 10520 3692 11060 3720
rect 8389 3655 8447 3661
rect 8389 3652 8401 3655
rect 7760 3624 8401 3652
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6503 3556 6684 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6104 3488 6561 3516
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 4356 3420 4936 3448
rect 6656 3448 6684 3556
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6972 3556 7113 3584
rect 6972 3544 6978 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 7558 3544 7564 3596
rect 7616 3544 7622 3596
rect 7650 3544 7656 3596
rect 7708 3544 7714 3596
rect 7760 3593 7788 3624
rect 8036 3593 8064 3624
rect 8389 3621 8401 3624
rect 8435 3652 8447 3655
rect 8435 3624 8616 3652
rect 8435 3621 8447 3624
rect 8389 3615 8447 3621
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3553 7987 3587
rect 7929 3547 7987 3553
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3553 8079 3587
rect 8021 3547 8079 3553
rect 7944 3516 7972 3547
rect 8202 3544 8208 3596
rect 8260 3544 8266 3596
rect 8294 3544 8300 3596
rect 8352 3544 8358 3596
rect 8478 3544 8484 3596
rect 8536 3544 8542 3596
rect 8588 3593 8616 3624
rect 8662 3612 8668 3664
rect 8720 3612 8726 3664
rect 9953 3655 10011 3661
rect 9953 3621 9965 3655
rect 9999 3652 10011 3655
rect 9999 3624 10364 3652
rect 9999 3621 10011 3624
rect 9953 3615 10011 3621
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3553 8631 3587
rect 8573 3547 8631 3553
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3553 8815 3587
rect 9766 3584 9772 3596
rect 8757 3547 8815 3553
rect 8864 3556 9772 3584
rect 8662 3516 8668 3528
rect 7944 3488 8668 3516
rect 7944 3448 7972 3488
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 6656 3420 7972 3448
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 8772 3448 8800 3547
rect 8260 3420 8800 3448
rect 8260 3408 8266 3420
rect 4706 3380 4712 3392
rect 4264 3352 4712 3380
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 7285 3383 7343 3389
rect 7285 3380 7297 3383
rect 7156 3352 7297 3380
rect 7156 3340 7162 3352
rect 7285 3349 7297 3352
rect 7331 3349 7343 3383
rect 7285 3343 7343 3349
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 8478 3380 8484 3392
rect 7708 3352 8484 3380
rect 7708 3340 7714 3352
rect 8478 3340 8484 3352
rect 8536 3380 8542 3392
rect 8864 3380 8892 3556
rect 9766 3544 9772 3556
rect 9824 3584 9830 3596
rect 10336 3593 10364 3624
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9824 3556 9873 3584
rect 9824 3544 9830 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9398 3516 9404 3528
rect 8996 3488 9404 3516
rect 8996 3476 9002 3488
rect 9398 3476 9404 3488
rect 9456 3516 9462 3528
rect 10152 3516 10180 3547
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 10520 3593 10548 3692
rect 11054 3680 11060 3692
rect 11112 3720 11118 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 11112 3692 12357 3720
rect 11112 3680 11118 3692
rect 12345 3689 12357 3692
rect 12391 3720 12403 3723
rect 14366 3720 14372 3732
rect 12391 3692 14372 3720
rect 12391 3689 12403 3692
rect 12345 3683 12403 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 26970 3680 26976 3732
rect 27028 3720 27034 3732
rect 27525 3723 27583 3729
rect 27525 3720 27537 3723
rect 27028 3692 27537 3720
rect 27028 3680 27034 3692
rect 27525 3689 27537 3692
rect 27571 3720 27583 3723
rect 28166 3720 28172 3732
rect 27571 3692 28172 3720
rect 27571 3689 27583 3692
rect 27525 3683 27583 3689
rect 28166 3680 28172 3692
rect 28224 3680 28230 3732
rect 28994 3680 29000 3732
rect 29052 3680 29058 3732
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 11210 3655 11268 3661
rect 11210 3652 11222 3655
rect 10827 3624 11222 3652
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 11210 3621 11222 3624
rect 11256 3621 11268 3655
rect 11210 3615 11268 3621
rect 20990 3612 20996 3664
rect 21048 3612 21054 3664
rect 28534 3612 28540 3664
rect 28592 3652 28598 3664
rect 28638 3655 28696 3661
rect 28638 3652 28650 3655
rect 28592 3624 28650 3652
rect 28592 3612 28598 3624
rect 28638 3621 28650 3624
rect 28684 3621 28696 3655
rect 28638 3615 28696 3621
rect 28810 3612 28816 3664
rect 28868 3652 28874 3664
rect 28868 3624 29316 3652
rect 28868 3612 28874 3624
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 10962 3544 10968 3596
rect 11020 3544 11026 3596
rect 11072 3556 14872 3584
rect 9456 3488 10180 3516
rect 9456 3476 9462 3488
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 11072 3516 11100 3556
rect 10284 3488 11100 3516
rect 10284 3476 10290 3488
rect 14844 3460 14872 3556
rect 16482 3544 16488 3596
rect 16540 3544 16546 3596
rect 19794 3544 19800 3596
rect 19852 3584 19858 3596
rect 19981 3587 20039 3593
rect 19981 3584 19993 3587
rect 19852 3556 19993 3584
rect 19852 3544 19858 3556
rect 19981 3553 19993 3556
rect 20027 3553 20039 3587
rect 19981 3547 20039 3553
rect 20346 3544 20352 3596
rect 20404 3584 20410 3596
rect 20441 3587 20499 3593
rect 20441 3584 20453 3587
rect 20404 3556 20453 3584
rect 20404 3544 20410 3556
rect 20441 3553 20453 3556
rect 20487 3584 20499 3587
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20487 3556 20821 3584
rect 20487 3553 20499 3556
rect 20441 3547 20499 3553
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 28902 3544 28908 3596
rect 28960 3544 28966 3596
rect 29086 3544 29092 3596
rect 29144 3584 29150 3596
rect 29288 3593 29316 3624
rect 29181 3587 29239 3593
rect 29181 3584 29193 3587
rect 29144 3556 29193 3584
rect 29144 3544 29150 3556
rect 29181 3553 29193 3556
rect 29227 3553 29239 3587
rect 29181 3547 29239 3553
rect 29273 3587 29331 3593
rect 29273 3553 29285 3587
rect 29319 3553 29331 3587
rect 29273 3547 29331 3553
rect 20717 3519 20775 3525
rect 20717 3485 20729 3519
rect 20763 3516 20775 3519
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20763 3488 21281 3516
rect 20763 3485 20775 3488
rect 20717 3479 20775 3485
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 21910 3476 21916 3528
rect 21968 3476 21974 3528
rect 28997 3519 29055 3525
rect 28997 3485 29009 3519
rect 29043 3485 29055 3519
rect 28997 3479 29055 3485
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 10008 3420 10732 3448
rect 10008 3408 10014 3420
rect 8536 3352 8892 3380
rect 10704 3380 10732 3420
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 16850 3448 16856 3460
rect 14884 3420 16856 3448
rect 14884 3408 14890 3420
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 15194 3380 15200 3392
rect 10704 3352 15200 3380
rect 8536 3340 8542 3352
rect 15194 3340 15200 3352
rect 15252 3340 15258 3392
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 16264 3352 16405 3380
rect 16264 3340 16270 3352
rect 16393 3349 16405 3352
rect 16439 3349 16451 3383
rect 16393 3343 16451 3349
rect 19702 3340 19708 3392
rect 19760 3380 19766 3392
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 19760 3352 19901 3380
rect 19760 3340 19766 3352
rect 19889 3349 19901 3352
rect 19935 3349 19947 3383
rect 19889 3343 19947 3349
rect 20254 3340 20260 3392
rect 20312 3340 20318 3392
rect 20622 3340 20628 3392
rect 20680 3340 20686 3392
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 25590 3380 25596 3392
rect 22152 3352 25596 3380
rect 22152 3340 22158 3352
rect 25590 3340 25596 3352
rect 25648 3380 25654 3392
rect 26602 3380 26608 3392
rect 25648 3352 26608 3380
rect 25648 3340 25654 3352
rect 26602 3340 26608 3352
rect 26660 3340 26666 3392
rect 27430 3340 27436 3392
rect 27488 3380 27494 3392
rect 29012 3380 29040 3479
rect 27488 3352 29040 3380
rect 27488 3340 27494 3352
rect 552 3290 31648 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 11436 3290
rect 11488 3238 11500 3290
rect 11552 3238 11564 3290
rect 11616 3238 11628 3290
rect 11680 3238 11692 3290
rect 11744 3238 19210 3290
rect 19262 3238 19274 3290
rect 19326 3238 19338 3290
rect 19390 3238 19402 3290
rect 19454 3238 19466 3290
rect 19518 3238 26984 3290
rect 27036 3238 27048 3290
rect 27100 3238 27112 3290
rect 27164 3238 27176 3290
rect 27228 3238 27240 3290
rect 27292 3238 31648 3290
rect 552 3216 31648 3238
rect 6638 3136 6644 3188
rect 6696 3136 6702 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 8202 3176 8208 3188
rect 7616 3148 8208 3176
rect 7616 3136 7622 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9824 3148 10609 3176
rect 9824 3136 9830 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 11204 3148 11253 3176
rect 11204 3136 11210 3148
rect 11241 3145 11253 3148
rect 11287 3145 11299 3179
rect 11241 3139 11299 3145
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 11882 3176 11888 3188
rect 11480 3148 11888 3176
rect 11480 3136 11486 3148
rect 9950 3068 9956 3120
rect 10008 3108 10014 3120
rect 10888 3108 10916 3136
rect 11808 3117 11836 3148
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 14918 3176 14924 3188
rect 12406 3148 14924 3176
rect 11793 3111 11851 3117
rect 10008 3080 11376 3108
rect 10008 3068 10014 3080
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6411 3012 6837 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 9732 3012 10364 3040
rect 9732 3000 9738 3012
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 7098 2981 7104 2984
rect 6273 2975 6331 2981
rect 6273 2972 6285 2975
rect 5684 2944 6285 2972
rect 5684 2932 5690 2944
rect 6273 2941 6285 2944
rect 6319 2972 6331 2975
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 6319 2944 6561 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 7092 2972 7104 2981
rect 7059 2944 7104 2972
rect 6549 2935 6607 2941
rect 7092 2935 7104 2944
rect 7098 2932 7104 2935
rect 7156 2932 7162 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 10137 2975 10195 2981
rect 10137 2972 10149 2975
rect 9916 2944 10149 2972
rect 9916 2932 9922 2944
rect 10137 2941 10149 2944
rect 10183 2941 10195 2975
rect 10137 2935 10195 2941
rect 10226 2932 10232 2984
rect 10284 2932 10290 2984
rect 10336 2981 10364 3012
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 11112 3012 11161 3040
rect 11112 3000 11118 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 10781 2975 10839 2981
rect 10781 2941 10793 2975
rect 10827 2972 10839 2975
rect 10962 2972 10968 2984
rect 10827 2944 10968 2972
rect 10827 2941 10839 2944
rect 10781 2935 10839 2941
rect 9953 2907 10011 2913
rect 9953 2873 9965 2907
rect 9999 2904 10011 2907
rect 10042 2904 10048 2916
rect 9999 2876 10048 2904
rect 9999 2873 10011 2876
rect 9953 2867 10011 2873
rect 10042 2864 10048 2876
rect 10100 2864 10106 2916
rect 10336 2904 10364 2935
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11348 2972 11376 3080
rect 11793 3077 11805 3111
rect 11839 3077 11851 3111
rect 11793 3071 11851 3077
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 11348 2944 11529 2972
rect 11517 2941 11529 2944
rect 11563 2972 11575 2975
rect 11790 2972 11796 2984
rect 11563 2944 11796 2972
rect 11563 2941 11575 2944
rect 11517 2935 11575 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 12406 2972 12434 3148
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 17770 3176 17776 3188
rect 15856 3148 17776 3176
rect 15856 3049 15884 3148
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 22094 3176 22100 3188
rect 21652 3148 22100 3176
rect 16114 3068 16120 3120
rect 16172 3108 16178 3120
rect 21652 3117 21680 3148
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 22833 3179 22891 3185
rect 22833 3176 22845 3179
rect 22244 3148 22845 3176
rect 22244 3136 22250 3148
rect 22833 3145 22845 3148
rect 22879 3145 22891 3179
rect 22833 3139 22891 3145
rect 24397 3179 24455 3185
rect 24397 3145 24409 3179
rect 24443 3176 24455 3179
rect 24854 3176 24860 3188
rect 24443 3148 24860 3176
rect 24443 3145 24455 3148
rect 24397 3139 24455 3145
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 27065 3179 27123 3185
rect 27065 3145 27077 3179
rect 27111 3176 27123 3179
rect 27154 3176 27160 3188
rect 27111 3148 27160 3176
rect 27111 3145 27123 3148
rect 27065 3139 27123 3145
rect 16209 3111 16267 3117
rect 16209 3108 16221 3111
rect 16172 3080 16221 3108
rect 16172 3068 16178 3080
rect 16209 3077 16221 3080
rect 16255 3077 16267 3111
rect 16209 3071 16267 3077
rect 20901 3111 20959 3117
rect 20901 3077 20913 3111
rect 20947 3108 20959 3111
rect 21637 3111 21695 3117
rect 20947 3080 21588 3108
rect 20947 3077 20959 3080
rect 20901 3071 20959 3077
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 21560 3040 21588 3080
rect 21637 3077 21649 3111
rect 21683 3077 21695 3111
rect 21637 3071 21695 3077
rect 25590 3068 25596 3120
rect 25648 3068 25654 3120
rect 27080 3108 27108 3139
rect 27154 3136 27160 3148
rect 27212 3136 27218 3188
rect 27433 3179 27491 3185
rect 27433 3145 27445 3179
rect 27479 3176 27491 3179
rect 27479 3148 29040 3176
rect 27479 3145 27491 3148
rect 27433 3139 27491 3145
rect 26068 3080 27108 3108
rect 21910 3040 21916 3052
rect 15841 3003 15899 3009
rect 16040 3012 16528 3040
rect 21560 3012 21916 3040
rect 16040 2984 16068 3012
rect 11900 2944 12434 2972
rect 11900 2904 11928 2944
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 13538 2972 13544 2984
rect 13228 2944 13544 2972
rect 13228 2932 13234 2944
rect 13538 2932 13544 2944
rect 13596 2972 13602 2984
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 13596 2944 13645 2972
rect 13596 2932 13602 2944
rect 13633 2941 13645 2944
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 15010 2972 15016 2984
rect 14231 2944 15016 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 10336 2876 11100 2904
rect 10505 2839 10563 2845
rect 10505 2805 10517 2839
rect 10551 2836 10563 2839
rect 10870 2836 10876 2848
rect 10551 2808 10876 2836
rect 10551 2805 10563 2808
rect 10505 2799 10563 2805
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 10962 2796 10968 2848
rect 11020 2796 11026 2848
rect 11072 2836 11100 2876
rect 11357 2876 11928 2904
rect 11357 2836 11385 2876
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 14200 2904 14228 2935
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 16022 2932 16028 2984
rect 16080 2932 16086 2984
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2972 16175 2975
rect 16390 2972 16396 2984
rect 16163 2944 16396 2972
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 16500 2981 16528 3012
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 22370 3040 22376 3052
rect 22235 3012 22376 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 22370 3000 22376 3012
rect 22428 3040 22434 3052
rect 25038 3040 25044 3052
rect 22428 3012 25044 3040
rect 22428 3000 22434 3012
rect 25038 3000 25044 3012
rect 25096 3000 25102 3052
rect 26068 3049 26096 3080
rect 27522 3068 27528 3120
rect 27580 3108 27586 3120
rect 27580 3080 28304 3108
rect 27580 3068 27586 3080
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 26510 3000 26516 3052
rect 26568 3040 26574 3052
rect 27341 3043 27399 3049
rect 27341 3040 27353 3043
rect 26568 3012 27353 3040
rect 26568 3000 26574 3012
rect 27341 3009 27353 3012
rect 27387 3040 27399 3043
rect 27430 3040 27436 3052
rect 27387 3012 27436 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 27982 3040 27988 3052
rect 27540 3012 27988 3040
rect 16485 2975 16543 2981
rect 16485 2941 16497 2975
rect 16531 2941 16543 2975
rect 16485 2935 16543 2941
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16816 2944 16865 2972
rect 16816 2932 16822 2944
rect 16853 2941 16865 2944
rect 16899 2972 16911 2975
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 16899 2944 17141 2972
rect 16899 2941 16911 2944
rect 16853 2935 16911 2941
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 17310 2932 17316 2984
rect 17368 2932 17374 2984
rect 19245 2975 19303 2981
rect 19245 2941 19257 2975
rect 19291 2941 19303 2975
rect 19245 2935 19303 2941
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19521 2975 19579 2981
rect 19521 2972 19533 2975
rect 19383 2944 19533 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19521 2941 19533 2944
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 19788 2975 19846 2981
rect 19788 2941 19800 2975
rect 19834 2972 19846 2975
rect 20254 2972 20260 2984
rect 19834 2944 20260 2972
rect 19834 2941 19846 2944
rect 19788 2935 19846 2941
rect 12492 2876 14228 2904
rect 15841 2907 15899 2913
rect 12492 2864 12498 2876
rect 15841 2873 15853 2907
rect 15887 2904 15899 2907
rect 16209 2907 16267 2913
rect 16209 2904 16221 2907
rect 15887 2876 16221 2904
rect 15887 2873 15899 2876
rect 15841 2867 15899 2873
rect 16209 2873 16221 2876
rect 16255 2873 16267 2907
rect 16669 2907 16727 2913
rect 16669 2904 16681 2907
rect 16209 2867 16267 2873
rect 16307 2876 16681 2904
rect 11072 2808 11385 2836
rect 11425 2839 11483 2845
rect 11425 2805 11437 2839
rect 11471 2836 11483 2839
rect 11514 2836 11520 2848
rect 11471 2808 11520 2836
rect 11471 2805 11483 2808
rect 11425 2799 11483 2805
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 11609 2839 11667 2845
rect 11609 2805 11621 2839
rect 11655 2836 11667 2839
rect 11974 2836 11980 2848
rect 11655 2808 11980 2836
rect 11655 2805 11667 2808
rect 11609 2799 11667 2805
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 13078 2796 13084 2848
rect 13136 2836 13142 2848
rect 13814 2836 13820 2848
rect 13136 2808 13820 2836
rect 13136 2796 13142 2808
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14090 2796 14096 2848
rect 14148 2796 14154 2848
rect 15010 2796 15016 2848
rect 15068 2836 15074 2848
rect 16307 2836 16335 2876
rect 16669 2873 16681 2876
rect 16715 2904 16727 2907
rect 17328 2904 17356 2932
rect 16715 2876 17356 2904
rect 19260 2904 19288 2935
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 20990 2932 20996 2984
rect 21048 2932 21054 2984
rect 21177 2975 21235 2981
rect 21177 2941 21189 2975
rect 21223 2941 21235 2975
rect 21177 2935 21235 2941
rect 19610 2904 19616 2916
rect 19260 2876 19616 2904
rect 16715 2873 16727 2876
rect 16669 2867 16727 2873
rect 19610 2864 19616 2876
rect 19668 2864 19674 2916
rect 15068 2808 16335 2836
rect 15068 2796 15074 2808
rect 16390 2796 16396 2848
rect 16448 2836 16454 2848
rect 16942 2836 16948 2848
rect 16448 2808 16948 2836
rect 16448 2796 16454 2808
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17034 2796 17040 2848
rect 17092 2796 17098 2848
rect 17494 2796 17500 2848
rect 17552 2796 17558 2848
rect 21192 2836 21220 2935
rect 22002 2932 22008 2984
rect 22060 2981 22066 2984
rect 22060 2975 22088 2981
rect 22076 2941 22088 2975
rect 22060 2935 22088 2941
rect 22060 2932 22066 2935
rect 23658 2932 23664 2984
rect 23716 2972 23722 2984
rect 25222 2981 25228 2984
rect 24029 2975 24087 2981
rect 24029 2972 24041 2975
rect 23716 2944 24041 2972
rect 23716 2932 23722 2944
rect 24029 2941 24041 2944
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 25200 2975 25228 2981
rect 25200 2941 25212 2975
rect 25200 2935 25228 2941
rect 25222 2932 25228 2935
rect 25280 2932 25286 2984
rect 25314 2932 25320 2984
rect 25372 2932 25378 2984
rect 26234 2932 26240 2984
rect 26292 2932 26298 2984
rect 26694 2932 26700 2984
rect 26752 2932 26758 2984
rect 26786 2932 26792 2984
rect 26844 2932 26850 2984
rect 27062 2932 27068 2984
rect 27120 2972 27126 2984
rect 27540 2981 27568 3012
rect 27982 3000 27988 3012
rect 28040 3000 28046 3052
rect 28276 3049 28304 3080
rect 28261 3043 28319 3049
rect 28261 3009 28273 3043
rect 28307 3040 28319 3043
rect 28445 3043 28503 3049
rect 28445 3040 28457 3043
rect 28307 3012 28457 3040
rect 28307 3009 28319 3012
rect 28261 3003 28319 3009
rect 28445 3009 28457 3012
rect 28491 3009 28503 3043
rect 28445 3003 28503 3009
rect 27525 2975 27583 2981
rect 27525 2972 27537 2975
rect 27120 2944 27537 2972
rect 27120 2932 27126 2944
rect 27525 2941 27537 2944
rect 27571 2941 27583 2975
rect 27525 2935 27583 2941
rect 27617 2975 27675 2981
rect 27617 2941 27629 2975
rect 27663 2972 27675 2975
rect 27709 2975 27767 2981
rect 27709 2972 27721 2975
rect 27663 2944 27721 2972
rect 27663 2941 27675 2944
rect 27617 2935 27675 2941
rect 27709 2941 27721 2944
rect 27755 2941 27767 2975
rect 28000 2972 28028 3000
rect 28629 2975 28687 2981
rect 28629 2972 28641 2975
rect 28000 2944 28641 2972
rect 27709 2935 27767 2941
rect 28629 2941 28641 2944
rect 28675 2941 28687 2975
rect 28629 2935 28687 2941
rect 28810 2932 28816 2984
rect 28868 2932 28874 2984
rect 29012 2981 29040 3148
rect 28997 2975 29055 2981
rect 28997 2941 29009 2975
rect 29043 2941 29055 2975
rect 28997 2935 29055 2941
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29181 2975 29239 2981
rect 29181 2972 29193 2975
rect 29144 2944 29193 2972
rect 29144 2932 29150 2944
rect 29181 2941 29193 2944
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 29457 2975 29515 2981
rect 29457 2941 29469 2975
rect 29503 2972 29515 2975
rect 30926 2972 30932 2984
rect 29503 2944 30932 2972
rect 29503 2941 29515 2944
rect 29457 2935 29515 2941
rect 27249 2907 27307 2913
rect 27249 2873 27261 2907
rect 27295 2904 27307 2907
rect 27338 2904 27344 2916
rect 27295 2876 27344 2904
rect 27295 2873 27307 2876
rect 27249 2867 27307 2873
rect 27338 2864 27344 2876
rect 27396 2864 27402 2916
rect 27430 2864 27436 2916
rect 27488 2904 27494 2916
rect 29472 2904 29500 2935
rect 30926 2932 30932 2944
rect 30984 2932 30990 2984
rect 27488 2876 29500 2904
rect 27488 2864 27494 2876
rect 21634 2836 21640 2848
rect 21192 2808 21640 2836
rect 21634 2796 21640 2808
rect 21692 2836 21698 2848
rect 22186 2836 22192 2848
rect 21692 2808 22192 2836
rect 21692 2796 21698 2808
rect 22186 2796 22192 2808
rect 22244 2796 22250 2848
rect 23750 2796 23756 2848
rect 23808 2836 23814 2848
rect 23937 2839 23995 2845
rect 23937 2836 23949 2839
rect 23808 2808 23949 2836
rect 23808 2796 23814 2808
rect 23937 2805 23949 2808
rect 23983 2805 23995 2839
rect 23937 2799 23995 2805
rect 26513 2839 26571 2845
rect 26513 2805 26525 2839
rect 26559 2836 26571 2839
rect 26694 2836 26700 2848
rect 26559 2808 26700 2836
rect 26559 2805 26571 2808
rect 26513 2799 26571 2805
rect 26694 2796 26700 2808
rect 26752 2796 26758 2848
rect 26878 2796 26884 2848
rect 26936 2796 26942 2848
rect 27062 2845 27068 2848
rect 27049 2839 27068 2845
rect 27049 2805 27061 2839
rect 27049 2799 27068 2805
rect 27062 2796 27068 2799
rect 27120 2796 27126 2848
rect 28810 2796 28816 2848
rect 28868 2836 28874 2848
rect 28994 2836 29000 2848
rect 28868 2808 29000 2836
rect 28868 2796 28874 2808
rect 28994 2796 29000 2808
rect 29052 2796 29058 2848
rect 29086 2796 29092 2848
rect 29144 2796 29150 2848
rect 29362 2796 29368 2848
rect 29420 2796 29426 2848
rect 552 2746 31648 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 12096 2746
rect 12148 2694 12160 2746
rect 12212 2694 12224 2746
rect 12276 2694 12288 2746
rect 12340 2694 12352 2746
rect 12404 2694 19870 2746
rect 19922 2694 19934 2746
rect 19986 2694 19998 2746
rect 20050 2694 20062 2746
rect 20114 2694 20126 2746
rect 20178 2694 27644 2746
rect 27696 2694 27708 2746
rect 27760 2694 27772 2746
rect 27824 2694 27836 2746
rect 27888 2694 27900 2746
rect 27952 2694 31648 2746
rect 552 2672 31648 2694
rect 11238 2632 11244 2644
rect 9600 2604 11244 2632
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 9600 2505 9628 2604
rect 11238 2592 11244 2604
rect 11296 2632 11302 2644
rect 11296 2604 12480 2632
rect 11296 2592 11302 2604
rect 10551 2533 10609 2539
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 9548 2468 9597 2496
rect 9548 2456 9554 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10137 2499 10195 2505
rect 9907 2468 10088 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 10060 2428 10088 2468
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 10226 2496 10232 2508
rect 10183 2468 10232 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 10551 2499 10563 2533
rect 10597 2530 10609 2533
rect 10597 2499 10624 2530
rect 10686 2524 10692 2576
rect 10744 2564 10750 2576
rect 11146 2573 11152 2576
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 10744 2536 10793 2564
rect 10744 2524 10750 2536
rect 10781 2533 10793 2536
rect 10827 2533 10839 2567
rect 10781 2527 10839 2533
rect 11133 2567 11152 2573
rect 11133 2533 11145 2567
rect 11133 2527 11152 2533
rect 11146 2524 11152 2527
rect 11204 2524 11210 2576
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 11379 2536 11560 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 10551 2496 10624 2499
rect 10870 2496 10876 2508
rect 10551 2493 10876 2496
rect 10596 2468 10876 2493
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 11348 2496 11376 2527
rect 11020 2468 11376 2496
rect 11020 2456 11026 2468
rect 10410 2428 10416 2440
rect 10060 2400 10416 2428
rect 10410 2388 10416 2400
rect 10468 2428 10474 2440
rect 10468 2400 11008 2428
rect 10468 2388 10474 2400
rect 10321 2363 10379 2369
rect 10321 2329 10333 2363
rect 10367 2360 10379 2363
rect 10686 2360 10692 2372
rect 10367 2332 10692 2360
rect 10367 2329 10379 2332
rect 10321 2323 10379 2329
rect 10686 2320 10692 2332
rect 10744 2320 10750 2372
rect 10980 2369 11008 2400
rect 10965 2363 11023 2369
rect 10965 2329 10977 2363
rect 11011 2329 11023 2363
rect 10965 2323 11023 2329
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 9364 2264 9505 2292
rect 9364 2252 9370 2264
rect 9493 2261 9505 2264
rect 9539 2261 9551 2295
rect 9493 2255 9551 2261
rect 9766 2252 9772 2304
rect 9824 2252 9830 2304
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 10284 2264 10425 2292
rect 10284 2252 10290 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 10597 2295 10655 2301
rect 10597 2261 10609 2295
rect 10643 2292 10655 2295
rect 11072 2292 11100 2468
rect 11532 2428 11560 2536
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11664 2468 11989 2496
rect 11664 2456 11670 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 12452 2505 12480 2604
rect 15194 2592 15200 2644
rect 15252 2592 15258 2644
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 17000 2604 17693 2632
rect 17000 2592 17006 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 17681 2595 17739 2601
rect 23658 2592 23664 2644
rect 23716 2632 23722 2644
rect 27430 2632 27436 2644
rect 23716 2604 27436 2632
rect 23716 2592 23722 2604
rect 27430 2592 27436 2604
rect 27488 2592 27494 2644
rect 13078 2524 13084 2576
rect 13136 2524 13142 2576
rect 14090 2564 14096 2576
rect 13372 2536 14096 2564
rect 13372 2505 13400 2536
rect 14090 2524 14096 2536
rect 14148 2524 14154 2576
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 15749 2567 15807 2573
rect 15749 2564 15761 2567
rect 14884 2536 15761 2564
rect 14884 2524 14890 2536
rect 15749 2533 15761 2536
rect 15795 2533 15807 2567
rect 15749 2527 15807 2533
rect 15933 2567 15991 2573
rect 15933 2533 15945 2567
rect 15979 2564 15991 2567
rect 17494 2564 17500 2576
rect 15979 2536 17500 2564
rect 15979 2533 15991 2536
rect 15933 2527 15991 2533
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 19794 2524 19800 2576
rect 19852 2564 19858 2576
rect 19852 2536 21956 2564
rect 19852 2524 19858 2536
rect 12437 2499 12495 2505
rect 12437 2496 12449 2499
rect 12400 2468 12449 2496
rect 12400 2456 12406 2468
rect 12437 2465 12449 2468
rect 12483 2465 12495 2499
rect 12437 2459 12495 2465
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2465 13415 2499
rect 13613 2499 13671 2505
rect 13613 2496 13625 2499
rect 13357 2459 13415 2465
rect 13464 2468 13625 2496
rect 11698 2428 11704 2440
rect 11532 2400 11704 2428
rect 11698 2388 11704 2400
rect 11756 2428 11762 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11756 2400 11805 2428
rect 11756 2388 11762 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 12161 2431 12219 2437
rect 12161 2428 12173 2431
rect 12124 2400 12173 2428
rect 12124 2388 12130 2400
rect 12161 2397 12173 2400
rect 12207 2428 12219 2431
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12207 2400 12725 2428
rect 12207 2397 12219 2400
rect 12161 2391 12219 2397
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 13464 2428 13492 2468
rect 13613 2465 13625 2468
rect 13659 2465 13671 2499
rect 13613 2459 13671 2465
rect 13998 2456 14004 2508
rect 14056 2496 14062 2508
rect 15013 2499 15071 2505
rect 15013 2496 15025 2499
rect 14056 2468 15025 2496
rect 14056 2456 14062 2468
rect 12713 2391 12771 2397
rect 13280 2400 13492 2428
rect 11882 2320 11888 2372
rect 11940 2360 11946 2372
rect 13280 2369 13308 2400
rect 12345 2363 12403 2369
rect 12345 2360 12357 2363
rect 11940 2332 12357 2360
rect 11940 2320 11946 2332
rect 12345 2329 12357 2332
rect 12391 2329 12403 2363
rect 12345 2323 12403 2329
rect 13265 2363 13323 2369
rect 13265 2329 13277 2363
rect 13311 2329 13323 2363
rect 14829 2363 14887 2369
rect 14829 2360 14841 2363
rect 13265 2323 13323 2329
rect 14292 2332 14841 2360
rect 10643 2264 11100 2292
rect 10643 2261 10655 2264
rect 10597 2255 10655 2261
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11606 2292 11612 2304
rect 11204 2264 11612 2292
rect 11204 2252 11210 2264
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 13081 2295 13139 2301
rect 13081 2261 13093 2295
rect 13127 2292 13139 2295
rect 14292 2292 14320 2332
rect 14829 2329 14841 2332
rect 14875 2329 14887 2363
rect 14829 2323 14887 2329
rect 13127 2264 14320 2292
rect 14737 2295 14795 2301
rect 13127 2261 13139 2264
rect 13081 2255 13139 2261
rect 14737 2261 14749 2295
rect 14783 2292 14795 2295
rect 14936 2292 14964 2468
rect 15013 2465 15025 2468
rect 15059 2465 15071 2499
rect 15013 2459 15071 2465
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 15378 2496 15384 2508
rect 15335 2468 15384 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 15378 2456 15384 2468
rect 15436 2496 15442 2508
rect 16022 2496 16028 2508
rect 15436 2468 16028 2496
rect 15436 2456 15442 2468
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16206 2456 16212 2508
rect 16264 2456 16270 2508
rect 16465 2499 16523 2505
rect 16465 2496 16477 2499
rect 16316 2468 16477 2496
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16316 2428 16344 2468
rect 16465 2465 16477 2468
rect 16511 2465 16523 2499
rect 16465 2459 16523 2465
rect 18230 2456 18236 2508
rect 18288 2456 18294 2508
rect 19702 2456 19708 2508
rect 19760 2456 19766 2508
rect 19978 2505 19984 2508
rect 19972 2459 19984 2505
rect 19978 2456 19984 2459
rect 20036 2456 20042 2508
rect 20990 2456 20996 2508
rect 21048 2496 21054 2508
rect 21545 2499 21603 2505
rect 21545 2496 21557 2499
rect 21048 2468 21557 2496
rect 21048 2456 21054 2468
rect 21545 2465 21557 2468
rect 21591 2465 21603 2499
rect 21545 2459 21603 2465
rect 21634 2456 21640 2508
rect 21692 2456 21698 2508
rect 21928 2505 21956 2536
rect 24118 2524 24124 2576
rect 24176 2564 24182 2576
rect 26510 2564 26516 2576
rect 24176 2536 26516 2564
rect 24176 2524 24182 2536
rect 26510 2524 26516 2536
rect 26568 2524 26574 2576
rect 26605 2567 26663 2573
rect 26605 2533 26617 2567
rect 26651 2564 26663 2567
rect 26786 2564 26792 2576
rect 26651 2536 26792 2564
rect 26651 2533 26663 2536
rect 26605 2527 26663 2533
rect 26786 2524 26792 2536
rect 26844 2524 26850 2576
rect 28476 2567 28534 2573
rect 28476 2533 28488 2567
rect 28522 2564 28534 2567
rect 29086 2564 29092 2576
rect 28522 2536 29092 2564
rect 28522 2533 28534 2536
rect 28476 2527 28534 2533
rect 29086 2524 29092 2536
rect 29144 2524 29150 2576
rect 21913 2499 21971 2505
rect 21913 2465 21925 2499
rect 21959 2465 21971 2499
rect 21913 2459 21971 2465
rect 22557 2499 22615 2505
rect 22557 2465 22569 2499
rect 22603 2496 22615 2499
rect 22646 2496 22652 2508
rect 22603 2468 22652 2496
rect 22603 2465 22615 2468
rect 22557 2459 22615 2465
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 23750 2456 23756 2508
rect 23808 2456 23814 2508
rect 23842 2456 23848 2508
rect 23900 2496 23906 2508
rect 24009 2499 24067 2505
rect 24009 2496 24021 2499
rect 23900 2468 24021 2496
rect 23900 2456 23906 2468
rect 24009 2465 24021 2468
rect 24055 2465 24067 2499
rect 24009 2459 24067 2465
rect 25222 2456 25228 2508
rect 25280 2496 25286 2508
rect 25501 2499 25559 2505
rect 25501 2496 25513 2499
rect 25280 2468 25513 2496
rect 25280 2456 25286 2468
rect 25501 2465 25513 2468
rect 25547 2465 25559 2499
rect 25501 2459 25559 2465
rect 25593 2499 25651 2505
rect 25593 2465 25605 2499
rect 25639 2496 25651 2499
rect 25774 2496 25780 2508
rect 25639 2468 25780 2496
rect 25639 2465 25651 2468
rect 25593 2459 25651 2465
rect 25774 2456 25780 2468
rect 25832 2496 25838 2508
rect 26234 2496 26240 2508
rect 25832 2468 26240 2496
rect 25832 2456 25838 2468
rect 26234 2456 26240 2468
rect 26292 2456 26298 2508
rect 27154 2456 27160 2508
rect 27212 2496 27218 2508
rect 27338 2496 27344 2508
rect 27212 2468 27344 2496
rect 27212 2456 27218 2468
rect 27338 2456 27344 2468
rect 27396 2456 27402 2508
rect 28721 2499 28779 2505
rect 28721 2465 28733 2499
rect 28767 2496 28779 2499
rect 29362 2496 29368 2508
rect 28767 2468 29368 2496
rect 28767 2465 28779 2468
rect 28721 2459 28779 2465
rect 29362 2456 29368 2468
rect 29420 2456 29426 2508
rect 15988 2400 16344 2428
rect 15988 2388 15994 2400
rect 21450 2388 21456 2440
rect 21508 2388 21514 2440
rect 21729 2431 21787 2437
rect 21729 2397 21741 2431
rect 21775 2428 21787 2431
rect 22002 2428 22008 2440
rect 21775 2400 22008 2428
rect 21775 2397 21787 2400
rect 21729 2391 21787 2397
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 21085 2363 21143 2369
rect 15252 2332 15884 2360
rect 15252 2320 15258 2332
rect 14783 2264 14964 2292
rect 15565 2295 15623 2301
rect 14783 2261 14795 2264
rect 14737 2255 14795 2261
rect 15565 2261 15577 2295
rect 15611 2292 15623 2295
rect 15746 2292 15752 2304
rect 15611 2264 15752 2292
rect 15611 2261 15623 2264
rect 15565 2255 15623 2261
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 15856 2292 15884 2332
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21744 2360 21772 2391
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22278 2388 22284 2440
rect 22336 2388 22342 2440
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25409 2391 25467 2397
rect 25516 2400 25697 2428
rect 21131 2332 21772 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 22094 2320 22100 2372
rect 22152 2360 22158 2372
rect 25133 2363 25191 2369
rect 22152 2332 22508 2360
rect 22152 2320 22158 2332
rect 16574 2292 16580 2304
rect 15856 2264 16580 2292
rect 16574 2252 16580 2264
rect 16632 2252 16638 2304
rect 16850 2252 16856 2304
rect 16908 2292 16914 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 16908 2264 17601 2292
rect 16908 2252 16914 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 21266 2252 21272 2304
rect 21324 2252 21330 2304
rect 21358 2252 21364 2304
rect 21416 2292 21422 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21416 2264 22017 2292
rect 21416 2252 21422 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22370 2252 22376 2304
rect 22428 2252 22434 2304
rect 22480 2301 22508 2332
rect 25133 2329 25145 2363
rect 25179 2360 25191 2363
rect 25314 2360 25320 2372
rect 25179 2332 25320 2360
rect 25179 2329 25191 2332
rect 25133 2323 25191 2329
rect 25314 2320 25320 2332
rect 25372 2320 25378 2372
rect 22465 2295 22523 2301
rect 22465 2261 22477 2295
rect 22511 2292 22523 2295
rect 24394 2292 24400 2304
rect 22511 2264 24400 2292
rect 22511 2261 22523 2264
rect 22465 2255 22523 2261
rect 24394 2252 24400 2264
rect 24452 2252 24458 2304
rect 25222 2252 25228 2304
rect 25280 2252 25286 2304
rect 25424 2292 25452 2391
rect 25516 2372 25544 2400
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 25498 2320 25504 2372
rect 25556 2320 25562 2372
rect 27246 2320 27252 2372
rect 27304 2360 27310 2372
rect 27341 2363 27399 2369
rect 27341 2360 27353 2363
rect 27304 2332 27353 2360
rect 27304 2320 27310 2332
rect 27341 2329 27353 2332
rect 27387 2360 27399 2363
rect 27522 2360 27528 2372
rect 27387 2332 27528 2360
rect 27387 2329 27399 2332
rect 27341 2323 27399 2329
rect 27522 2320 27528 2332
rect 27580 2320 27586 2372
rect 25866 2292 25872 2304
rect 25424 2264 25872 2292
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 552 2202 31648 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 11436 2202
rect 11488 2150 11500 2202
rect 11552 2150 11564 2202
rect 11616 2150 11628 2202
rect 11680 2150 11692 2202
rect 11744 2150 19210 2202
rect 19262 2150 19274 2202
rect 19326 2150 19338 2202
rect 19390 2150 19402 2202
rect 19454 2150 19466 2202
rect 19518 2150 26984 2202
rect 27036 2150 27048 2202
rect 27100 2150 27112 2202
rect 27164 2150 27176 2202
rect 27228 2150 27240 2202
rect 27292 2150 31648 2202
rect 552 2128 31648 2150
rect 9766 2048 9772 2100
rect 9824 2088 9830 2100
rect 9824 2060 11560 2088
rect 9824 2048 9830 2060
rect 10781 2023 10839 2029
rect 10781 1989 10793 2023
rect 10827 2020 10839 2023
rect 11330 2020 11336 2032
rect 10827 1992 11336 2020
rect 10827 1989 10839 1992
rect 10781 1983 10839 1989
rect 11330 1980 11336 1992
rect 11388 1980 11394 2032
rect 9217 1955 9275 1961
rect 9217 1921 9229 1955
rect 9263 1952 9275 1955
rect 9401 1955 9459 1961
rect 9401 1952 9413 1955
rect 9263 1924 9413 1952
rect 9263 1921 9275 1924
rect 9217 1915 9275 1921
rect 9401 1921 9413 1924
rect 9447 1921 9459 1955
rect 11348 1952 11376 1980
rect 9401 1915 9459 1921
rect 11164 1924 11376 1952
rect 9309 1887 9367 1893
rect 9309 1853 9321 1887
rect 9355 1884 9367 1887
rect 9490 1884 9496 1896
rect 9355 1856 9496 1884
rect 9355 1853 9367 1856
rect 9309 1847 9367 1853
rect 9490 1844 9496 1856
rect 9548 1844 9554 1896
rect 11164 1893 11192 1924
rect 11149 1887 11207 1893
rect 11149 1853 11161 1887
rect 11195 1853 11207 1887
rect 11149 1847 11207 1853
rect 11238 1844 11244 1896
rect 11296 1844 11302 1896
rect 11333 1887 11391 1893
rect 11333 1853 11345 1887
rect 11379 1884 11391 1887
rect 11422 1884 11428 1896
rect 11379 1856 11428 1884
rect 11379 1853 11391 1856
rect 11333 1847 11391 1853
rect 11422 1844 11428 1856
rect 11480 1844 11486 1896
rect 11532 1893 11560 2060
rect 11790 2048 11796 2100
rect 11848 2048 11854 2100
rect 12437 2091 12495 2097
rect 12437 2057 12449 2091
rect 12483 2088 12495 2091
rect 12897 2091 12955 2097
rect 12897 2088 12909 2091
rect 12483 2060 12909 2088
rect 12483 2057 12495 2060
rect 12437 2051 12495 2057
rect 12897 2057 12909 2060
rect 12943 2057 12955 2091
rect 12897 2051 12955 2057
rect 14918 2048 14924 2100
rect 14976 2088 14982 2100
rect 15013 2091 15071 2097
rect 15013 2088 15025 2091
rect 14976 2060 15025 2088
rect 14976 2048 14982 2060
rect 15013 2057 15025 2060
rect 15059 2057 15071 2091
rect 15013 2051 15071 2057
rect 15746 2048 15752 2100
rect 15804 2048 15810 2100
rect 15930 2048 15936 2100
rect 15988 2048 15994 2100
rect 16666 2048 16672 2100
rect 16724 2088 16730 2100
rect 16724 2060 16988 2088
rect 16724 2048 16730 2060
rect 11606 1980 11612 2032
rect 11664 1980 11670 2032
rect 12529 2023 12587 2029
rect 12529 2020 12541 2023
rect 11808 1992 12541 2020
rect 11808 1964 11836 1992
rect 12529 1989 12541 1992
rect 12575 1989 12587 2023
rect 12529 1983 12587 1989
rect 15197 2023 15255 2029
rect 15197 1989 15209 2023
rect 15243 2020 15255 2023
rect 15378 2020 15384 2032
rect 15243 1992 15384 2020
rect 15243 1989 15255 1992
rect 15197 1983 15255 1989
rect 15378 1980 15384 1992
rect 15436 1980 15442 2032
rect 16960 2020 16988 2060
rect 17034 2048 17040 2100
rect 17092 2088 17098 2100
rect 17773 2091 17831 2097
rect 17773 2088 17785 2091
rect 17092 2060 17785 2088
rect 17092 2048 17098 2060
rect 17773 2057 17785 2060
rect 17819 2057 17831 2091
rect 17773 2051 17831 2057
rect 19978 2048 19984 2100
rect 20036 2048 20042 2100
rect 20165 2091 20223 2097
rect 20165 2057 20177 2091
rect 20211 2088 20223 2091
rect 20254 2088 20260 2100
rect 20211 2060 20260 2088
rect 20211 2057 20223 2060
rect 20165 2051 20223 2057
rect 20254 2048 20260 2060
rect 20312 2048 20318 2100
rect 20806 2088 20812 2100
rect 20456 2060 20812 2088
rect 17405 2023 17463 2029
rect 17405 2020 17417 2023
rect 16960 1992 17417 2020
rect 17405 1989 17417 1992
rect 17451 1989 17463 2023
rect 17405 1983 17463 1989
rect 11790 1912 11796 1964
rect 11848 1912 11854 1964
rect 11974 1912 11980 1964
rect 12032 1952 12038 1964
rect 12032 1924 12296 1952
rect 12032 1912 12038 1924
rect 11517 1887 11575 1893
rect 11517 1853 11529 1887
rect 11563 1853 11575 1887
rect 11517 1847 11575 1853
rect 11698 1844 11704 1896
rect 11756 1881 11762 1896
rect 11756 1853 11928 1881
rect 11756 1844 11762 1853
rect 9668 1819 9726 1825
rect 9668 1785 9680 1819
rect 9714 1816 9726 1819
rect 10873 1819 10931 1825
rect 10873 1816 10885 1819
rect 9714 1788 10885 1816
rect 9714 1785 9726 1788
rect 9668 1779 9726 1785
rect 10873 1785 10885 1788
rect 10919 1785 10931 1819
rect 11256 1816 11284 1844
rect 11606 1816 11612 1828
rect 11256 1788 11612 1816
rect 10873 1779 10931 1785
rect 11606 1776 11612 1788
rect 11664 1776 11670 1828
rect 10226 1708 10232 1760
rect 10284 1748 10290 1760
rect 11790 1757 11796 1760
rect 11767 1751 11796 1757
rect 11767 1748 11779 1751
rect 10284 1720 11779 1748
rect 10284 1708 10290 1720
rect 11767 1717 11779 1720
rect 11767 1711 11796 1717
rect 11790 1708 11796 1711
rect 11848 1708 11854 1760
rect 11900 1748 11928 1853
rect 12066 1844 12072 1896
rect 12124 1844 12130 1896
rect 12268 1893 12296 1924
rect 12342 1912 12348 1964
rect 12400 1952 12406 1964
rect 12400 1924 13216 1952
rect 12400 1912 12406 1924
rect 12253 1887 12311 1893
rect 12253 1853 12265 1887
rect 12299 1884 12311 1887
rect 12986 1884 12992 1896
rect 12299 1856 12992 1884
rect 12299 1853 12311 1856
rect 12253 1847 12311 1853
rect 12986 1844 12992 1856
rect 13044 1844 13050 1896
rect 13188 1893 13216 1924
rect 13538 1912 13544 1964
rect 13596 1912 13602 1964
rect 17420 1952 17448 1983
rect 17494 1980 17500 2032
rect 17552 2020 17558 2032
rect 18141 2023 18199 2029
rect 18141 2020 18153 2023
rect 17552 1992 18153 2020
rect 17552 1980 17558 1992
rect 18141 1989 18153 1992
rect 18187 1989 18199 2023
rect 18141 1983 18199 1989
rect 19702 1980 19708 2032
rect 19760 2020 19766 2032
rect 19889 2023 19947 2029
rect 19889 2020 19901 2023
rect 19760 1992 19901 2020
rect 19760 1980 19766 1992
rect 19889 1989 19901 1992
rect 19935 1989 19947 2023
rect 20456 2020 20484 2060
rect 20806 2048 20812 2060
rect 20864 2088 20870 2100
rect 21545 2091 21603 2097
rect 20864 2060 21496 2088
rect 20864 2048 20870 2060
rect 21468 2032 21496 2060
rect 21545 2057 21557 2091
rect 21591 2088 21603 2091
rect 22002 2088 22008 2100
rect 21591 2060 22008 2088
rect 21591 2057 21603 2060
rect 21545 2051 21603 2057
rect 22002 2048 22008 2060
rect 22060 2048 22066 2100
rect 22278 2048 22284 2100
rect 22336 2088 22342 2100
rect 22336 2060 22600 2088
rect 22336 2048 22342 2060
rect 19889 1983 19947 1989
rect 19996 1992 20484 2020
rect 20533 2023 20591 2029
rect 18230 1952 18236 1964
rect 17420 1924 18236 1952
rect 18230 1912 18236 1924
rect 18288 1912 18294 1964
rect 19794 1952 19800 1964
rect 19352 1924 19800 1952
rect 13173 1887 13231 1893
rect 13173 1853 13185 1887
rect 13219 1853 13231 1887
rect 13173 1847 13231 1853
rect 13817 1887 13875 1893
rect 13817 1853 13829 1887
rect 13863 1884 13875 1887
rect 13863 1856 15148 1884
rect 13863 1853 13875 1856
rect 13817 1847 13875 1853
rect 11974 1776 11980 1828
rect 12032 1816 12038 1828
rect 12158 1816 12164 1828
rect 12032 1788 12164 1816
rect 12032 1776 12038 1788
rect 12158 1776 12164 1788
rect 12216 1776 12222 1828
rect 12897 1819 12955 1825
rect 12897 1785 12909 1819
rect 12943 1816 12955 1819
rect 13832 1816 13860 1847
rect 12943 1788 13860 1816
rect 12943 1785 12955 1788
rect 12897 1779 12955 1785
rect 12912 1748 12940 1779
rect 14826 1776 14832 1828
rect 14884 1776 14890 1828
rect 15010 1776 15016 1828
rect 15068 1825 15074 1828
rect 15068 1819 15087 1825
rect 15075 1785 15087 1819
rect 15120 1816 15148 1856
rect 16022 1844 16028 1896
rect 16080 1844 16086 1896
rect 16114 1844 16120 1896
rect 16172 1884 16178 1896
rect 16292 1887 16350 1893
rect 16292 1884 16304 1887
rect 16172 1856 16304 1884
rect 16172 1844 16178 1856
rect 16292 1853 16304 1856
rect 16338 1853 16350 1887
rect 17770 1884 17776 1896
rect 16292 1847 16350 1853
rect 16408 1856 17776 1884
rect 16408 1816 16436 1856
rect 17770 1844 17776 1856
rect 17828 1844 17834 1896
rect 19352 1893 19380 1924
rect 19794 1912 19800 1924
rect 19852 1912 19858 1964
rect 18417 1887 18475 1893
rect 18417 1853 18429 1887
rect 18463 1884 18475 1887
rect 19337 1887 19395 1893
rect 19337 1884 19349 1887
rect 18463 1856 19349 1884
rect 18463 1853 18475 1856
rect 18417 1847 18475 1853
rect 19337 1853 19349 1856
rect 19383 1853 19395 1887
rect 19337 1847 19395 1853
rect 19613 1887 19671 1893
rect 19613 1853 19625 1887
rect 19659 1884 19671 1887
rect 19996 1884 20024 1992
rect 20533 1989 20545 2023
rect 20579 2020 20591 2023
rect 20622 2020 20628 2032
rect 20579 1992 20628 2020
rect 20579 1989 20591 1992
rect 20533 1983 20591 1989
rect 20622 1980 20628 1992
rect 20680 2020 20686 2032
rect 21361 2023 21419 2029
rect 21361 2020 21373 2023
rect 20680 1992 21373 2020
rect 20680 1980 20686 1992
rect 21361 1989 21373 1992
rect 21407 1989 21419 2023
rect 21361 1983 21419 1989
rect 21450 1980 21456 2032
rect 21508 2020 21514 2032
rect 21821 2023 21879 2029
rect 21821 2020 21833 2023
rect 21508 1992 21833 2020
rect 21508 1980 21514 1992
rect 21821 1989 21833 1992
rect 21867 2020 21879 2023
rect 22373 2023 22431 2029
rect 22373 2020 22385 2023
rect 21867 1992 22385 2020
rect 21867 1989 21879 1992
rect 21821 1983 21879 1989
rect 22373 1989 22385 1992
rect 22419 1989 22431 2023
rect 22373 1983 22431 1989
rect 22465 2023 22523 2029
rect 22465 1989 22477 2023
rect 22511 1989 22523 2023
rect 22465 1983 22523 1989
rect 22112 1952 22232 1960
rect 22480 1952 22508 1983
rect 22572 1961 22600 2060
rect 22646 2048 22652 2100
rect 22704 2048 22710 2100
rect 24029 2091 24087 2097
rect 24029 2088 24041 2091
rect 23584 2060 24041 2088
rect 20456 1932 22508 1952
rect 20456 1924 22140 1932
rect 22204 1924 22508 1932
rect 22557 1955 22615 1961
rect 20456 1884 20484 1924
rect 22557 1921 22569 1955
rect 22603 1952 22615 1955
rect 23584 1952 23612 2060
rect 24029 2057 24041 2060
rect 24075 2088 24087 2091
rect 24118 2088 24124 2100
rect 24075 2060 24124 2088
rect 24075 2057 24087 2060
rect 24029 2051 24087 2057
rect 24118 2048 24124 2060
rect 24176 2048 24182 2100
rect 24394 2048 24400 2100
rect 24452 2088 24458 2100
rect 25225 2091 25283 2097
rect 25225 2088 25237 2091
rect 24452 2060 25237 2088
rect 24452 2048 24458 2060
rect 25225 2057 25237 2060
rect 25271 2057 25283 2091
rect 25225 2051 25283 2057
rect 25314 2048 25320 2100
rect 25372 2088 25378 2100
rect 25409 2091 25467 2097
rect 25409 2088 25421 2091
rect 25372 2060 25421 2088
rect 25372 2048 25378 2060
rect 25409 2057 25421 2060
rect 25455 2057 25467 2091
rect 25409 2051 25467 2057
rect 25866 2048 25872 2100
rect 25924 2088 25930 2100
rect 26697 2091 26755 2097
rect 26697 2088 26709 2091
rect 25924 2060 26709 2088
rect 25924 2048 25930 2060
rect 26697 2057 26709 2060
rect 26743 2088 26755 2091
rect 26878 2088 26884 2100
rect 26743 2060 26884 2088
rect 26743 2057 26755 2060
rect 26697 2051 26755 2057
rect 26878 2048 26884 2060
rect 26936 2048 26942 2100
rect 27065 2091 27123 2097
rect 27065 2057 27077 2091
rect 27111 2088 27123 2091
rect 27338 2088 27344 2100
rect 27111 2060 27344 2088
rect 27111 2057 27123 2060
rect 27065 2051 27123 2057
rect 27338 2048 27344 2060
rect 27396 2048 27402 2100
rect 23661 2023 23719 2029
rect 23661 1989 23673 2023
rect 23707 2020 23719 2023
rect 23750 2020 23756 2032
rect 23707 1992 23756 2020
rect 23707 1989 23719 1992
rect 23661 1983 23719 1989
rect 23750 1980 23756 1992
rect 23808 1980 23814 2032
rect 23842 1980 23848 2032
rect 23900 1980 23906 2032
rect 23934 1980 23940 2032
rect 23992 2020 23998 2032
rect 24489 2023 24547 2029
rect 24489 2020 24501 2023
rect 23992 1992 24501 2020
rect 23992 1980 23998 1992
rect 24489 1989 24501 1992
rect 24535 2020 24547 2023
rect 24535 1992 26096 2020
rect 24535 1989 24547 1992
rect 24489 1983 24547 1989
rect 22603 1924 23612 1952
rect 23952 1924 25728 1952
rect 22603 1921 22615 1924
rect 22557 1915 22615 1921
rect 19659 1856 20024 1884
rect 20088 1856 20484 1884
rect 19659 1853 19671 1856
rect 19613 1847 19671 1853
rect 15120 1788 16436 1816
rect 15068 1779 15087 1785
rect 15068 1776 15074 1779
rect 16482 1776 16488 1828
rect 16540 1816 16546 1828
rect 18432 1816 18460 1847
rect 16540 1788 18460 1816
rect 19889 1819 19947 1825
rect 16540 1776 16546 1788
rect 19889 1785 19901 1819
rect 19935 1816 19947 1819
rect 20088 1816 20116 1856
rect 20990 1844 20996 1896
rect 21048 1884 21054 1896
rect 21177 1887 21235 1893
rect 21177 1884 21189 1887
rect 21048 1856 21189 1884
rect 21048 1844 21054 1856
rect 21177 1853 21189 1856
rect 21223 1853 21235 1887
rect 22002 1884 22008 1896
rect 21965 1856 22008 1884
rect 21177 1847 21235 1853
rect 22002 1844 22008 1856
rect 22060 1844 22066 1896
rect 22097 1887 22155 1893
rect 22097 1853 22109 1887
rect 22143 1886 22155 1887
rect 22186 1886 22192 1896
rect 22143 1858 22192 1886
rect 22143 1853 22155 1858
rect 22097 1847 22155 1853
rect 22186 1844 22192 1858
rect 22244 1844 22250 1896
rect 22281 1887 22339 1893
rect 22281 1853 22293 1887
rect 22327 1878 22339 1887
rect 22327 1853 22407 1878
rect 22281 1850 22407 1853
rect 22281 1847 22339 1850
rect 19935 1788 20116 1816
rect 20165 1819 20223 1825
rect 19935 1785 19947 1788
rect 19889 1779 19947 1785
rect 20165 1785 20177 1819
rect 20211 1816 20223 1819
rect 21266 1816 21272 1828
rect 20211 1788 21272 1816
rect 20211 1785 20223 1788
rect 20165 1779 20223 1785
rect 21266 1776 21272 1788
rect 21324 1776 21330 1828
rect 21450 1776 21456 1828
rect 21508 1825 21514 1828
rect 21508 1819 21571 1825
rect 21508 1785 21525 1819
rect 21559 1785 21571 1819
rect 21508 1779 21571 1785
rect 21508 1776 21514 1779
rect 21726 1776 21732 1828
rect 21784 1776 21790 1828
rect 11900 1720 12940 1748
rect 13078 1708 13084 1760
rect 13136 1708 13142 1760
rect 13262 1708 13268 1760
rect 13320 1708 13326 1760
rect 13814 1708 13820 1760
rect 13872 1748 13878 1760
rect 15749 1751 15807 1757
rect 15749 1748 15761 1751
rect 13872 1720 15761 1748
rect 13872 1708 13878 1720
rect 15749 1717 15761 1720
rect 15795 1717 15807 1751
rect 15749 1711 15807 1717
rect 17586 1708 17592 1760
rect 17644 1708 17650 1760
rect 17770 1708 17776 1760
rect 17828 1708 17834 1760
rect 18322 1708 18328 1760
rect 18380 1708 18386 1760
rect 19426 1708 19432 1760
rect 19484 1708 19490 1760
rect 19705 1751 19763 1757
rect 19705 1717 19717 1751
rect 19751 1748 19763 1751
rect 20625 1751 20683 1757
rect 20625 1748 20637 1751
rect 19751 1720 20637 1748
rect 19751 1717 19763 1720
rect 19705 1711 19763 1717
rect 20625 1717 20637 1720
rect 20671 1748 20683 1751
rect 22379 1748 22407 1850
rect 23198 1844 23204 1896
rect 23256 1844 23262 1896
rect 23385 1887 23443 1893
rect 23385 1853 23397 1887
rect 23431 1853 23443 1887
rect 23385 1847 23443 1853
rect 23661 1887 23719 1893
rect 23661 1853 23673 1887
rect 23707 1884 23719 1887
rect 23952 1884 23980 1924
rect 23707 1856 23980 1884
rect 23707 1853 23719 1856
rect 23661 1847 23719 1853
rect 20671 1720 22407 1748
rect 23400 1748 23428 1847
rect 24394 1844 24400 1896
rect 24452 1844 24458 1896
rect 25130 1844 25136 1896
rect 25188 1844 25194 1896
rect 25222 1844 25228 1896
rect 25280 1844 25286 1896
rect 23477 1819 23535 1825
rect 23477 1785 23489 1819
rect 23523 1816 23535 1819
rect 23934 1816 23940 1828
rect 23523 1788 23940 1816
rect 23523 1785 23535 1788
rect 23477 1779 23535 1785
rect 23934 1776 23940 1788
rect 23992 1776 23998 1828
rect 24029 1819 24087 1825
rect 24029 1785 24041 1819
rect 24075 1816 24087 1819
rect 25240 1816 25268 1844
rect 24075 1788 25268 1816
rect 24075 1785 24087 1788
rect 24029 1779 24087 1785
rect 25590 1776 25596 1828
rect 25648 1776 25654 1828
rect 25700 1816 25728 1924
rect 25774 1844 25780 1896
rect 25832 1844 25838 1896
rect 25866 1844 25872 1896
rect 25924 1844 25930 1896
rect 26068 1884 26096 1992
rect 26142 1980 26148 2032
rect 26200 2020 26206 2032
rect 26237 2023 26295 2029
rect 26237 2020 26249 2023
rect 26200 1992 26249 2020
rect 26200 1980 26206 1992
rect 26237 1989 26249 1992
rect 26283 1989 26295 2023
rect 26237 1983 26295 1989
rect 26421 1955 26479 1961
rect 26421 1921 26433 1955
rect 26467 1952 26479 1955
rect 26510 1952 26516 1964
rect 26467 1924 26516 1952
rect 26467 1921 26479 1924
rect 26421 1915 26479 1921
rect 26510 1912 26516 1924
rect 26568 1912 26574 1964
rect 26145 1887 26203 1893
rect 26145 1884 26157 1887
rect 26068 1856 26157 1884
rect 26145 1853 26157 1856
rect 26191 1853 26203 1887
rect 26145 1847 26203 1853
rect 26789 1887 26847 1893
rect 26789 1853 26801 1887
rect 26835 1884 26847 1887
rect 27062 1884 27068 1896
rect 26835 1856 27068 1884
rect 26835 1853 26847 1856
rect 26789 1847 26847 1853
rect 27062 1844 27068 1856
rect 27120 1844 27126 1896
rect 28442 1844 28448 1896
rect 28500 1844 28506 1896
rect 26421 1819 26479 1825
rect 26421 1816 26433 1819
rect 25700 1788 26433 1816
rect 26421 1785 26433 1788
rect 26467 1785 26479 1819
rect 26421 1779 26479 1785
rect 27982 1776 27988 1828
rect 28040 1816 28046 1828
rect 28178 1819 28236 1825
rect 28178 1816 28190 1819
rect 28040 1788 28190 1816
rect 28040 1776 28046 1788
rect 28178 1785 28190 1788
rect 28224 1785 28236 1819
rect 28178 1779 28236 1785
rect 25406 1757 25412 1760
rect 25383 1751 25412 1757
rect 25383 1748 25395 1751
rect 23400 1720 25395 1748
rect 20671 1717 20683 1720
rect 20625 1711 20683 1717
rect 25383 1717 25395 1720
rect 25464 1748 25470 1760
rect 26053 1751 26111 1757
rect 26053 1748 26065 1751
rect 25464 1720 26065 1748
rect 25383 1711 25412 1717
rect 25406 1708 25412 1711
rect 25464 1708 25470 1720
rect 26053 1717 26065 1720
rect 26099 1748 26111 1751
rect 26142 1748 26148 1760
rect 26099 1720 26148 1748
rect 26099 1717 26111 1720
rect 26053 1711 26111 1717
rect 26142 1708 26148 1720
rect 26200 1708 26206 1760
rect 26510 1708 26516 1760
rect 26568 1708 26574 1760
rect 552 1658 31648 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 12096 1658
rect 12148 1606 12160 1658
rect 12212 1606 12224 1658
rect 12276 1606 12288 1658
rect 12340 1606 12352 1658
rect 12404 1606 19870 1658
rect 19922 1606 19934 1658
rect 19986 1606 19998 1658
rect 20050 1606 20062 1658
rect 20114 1606 20126 1658
rect 20178 1606 27644 1658
rect 27696 1606 27708 1658
rect 27760 1606 27772 1658
rect 27824 1606 27836 1658
rect 27888 1606 27900 1658
rect 27952 1606 31648 1658
rect 552 1584 31648 1606
rect 9950 1504 9956 1556
rect 10008 1544 10014 1556
rect 10689 1547 10747 1553
rect 10689 1544 10701 1547
rect 10008 1516 10701 1544
rect 10008 1504 10014 1516
rect 10689 1513 10701 1516
rect 10735 1513 10747 1547
rect 10689 1507 10747 1513
rect 11517 1547 11575 1553
rect 11517 1513 11529 1547
rect 11563 1544 11575 1547
rect 11606 1544 11612 1556
rect 11563 1516 11612 1544
rect 11563 1513 11575 1516
rect 11517 1507 11575 1513
rect 11606 1504 11612 1516
rect 11664 1504 11670 1556
rect 11701 1547 11759 1553
rect 11701 1513 11713 1547
rect 11747 1513 11759 1547
rect 11701 1507 11759 1513
rect 11716 1476 11744 1507
rect 11974 1504 11980 1556
rect 12032 1544 12038 1556
rect 13265 1547 13323 1553
rect 13265 1544 13277 1547
rect 12032 1516 13277 1544
rect 12032 1504 12038 1516
rect 13265 1513 13277 1516
rect 13311 1513 13323 1547
rect 13265 1507 13323 1513
rect 16022 1504 16028 1556
rect 16080 1544 16086 1556
rect 16209 1547 16267 1553
rect 16209 1544 16221 1547
rect 16080 1516 16221 1544
rect 16080 1504 16086 1516
rect 16209 1513 16221 1516
rect 16255 1513 16267 1547
rect 16209 1507 16267 1513
rect 16485 1547 16543 1553
rect 16485 1513 16497 1547
rect 16531 1544 16543 1547
rect 16758 1544 16764 1556
rect 16531 1516 16764 1544
rect 16531 1513 16543 1516
rect 16485 1507 16543 1513
rect 12130 1479 12188 1485
rect 12130 1476 12142 1479
rect 11716 1448 12142 1476
rect 12130 1445 12142 1448
rect 12176 1445 12188 1479
rect 12130 1439 12188 1445
rect 13078 1436 13084 1488
rect 13136 1476 13142 1488
rect 13602 1479 13660 1485
rect 13602 1476 13614 1479
rect 13136 1448 13614 1476
rect 13136 1436 13142 1448
rect 13602 1445 13614 1448
rect 13648 1445 13660 1479
rect 13602 1439 13660 1445
rect 14918 1436 14924 1488
rect 14976 1476 14982 1488
rect 16500 1476 16528 1507
rect 16758 1504 16764 1516
rect 16816 1504 16822 1556
rect 19702 1504 19708 1556
rect 19760 1504 19766 1556
rect 20990 1504 20996 1556
rect 21048 1544 21054 1556
rect 21085 1547 21143 1553
rect 21085 1544 21097 1547
rect 21048 1516 21097 1544
rect 21048 1504 21054 1516
rect 21085 1513 21097 1516
rect 21131 1544 21143 1547
rect 21726 1544 21732 1556
rect 21131 1516 21732 1544
rect 21131 1513 21143 1516
rect 21085 1507 21143 1513
rect 21726 1504 21732 1516
rect 21784 1504 21790 1556
rect 22186 1504 22192 1556
rect 22244 1544 22250 1556
rect 22649 1547 22707 1553
rect 22649 1544 22661 1547
rect 22244 1516 22661 1544
rect 22244 1504 22250 1516
rect 22649 1513 22661 1516
rect 22695 1544 22707 1547
rect 23198 1544 23204 1556
rect 22695 1516 23204 1544
rect 22695 1513 22707 1516
rect 22649 1507 22707 1513
rect 23198 1504 23204 1516
rect 23256 1504 23262 1556
rect 25130 1504 25136 1556
rect 25188 1544 25194 1556
rect 25317 1547 25375 1553
rect 25317 1544 25329 1547
rect 25188 1516 25329 1544
rect 25188 1504 25194 1516
rect 25317 1513 25329 1516
rect 25363 1544 25375 1547
rect 25590 1544 25596 1556
rect 25363 1516 25596 1544
rect 25363 1513 25375 1516
rect 25317 1507 25375 1513
rect 25590 1504 25596 1516
rect 25648 1504 25654 1556
rect 27062 1504 27068 1556
rect 27120 1504 27126 1556
rect 27525 1547 27583 1553
rect 27525 1513 27537 1547
rect 27571 1544 27583 1547
rect 28442 1544 28448 1556
rect 27571 1516 28448 1544
rect 27571 1513 27583 1516
rect 27525 1507 27583 1513
rect 28442 1504 28448 1516
rect 28500 1504 28506 1556
rect 14976 1448 16528 1476
rect 14976 1436 14982 1448
rect 17586 1436 17592 1488
rect 17644 1485 17650 1488
rect 17644 1476 17656 1485
rect 19720 1476 19748 1504
rect 19950 1479 20008 1485
rect 19950 1476 19962 1479
rect 17644 1448 17689 1476
rect 19720 1448 19962 1476
rect 17644 1439 17656 1448
rect 19950 1445 19962 1448
rect 19996 1445 20008 1479
rect 19950 1439 20008 1445
rect 17644 1436 17650 1439
rect 20254 1436 20260 1488
rect 20312 1476 20318 1488
rect 22278 1476 22284 1488
rect 20312 1448 22284 1476
rect 20312 1436 20318 1448
rect 22278 1436 22284 1448
rect 22336 1436 22342 1488
rect 23750 1436 23756 1488
rect 23808 1476 23814 1488
rect 24204 1479 24262 1485
rect 24204 1476 24216 1479
rect 23808 1448 24216 1476
rect 23808 1436 23814 1448
rect 24204 1445 24216 1448
rect 24250 1445 24262 1479
rect 24204 1439 24262 1445
rect 26694 1436 26700 1488
rect 26752 1476 26758 1488
rect 26752 1448 27384 1476
rect 26752 1436 26758 1448
rect 9306 1368 9312 1420
rect 9364 1368 9370 1420
rect 9582 1417 9588 1420
rect 9576 1371 9588 1417
rect 9582 1368 9588 1371
rect 9640 1368 9646 1420
rect 11149 1411 11207 1417
rect 11149 1377 11161 1411
rect 11195 1408 11207 1411
rect 11238 1408 11244 1420
rect 11195 1380 11244 1408
rect 11195 1377 11207 1380
rect 11149 1371 11207 1377
rect 11238 1368 11244 1380
rect 11296 1368 11302 1420
rect 11882 1368 11888 1420
rect 11940 1368 11946 1420
rect 13262 1368 13268 1420
rect 13320 1408 13326 1420
rect 13357 1411 13415 1417
rect 13357 1408 13369 1411
rect 13320 1380 13369 1408
rect 13320 1368 13326 1380
rect 13357 1377 13369 1380
rect 13403 1377 13415 1411
rect 13357 1371 13415 1377
rect 16301 1411 16359 1417
rect 16301 1377 16313 1411
rect 16347 1408 16359 1411
rect 16482 1408 16488 1420
rect 16347 1380 16488 1408
rect 16347 1377 16359 1380
rect 16301 1371 16359 1377
rect 16482 1368 16488 1380
rect 16540 1368 16546 1420
rect 19426 1368 19432 1420
rect 19484 1408 19490 1420
rect 19705 1411 19763 1417
rect 19705 1408 19717 1411
rect 19484 1380 19717 1408
rect 19484 1368 19490 1380
rect 19705 1377 19717 1380
rect 19751 1377 19763 1411
rect 19705 1371 19763 1377
rect 21269 1411 21327 1417
rect 21269 1377 21281 1411
rect 21315 1408 21327 1411
rect 21358 1408 21364 1420
rect 21315 1380 21364 1408
rect 21315 1377 21327 1380
rect 21269 1371 21327 1377
rect 21358 1368 21364 1380
rect 21416 1368 21422 1420
rect 21542 1417 21548 1420
rect 21536 1371 21548 1417
rect 21542 1368 21548 1371
rect 21600 1368 21606 1420
rect 23293 1411 23351 1417
rect 23293 1377 23305 1411
rect 23339 1408 23351 1411
rect 23658 1408 23664 1420
rect 23339 1380 23664 1408
rect 23339 1377 23351 1380
rect 23293 1371 23351 1377
rect 23658 1368 23664 1380
rect 23716 1368 23722 1420
rect 25406 1368 25412 1420
rect 25464 1368 25470 1420
rect 25593 1411 25651 1417
rect 25593 1377 25605 1411
rect 25639 1408 25651 1411
rect 26510 1408 26516 1420
rect 25639 1380 26516 1408
rect 25639 1377 25651 1380
rect 25593 1371 25651 1377
rect 26510 1368 26516 1380
rect 26568 1368 26574 1420
rect 26878 1368 26884 1420
rect 26936 1408 26942 1420
rect 27356 1417 27384 1448
rect 27157 1411 27215 1417
rect 27157 1408 27169 1411
rect 26936 1380 27169 1408
rect 26936 1368 26942 1380
rect 27157 1377 27169 1380
rect 27203 1377 27215 1411
rect 27157 1371 27215 1377
rect 27341 1411 27399 1417
rect 27341 1377 27353 1411
rect 27387 1377 27399 1411
rect 27341 1371 27399 1377
rect 27430 1368 27436 1420
rect 27488 1368 27494 1420
rect 17865 1343 17923 1349
rect 17865 1309 17877 1343
rect 17911 1340 17923 1343
rect 18322 1340 18328 1352
rect 17911 1312 18328 1340
rect 17911 1309 17923 1312
rect 17865 1303 17923 1309
rect 18322 1300 18328 1312
rect 18380 1300 18386 1352
rect 23201 1343 23259 1349
rect 23201 1309 23213 1343
rect 23247 1340 23259 1343
rect 23937 1343 23995 1349
rect 23937 1340 23949 1343
rect 23247 1312 23949 1340
rect 23247 1309 23259 1312
rect 23201 1303 23259 1309
rect 23937 1309 23949 1312
rect 23983 1309 23995 1343
rect 23937 1303 23995 1309
rect 26234 1300 26240 1352
rect 26292 1340 26298 1352
rect 26421 1343 26479 1349
rect 26421 1340 26433 1343
rect 26292 1312 26433 1340
rect 26292 1300 26298 1312
rect 26421 1309 26433 1312
rect 26467 1309 26479 1343
rect 26421 1303 26479 1309
rect 27341 1275 27399 1281
rect 27341 1241 27353 1275
rect 27387 1272 27399 1275
rect 27982 1272 27988 1284
rect 27387 1244 27988 1272
rect 27387 1241 27399 1244
rect 27341 1235 27399 1241
rect 27982 1232 27988 1244
rect 28040 1232 28046 1284
rect 11330 1164 11336 1216
rect 11388 1204 11394 1216
rect 11517 1207 11575 1213
rect 11517 1204 11529 1207
rect 11388 1176 11529 1204
rect 11388 1164 11394 1176
rect 11517 1173 11529 1176
rect 11563 1173 11575 1207
rect 11517 1167 11575 1173
rect 12986 1164 12992 1216
rect 13044 1204 13050 1216
rect 14737 1207 14795 1213
rect 14737 1204 14749 1207
rect 13044 1176 14749 1204
rect 13044 1164 13050 1176
rect 14737 1173 14749 1176
rect 14783 1173 14795 1207
rect 14737 1167 14795 1173
rect 25590 1164 25596 1216
rect 25648 1164 25654 1216
rect 552 1114 31648 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 11436 1114
rect 11488 1062 11500 1114
rect 11552 1062 11564 1114
rect 11616 1062 11628 1114
rect 11680 1062 11692 1114
rect 11744 1062 19210 1114
rect 19262 1062 19274 1114
rect 19326 1062 19338 1114
rect 19390 1062 19402 1114
rect 19454 1062 19466 1114
rect 19518 1062 26984 1114
rect 27036 1062 27048 1114
rect 27100 1062 27112 1114
rect 27164 1062 27176 1114
rect 27228 1062 27240 1114
rect 27292 1062 31648 1114
rect 552 1040 31648 1062
rect 9582 960 9588 1012
rect 9640 1000 9646 1012
rect 10505 1003 10563 1009
rect 10505 1000 10517 1003
rect 9640 972 10517 1000
rect 9640 960 9646 972
rect 10505 969 10517 972
rect 10551 969 10563 1003
rect 10505 963 10563 969
rect 11330 960 11336 1012
rect 11388 960 11394 1012
rect 20993 1003 21051 1009
rect 20993 969 21005 1003
rect 21039 1000 21051 1003
rect 21542 1000 21548 1012
rect 21039 972 21548 1000
rect 21039 969 21051 972
rect 20993 963 21051 969
rect 21542 960 21548 972
rect 21600 960 21606 1012
rect 25685 1003 25743 1009
rect 25685 969 25697 1003
rect 25731 1000 25743 1003
rect 26234 1000 26240 1012
rect 25731 972 26240 1000
rect 25731 969 25743 972
rect 25685 963 25743 969
rect 26234 960 26240 972
rect 26292 960 26298 1012
rect 10226 892 10232 944
rect 10284 892 10290 944
rect 9398 824 9404 876
rect 9456 864 9462 876
rect 10413 867 10471 873
rect 10413 864 10425 867
rect 9456 836 10425 864
rect 9456 824 9462 836
rect 10413 833 10425 836
rect 10459 864 10471 867
rect 13814 864 13820 876
rect 10459 836 13820 864
rect 10459 833 10471 836
rect 10413 827 10471 833
rect 13814 824 13820 836
rect 13872 824 13878 876
rect 9950 756 9956 808
rect 10008 796 10014 808
rect 10137 799 10195 805
rect 10137 796 10149 799
rect 10008 768 10149 796
rect 10008 756 10014 768
rect 10137 765 10149 768
rect 10183 765 10195 799
rect 10505 799 10563 805
rect 10505 796 10517 799
rect 10137 759 10195 765
rect 10428 768 10517 796
rect 10428 737 10456 768
rect 10505 765 10517 768
rect 10551 765 10563 799
rect 10505 759 10563 765
rect 10686 756 10692 808
rect 10744 796 10750 808
rect 10965 799 11023 805
rect 10965 796 10977 799
rect 10744 768 10977 796
rect 10744 756 10750 768
rect 10965 765 10977 768
rect 11011 765 11023 799
rect 10965 759 11023 765
rect 11149 799 11207 805
rect 11149 765 11161 799
rect 11195 796 11207 799
rect 11974 796 11980 808
rect 11195 768 11980 796
rect 11195 765 11207 768
rect 11149 759 11207 765
rect 11974 756 11980 768
rect 12032 756 12038 808
rect 20806 756 20812 808
rect 20864 756 20870 808
rect 20993 799 21051 805
rect 20993 765 21005 799
rect 21039 796 21051 799
rect 22370 796 22376 808
rect 21039 768 22376 796
rect 21039 765 21051 768
rect 20993 759 21051 765
rect 22370 756 22376 768
rect 22428 756 22434 808
rect 23658 756 23664 808
rect 23716 796 23722 808
rect 24029 799 24087 805
rect 24029 796 24041 799
rect 23716 768 24041 796
rect 23716 756 23722 768
rect 24029 765 24041 768
rect 24075 765 24087 799
rect 24029 759 24087 765
rect 24121 799 24179 805
rect 24121 765 24133 799
rect 24167 796 24179 799
rect 24305 799 24363 805
rect 24305 796 24317 799
rect 24167 768 24317 796
rect 24167 765 24179 768
rect 24121 759 24179 765
rect 24305 765 24317 768
rect 24351 765 24363 799
rect 24305 759 24363 765
rect 24572 799 24630 805
rect 24572 765 24584 799
rect 24618 796 24630 799
rect 25590 796 25596 808
rect 24618 768 25596 796
rect 24618 765 24630 768
rect 24572 759 24630 765
rect 25590 756 25596 768
rect 25648 756 25654 808
rect 10413 731 10471 737
rect 10413 697 10425 731
rect 10459 697 10471 731
rect 10413 691 10471 697
rect 552 570 31648 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 12096 570
rect 12148 518 12160 570
rect 12212 518 12224 570
rect 12276 518 12288 570
rect 12340 518 12352 570
rect 12404 518 19870 570
rect 19922 518 19934 570
rect 19986 518 19998 570
rect 20050 518 20062 570
rect 20114 518 20126 570
rect 20178 518 27644 570
rect 27696 518 27708 570
rect 27760 518 27772 570
rect 27824 518 27836 570
rect 27888 518 27900 570
rect 27952 518 31648 570
rect 552 496 31648 518
<< via1 >>
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 11436 21734 11488 21786
rect 11500 21734 11552 21786
rect 11564 21734 11616 21786
rect 11628 21734 11680 21786
rect 11692 21734 11744 21786
rect 19210 21734 19262 21786
rect 19274 21734 19326 21786
rect 19338 21734 19390 21786
rect 19402 21734 19454 21786
rect 19466 21734 19518 21786
rect 26984 21734 27036 21786
rect 27048 21734 27100 21786
rect 27112 21734 27164 21786
rect 27176 21734 27228 21786
rect 27240 21734 27292 21786
rect 6460 21675 6512 21684
rect 6460 21641 6469 21675
rect 6469 21641 6503 21675
rect 6503 21641 6512 21675
rect 6460 21632 6512 21641
rect 7288 21675 7340 21684
rect 7288 21641 7297 21675
rect 7297 21641 7331 21675
rect 7331 21641 7340 21675
rect 7288 21632 7340 21641
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 8668 21675 8720 21684
rect 8668 21641 8677 21675
rect 8677 21641 8711 21675
rect 8711 21641 8720 21675
rect 8668 21632 8720 21641
rect 9956 21632 10008 21684
rect 10324 21675 10376 21684
rect 10324 21641 10333 21675
rect 10333 21641 10367 21675
rect 10367 21641 10376 21675
rect 10324 21632 10376 21641
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 27528 21632 27580 21684
rect 3332 21564 3384 21616
rect 4068 21564 4120 21616
rect 26884 21564 26936 21616
rect 2688 21428 2740 21480
rect 3240 21471 3292 21480
rect 3240 21437 3249 21471
rect 3249 21437 3283 21471
rect 3283 21437 3292 21471
rect 3240 21428 3292 21437
rect 3332 21471 3384 21480
rect 3332 21437 3341 21471
rect 3341 21437 3375 21471
rect 3375 21437 3384 21471
rect 3332 21428 3384 21437
rect 3516 21539 3568 21548
rect 3516 21505 3525 21539
rect 3525 21505 3559 21539
rect 3559 21505 3568 21539
rect 3516 21496 3568 21505
rect 4068 21471 4120 21480
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 4252 21471 4304 21480
rect 4252 21437 4261 21471
rect 4261 21437 4295 21471
rect 4295 21437 4304 21471
rect 4252 21428 4304 21437
rect 8024 21496 8076 21548
rect 6460 21428 6512 21480
rect 8300 21428 8352 21480
rect 2412 21360 2464 21412
rect 3424 21360 3476 21412
rect 2504 21292 2556 21344
rect 2780 21292 2832 21344
rect 4068 21335 4120 21344
rect 4068 21301 4077 21335
rect 4077 21301 4111 21335
rect 4111 21301 4120 21335
rect 4068 21292 4120 21301
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 6828 21292 6880 21344
rect 7012 21292 7064 21344
rect 9864 21471 9916 21480
rect 9864 21437 9873 21471
rect 9873 21437 9907 21471
rect 9907 21437 9916 21471
rect 9864 21428 9916 21437
rect 9772 21360 9824 21412
rect 10508 21471 10560 21480
rect 10508 21437 10517 21471
rect 10517 21437 10551 21471
rect 10551 21437 10560 21471
rect 10508 21428 10560 21437
rect 11336 21471 11388 21480
rect 11336 21437 11345 21471
rect 11345 21437 11379 21471
rect 11379 21437 11388 21471
rect 11336 21428 11388 21437
rect 13728 21428 13780 21480
rect 16580 21428 16632 21480
rect 16672 21471 16724 21480
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 18604 21428 18656 21480
rect 19432 21428 19484 21480
rect 17592 21360 17644 21412
rect 19248 21403 19300 21412
rect 19248 21369 19257 21403
rect 19257 21369 19291 21403
rect 19291 21369 19300 21403
rect 19248 21360 19300 21369
rect 19800 21471 19852 21480
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 21548 21428 21600 21480
rect 21640 21471 21692 21480
rect 21640 21437 21649 21471
rect 21649 21437 21683 21471
rect 21683 21437 21692 21471
rect 21640 21428 21692 21437
rect 23848 21471 23900 21480
rect 23848 21437 23857 21471
rect 23857 21437 23891 21471
rect 23891 21437 23900 21471
rect 23848 21428 23900 21437
rect 24400 21471 24452 21480
rect 24400 21437 24409 21471
rect 24409 21437 24443 21471
rect 24443 21437 24452 21471
rect 24400 21428 24452 21437
rect 24952 21471 25004 21480
rect 24952 21437 24961 21471
rect 24961 21437 24995 21471
rect 24995 21437 25004 21471
rect 24952 21428 25004 21437
rect 25504 21471 25556 21480
rect 25504 21437 25513 21471
rect 25513 21437 25547 21471
rect 25547 21437 25556 21471
rect 25504 21428 25556 21437
rect 26516 21496 26568 21548
rect 26056 21471 26108 21480
rect 26056 21437 26065 21471
rect 26065 21437 26099 21471
rect 26099 21437 26108 21471
rect 26056 21428 26108 21437
rect 29000 21539 29052 21548
rect 29000 21505 29009 21539
rect 29009 21505 29043 21539
rect 29043 21505 29052 21539
rect 29000 21496 29052 21505
rect 9956 21292 10008 21344
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 12808 21292 12860 21344
rect 15568 21335 15620 21344
rect 15568 21301 15577 21335
rect 15577 21301 15611 21335
rect 15611 21301 15620 21335
rect 15568 21292 15620 21301
rect 15752 21292 15804 21344
rect 16764 21292 16816 21344
rect 17776 21292 17828 21344
rect 18512 21292 18564 21344
rect 20260 21360 20312 21412
rect 19616 21292 19668 21344
rect 19708 21335 19760 21344
rect 19708 21301 19717 21335
rect 19717 21301 19751 21335
rect 19751 21301 19760 21335
rect 19708 21292 19760 21301
rect 21824 21335 21876 21344
rect 21824 21301 21833 21335
rect 21833 21301 21867 21335
rect 21867 21301 21876 21335
rect 21824 21292 21876 21301
rect 24032 21335 24084 21344
rect 24032 21301 24041 21335
rect 24041 21301 24075 21335
rect 24075 21301 24084 21335
rect 24032 21292 24084 21301
rect 24584 21335 24636 21344
rect 24584 21301 24593 21335
rect 24593 21301 24627 21335
rect 24627 21301 24636 21335
rect 24584 21292 24636 21301
rect 25136 21335 25188 21344
rect 25136 21301 25145 21335
rect 25145 21301 25179 21335
rect 25179 21301 25188 21335
rect 25136 21292 25188 21301
rect 28264 21471 28316 21480
rect 28264 21437 28273 21471
rect 28273 21437 28307 21471
rect 28307 21437 28316 21471
rect 28264 21428 28316 21437
rect 29184 21428 29236 21480
rect 26240 21335 26292 21344
rect 26240 21301 26249 21335
rect 26249 21301 26283 21335
rect 26283 21301 26292 21335
rect 26240 21292 26292 21301
rect 26516 21335 26568 21344
rect 26516 21301 26525 21335
rect 26525 21301 26559 21335
rect 26559 21301 26568 21335
rect 26516 21292 26568 21301
rect 27988 21292 28040 21344
rect 28172 21335 28224 21344
rect 28172 21301 28181 21335
rect 28181 21301 28215 21335
rect 28215 21301 28224 21335
rect 28172 21292 28224 21301
rect 30472 21292 30524 21344
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 12096 21190 12148 21242
rect 12160 21190 12212 21242
rect 12224 21190 12276 21242
rect 12288 21190 12340 21242
rect 12352 21190 12404 21242
rect 19870 21190 19922 21242
rect 19934 21190 19986 21242
rect 19998 21190 20050 21242
rect 20062 21190 20114 21242
rect 20126 21190 20178 21242
rect 27644 21190 27696 21242
rect 27708 21190 27760 21242
rect 27772 21190 27824 21242
rect 27836 21190 27888 21242
rect 27900 21190 27952 21242
rect 3240 21088 3292 21140
rect 3976 21088 4028 21140
rect 6276 21131 6328 21140
rect 6276 21097 6285 21131
rect 6285 21097 6319 21131
rect 6319 21097 6328 21131
rect 6276 21088 6328 21097
rect 8300 21088 8352 21140
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 9864 21088 9916 21140
rect 13820 21088 13872 21140
rect 16672 21088 16724 21140
rect 3516 21020 3568 21072
rect 5356 21020 5408 21072
rect 2320 20952 2372 21004
rect 2412 20995 2464 21004
rect 2412 20961 2421 20995
rect 2421 20961 2455 20995
rect 2455 20961 2464 20995
rect 2412 20952 2464 20961
rect 2504 20995 2556 21004
rect 2504 20961 2513 20995
rect 2513 20961 2547 20995
rect 2547 20961 2556 20995
rect 2504 20952 2556 20961
rect 4068 20952 4120 21004
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 4620 20995 4672 21004
rect 4620 20961 4629 20995
rect 4629 20961 4663 20995
rect 4663 20961 4672 20995
rect 4620 20952 4672 20961
rect 6184 21020 6236 21072
rect 6460 20995 6512 21004
rect 6460 20961 6469 20995
rect 6469 20961 6503 20995
rect 6503 20961 6512 20995
rect 6460 20952 6512 20961
rect 11704 21063 11756 21072
rect 11704 21029 11713 21063
rect 11713 21029 11747 21063
rect 11747 21029 11756 21063
rect 11704 21020 11756 21029
rect 17684 21020 17736 21072
rect 6828 20995 6880 21004
rect 6828 20961 6862 20995
rect 6862 20961 6880 20995
rect 6828 20952 6880 20961
rect 8300 20995 8352 21004
rect 8300 20961 8309 20995
rect 8309 20961 8343 20995
rect 8343 20961 8352 20995
rect 8300 20952 8352 20961
rect 8392 20952 8444 21004
rect 8208 20884 8260 20936
rect 10232 20952 10284 21004
rect 12072 20995 12124 21004
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 10324 20884 10376 20936
rect 11336 20884 11388 20936
rect 12808 20995 12860 21004
rect 12808 20961 12817 20995
rect 12817 20961 12851 20995
rect 12851 20961 12860 20995
rect 12808 20952 12860 20961
rect 13728 20952 13780 21004
rect 15292 20995 15344 21004
rect 15292 20961 15301 20995
rect 15301 20961 15335 20995
rect 15335 20961 15344 20995
rect 15292 20952 15344 20961
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 15752 20995 15804 21004
rect 15752 20961 15761 20995
rect 15761 20961 15795 20995
rect 15795 20961 15804 20995
rect 15752 20952 15804 20961
rect 16580 20952 16632 21004
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 17960 20952 18012 21004
rect 18236 20995 18288 21004
rect 18236 20961 18245 20995
rect 18245 20961 18279 20995
rect 18279 20961 18288 20995
rect 18236 20952 18288 20961
rect 19248 21088 19300 21140
rect 19892 21088 19944 21140
rect 21548 21020 21600 21072
rect 18512 20995 18564 21004
rect 18512 20961 18521 20995
rect 18521 20961 18555 20995
rect 18555 20961 18564 20995
rect 18512 20952 18564 20961
rect 19708 20952 19760 21004
rect 21824 20952 21876 21004
rect 24032 21020 24084 21072
rect 24584 20952 24636 21004
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 18972 20927 19024 20936
rect 18972 20893 18981 20927
rect 18981 20893 19015 20927
rect 19015 20893 19024 20927
rect 18972 20884 19024 20893
rect 26240 21020 26292 21072
rect 28172 21020 28224 21072
rect 30472 20995 30524 21004
rect 30472 20961 30490 20995
rect 30490 20961 30524 20995
rect 30472 20952 30524 20961
rect 25780 20884 25832 20936
rect 27804 20927 27856 20936
rect 27804 20893 27813 20927
rect 27813 20893 27847 20927
rect 27847 20893 27856 20927
rect 27804 20884 27856 20893
rect 29276 20927 29328 20936
rect 29276 20893 29285 20927
rect 29285 20893 29319 20927
rect 29319 20893 29328 20927
rect 29276 20884 29328 20893
rect 2228 20748 2280 20800
rect 2688 20748 2740 20800
rect 12900 20816 12952 20868
rect 13820 20816 13872 20868
rect 5448 20791 5500 20800
rect 5448 20757 5457 20791
rect 5457 20757 5491 20791
rect 5491 20757 5500 20791
rect 5448 20748 5500 20757
rect 6276 20748 6328 20800
rect 8668 20791 8720 20800
rect 8668 20757 8677 20791
rect 8677 20757 8711 20791
rect 8711 20757 8720 20791
rect 8668 20748 8720 20757
rect 13728 20791 13780 20800
rect 13728 20757 13737 20791
rect 13737 20757 13771 20791
rect 13771 20757 13780 20791
rect 13728 20748 13780 20757
rect 15752 20748 15804 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 17868 20791 17920 20800
rect 17868 20757 17877 20791
rect 17877 20757 17911 20791
rect 17911 20757 17920 20791
rect 17868 20748 17920 20757
rect 20812 20748 20864 20800
rect 22652 20748 22704 20800
rect 24216 20791 24268 20800
rect 24216 20757 24225 20791
rect 24225 20757 24259 20791
rect 24259 20757 24268 20791
rect 24216 20748 24268 20757
rect 26424 20791 26476 20800
rect 26424 20757 26433 20791
rect 26433 20757 26467 20791
rect 26467 20757 26476 20791
rect 26424 20748 26476 20757
rect 28080 20748 28132 20800
rect 29368 20791 29420 20800
rect 29368 20757 29377 20791
rect 29377 20757 29411 20791
rect 29411 20757 29420 20791
rect 29368 20748 29420 20757
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 11436 20646 11488 20698
rect 11500 20646 11552 20698
rect 11564 20646 11616 20698
rect 11628 20646 11680 20698
rect 11692 20646 11744 20698
rect 19210 20646 19262 20698
rect 19274 20646 19326 20698
rect 19338 20646 19390 20698
rect 19402 20646 19454 20698
rect 19466 20646 19518 20698
rect 26984 20646 27036 20698
rect 27048 20646 27100 20698
rect 27112 20646 27164 20698
rect 27176 20646 27228 20698
rect 27240 20646 27292 20698
rect 2320 20544 2372 20596
rect 4252 20544 4304 20596
rect 8576 20587 8628 20596
rect 8576 20553 8585 20587
rect 8585 20553 8619 20587
rect 8619 20553 8628 20587
rect 8576 20544 8628 20553
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 12072 20544 12124 20596
rect 16948 20587 17000 20596
rect 16948 20553 16957 20587
rect 16957 20553 16991 20587
rect 16991 20553 17000 20587
rect 16948 20544 17000 20553
rect 17500 20544 17552 20596
rect 20260 20587 20312 20596
rect 20260 20553 20269 20587
rect 20269 20553 20303 20587
rect 20303 20553 20312 20587
rect 20260 20544 20312 20553
rect 18052 20476 18104 20528
rect 4436 20408 4488 20460
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 3332 20340 3384 20392
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 5080 20408 5132 20460
rect 5448 20408 5500 20460
rect 6000 20408 6052 20460
rect 13728 20408 13780 20460
rect 15568 20408 15620 20460
rect 15844 20408 15896 20460
rect 18604 20476 18656 20528
rect 4620 20383 4672 20392
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 4804 20340 4856 20392
rect 4988 20383 5040 20392
rect 4988 20349 4997 20383
rect 4997 20349 5031 20383
rect 5031 20349 5040 20383
rect 4988 20340 5040 20349
rect 8024 20383 8076 20392
rect 8024 20349 8033 20383
rect 8033 20349 8067 20383
rect 8067 20349 8076 20383
rect 8024 20340 8076 20349
rect 8300 20340 8352 20392
rect 8944 20383 8996 20392
rect 8944 20349 8953 20383
rect 8953 20349 8987 20383
rect 8987 20349 8996 20383
rect 8944 20340 8996 20349
rect 10140 20340 10192 20392
rect 12624 20340 12676 20392
rect 13636 20340 13688 20392
rect 13820 20383 13872 20392
rect 13820 20349 13829 20383
rect 13829 20349 13863 20383
rect 13863 20349 13872 20383
rect 13820 20340 13872 20349
rect 15660 20383 15712 20392
rect 15660 20349 15669 20383
rect 15669 20349 15703 20383
rect 15703 20349 15712 20383
rect 15660 20340 15712 20349
rect 16764 20340 16816 20392
rect 3240 20272 3292 20324
rect 1952 20204 2004 20256
rect 3332 20204 3384 20256
rect 4896 20204 4948 20256
rect 7012 20272 7064 20324
rect 11060 20272 11112 20324
rect 17592 20383 17644 20392
rect 17592 20349 17601 20383
rect 17601 20349 17635 20383
rect 17635 20349 17644 20383
rect 17592 20340 17644 20349
rect 18880 20408 18932 20460
rect 18236 20383 18288 20392
rect 18236 20349 18245 20383
rect 18245 20349 18279 20383
rect 18279 20349 18288 20383
rect 18236 20340 18288 20349
rect 18328 20383 18380 20392
rect 18328 20349 18337 20383
rect 18337 20349 18371 20383
rect 18371 20349 18380 20383
rect 18328 20340 18380 20349
rect 18420 20340 18472 20392
rect 8484 20204 8536 20256
rect 13360 20204 13412 20256
rect 15200 20204 15252 20256
rect 16028 20204 16080 20256
rect 17040 20204 17092 20256
rect 17776 20204 17828 20256
rect 19064 20340 19116 20392
rect 19432 20340 19484 20392
rect 19800 20340 19852 20392
rect 20260 20340 20312 20392
rect 20904 20383 20956 20392
rect 20904 20349 20913 20383
rect 20913 20349 20947 20383
rect 20947 20349 20956 20383
rect 20904 20340 20956 20349
rect 29368 20544 29420 20596
rect 22468 20408 22520 20460
rect 22744 20408 22796 20460
rect 22376 20340 22428 20392
rect 19708 20272 19760 20324
rect 22100 20315 22152 20324
rect 22100 20281 22109 20315
rect 22109 20281 22143 20315
rect 22143 20281 22152 20315
rect 22100 20272 22152 20281
rect 22192 20315 22244 20324
rect 22192 20281 22201 20315
rect 22201 20281 22235 20315
rect 22235 20281 22244 20315
rect 22192 20272 22244 20281
rect 19340 20204 19392 20256
rect 19616 20204 19668 20256
rect 19892 20204 19944 20256
rect 20260 20204 20312 20256
rect 22468 20247 22520 20256
rect 22468 20213 22477 20247
rect 22477 20213 22511 20247
rect 22511 20213 22520 20247
rect 22468 20204 22520 20213
rect 22928 20383 22980 20392
rect 22928 20349 22937 20383
rect 22937 20349 22971 20383
rect 22971 20349 22980 20383
rect 22928 20340 22980 20349
rect 23756 20340 23808 20392
rect 25136 20340 25188 20392
rect 25780 20383 25832 20392
rect 25780 20349 25789 20383
rect 25789 20349 25823 20383
rect 25823 20349 25832 20383
rect 25780 20340 25832 20349
rect 27804 20340 27856 20392
rect 29276 20383 29328 20392
rect 29276 20349 29285 20383
rect 29285 20349 29319 20383
rect 29319 20349 29328 20383
rect 29276 20340 29328 20349
rect 26516 20272 26568 20324
rect 26884 20272 26936 20324
rect 29460 20272 29512 20324
rect 22928 20204 22980 20256
rect 23480 20204 23532 20256
rect 24124 20204 24176 20256
rect 25872 20247 25924 20256
rect 25872 20213 25881 20247
rect 25881 20213 25915 20247
rect 25915 20213 25924 20247
rect 25872 20204 25924 20213
rect 29552 20204 29604 20256
rect 29644 20204 29696 20256
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 12096 20102 12148 20154
rect 12160 20102 12212 20154
rect 12224 20102 12276 20154
rect 12288 20102 12340 20154
rect 12352 20102 12404 20154
rect 19870 20102 19922 20154
rect 19934 20102 19986 20154
rect 19998 20102 20050 20154
rect 20062 20102 20114 20154
rect 20126 20102 20178 20154
rect 27644 20102 27696 20154
rect 27708 20102 27760 20154
rect 27772 20102 27824 20154
rect 27836 20102 27888 20154
rect 27900 20102 27952 20154
rect 4988 20000 5040 20052
rect 5356 20000 5408 20052
rect 7104 20000 7156 20052
rect 8392 20000 8444 20052
rect 8944 20000 8996 20052
rect 10232 20000 10284 20052
rect 11060 20043 11112 20052
rect 11060 20009 11069 20043
rect 11069 20009 11103 20043
rect 11103 20009 11112 20043
rect 11060 20000 11112 20009
rect 14740 20000 14792 20052
rect 15476 20000 15528 20052
rect 2412 19932 2464 19984
rect 4712 19932 4764 19984
rect 1952 19907 2004 19916
rect 1952 19873 1961 19907
rect 1961 19873 1995 19907
rect 1995 19873 2004 19907
rect 1952 19864 2004 19873
rect 3424 19907 3476 19916
rect 3424 19873 3433 19907
rect 3433 19873 3467 19907
rect 3467 19873 3476 19907
rect 3424 19864 3476 19873
rect 3516 19864 3568 19916
rect 5356 19864 5408 19916
rect 7196 19932 7248 19984
rect 8208 19932 8260 19984
rect 8668 19932 8720 19984
rect 6000 19907 6052 19916
rect 6000 19873 6009 19907
rect 6009 19873 6043 19907
rect 6043 19873 6052 19907
rect 6000 19864 6052 19873
rect 4804 19796 4856 19848
rect 6276 19907 6328 19916
rect 6276 19873 6285 19907
rect 6285 19873 6319 19907
rect 6319 19873 6328 19907
rect 6276 19864 6328 19873
rect 6460 19864 6512 19916
rect 7656 19864 7708 19916
rect 8024 19864 8076 19916
rect 8484 19864 8536 19916
rect 11060 19864 11112 19916
rect 11888 19932 11940 19984
rect 15292 19932 15344 19984
rect 15568 19975 15620 19984
rect 15568 19941 15577 19975
rect 15577 19941 15611 19975
rect 15611 19941 15620 19975
rect 15568 19932 15620 19941
rect 15936 19932 15988 19984
rect 16580 20000 16632 20052
rect 17684 20000 17736 20052
rect 17960 20000 18012 20052
rect 18420 20000 18472 20052
rect 18972 20000 19024 20052
rect 4896 19728 4948 19780
rect 6000 19728 6052 19780
rect 4068 19660 4120 19712
rect 4160 19660 4212 19712
rect 7012 19796 7064 19848
rect 7196 19839 7248 19848
rect 7196 19805 7205 19839
rect 7205 19805 7239 19839
rect 7239 19805 7248 19839
rect 7196 19796 7248 19805
rect 6552 19728 6604 19780
rect 11244 19796 11296 19848
rect 11152 19728 11204 19780
rect 13360 19907 13412 19916
rect 13360 19873 13369 19907
rect 13369 19873 13403 19907
rect 13403 19873 13412 19907
rect 13360 19864 13412 19873
rect 14556 19796 14608 19848
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 16028 19864 16080 19916
rect 17132 19932 17184 19984
rect 16304 19907 16356 19916
rect 16304 19873 16311 19907
rect 16311 19873 16356 19907
rect 16304 19864 16356 19873
rect 16396 19907 16448 19916
rect 16396 19873 16405 19907
rect 16405 19873 16439 19907
rect 16439 19873 16448 19907
rect 16396 19864 16448 19873
rect 16672 19864 16724 19916
rect 16948 19864 17000 19916
rect 17592 19975 17644 19984
rect 17592 19941 17601 19975
rect 17601 19941 17635 19975
rect 17635 19941 17644 19975
rect 17592 19932 17644 19941
rect 19432 20000 19484 20052
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 18512 19864 18564 19916
rect 18696 19864 18748 19916
rect 16580 19728 16632 19780
rect 17592 19728 17644 19780
rect 9772 19660 9824 19712
rect 15292 19660 15344 19712
rect 15476 19660 15528 19712
rect 16396 19660 16448 19712
rect 16488 19660 16540 19712
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 19616 19907 19668 19916
rect 19616 19873 19625 19907
rect 19625 19873 19659 19907
rect 19659 19873 19668 19907
rect 19616 19864 19668 19873
rect 19064 19728 19116 19780
rect 20352 20000 20404 20052
rect 22192 20000 22244 20052
rect 26424 20000 26476 20052
rect 22836 19932 22888 19984
rect 20904 19864 20956 19916
rect 21548 19907 21600 19916
rect 21548 19873 21557 19907
rect 21557 19873 21591 19907
rect 21591 19873 21600 19907
rect 21548 19864 21600 19873
rect 22192 19864 22244 19916
rect 22284 19728 22336 19780
rect 23112 19907 23164 19916
rect 23112 19873 23121 19907
rect 23121 19873 23155 19907
rect 23155 19873 23164 19907
rect 23112 19864 23164 19873
rect 23204 19907 23256 19916
rect 23204 19873 23213 19907
rect 23213 19873 23247 19907
rect 23247 19873 23256 19907
rect 23204 19864 23256 19873
rect 24216 19932 24268 19984
rect 27528 19932 27580 19984
rect 29184 20000 29236 20052
rect 29460 20043 29512 20052
rect 29460 20009 29469 20043
rect 29469 20009 29503 20043
rect 29503 20009 29512 20043
rect 29460 20000 29512 20009
rect 23480 19907 23532 19916
rect 23480 19873 23489 19907
rect 23489 19873 23523 19907
rect 23523 19873 23532 19907
rect 23480 19864 23532 19873
rect 23756 19907 23808 19916
rect 23756 19873 23765 19907
rect 23765 19873 23799 19907
rect 23799 19873 23808 19907
rect 23756 19864 23808 19873
rect 22744 19796 22796 19848
rect 22836 19796 22888 19848
rect 24124 19907 24176 19916
rect 24124 19873 24133 19907
rect 24133 19873 24167 19907
rect 24167 19873 24176 19907
rect 24124 19864 24176 19873
rect 25780 19864 25832 19916
rect 27988 19864 28040 19916
rect 28816 19907 28868 19916
rect 28816 19873 28825 19907
rect 28825 19873 28859 19907
rect 28859 19873 28868 19907
rect 28816 19864 28868 19873
rect 29644 19932 29696 19984
rect 25596 19796 25648 19848
rect 25872 19728 25924 19780
rect 21272 19660 21324 19712
rect 22744 19660 22796 19712
rect 23020 19660 23072 19712
rect 25136 19703 25188 19712
rect 25136 19669 25145 19703
rect 25145 19669 25179 19703
rect 25179 19669 25188 19703
rect 25136 19660 25188 19669
rect 27436 19660 27488 19712
rect 27988 19703 28040 19712
rect 27988 19669 27997 19703
rect 27997 19669 28031 19703
rect 28031 19669 28040 19703
rect 27988 19660 28040 19669
rect 29552 19907 29604 19916
rect 29552 19873 29561 19907
rect 29561 19873 29595 19907
rect 29595 19873 29604 19907
rect 29552 19864 29604 19873
rect 29828 19907 29880 19916
rect 29828 19873 29862 19907
rect 29862 19873 29880 19907
rect 29828 19864 29880 19873
rect 29368 19796 29420 19848
rect 29736 19660 29788 19712
rect 29920 19660 29972 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 11436 19558 11488 19610
rect 11500 19558 11552 19610
rect 11564 19558 11616 19610
rect 11628 19558 11680 19610
rect 11692 19558 11744 19610
rect 19210 19558 19262 19610
rect 19274 19558 19326 19610
rect 19338 19558 19390 19610
rect 19402 19558 19454 19610
rect 19466 19558 19518 19610
rect 26984 19558 27036 19610
rect 27048 19558 27100 19610
rect 27112 19558 27164 19610
rect 27176 19558 27228 19610
rect 27240 19558 27292 19610
rect 2412 19499 2464 19508
rect 2412 19465 2421 19499
rect 2421 19465 2455 19499
rect 2455 19465 2464 19499
rect 2412 19456 2464 19465
rect 6276 19456 6328 19508
rect 6460 19499 6512 19508
rect 6460 19465 6469 19499
rect 6469 19465 6503 19499
rect 6503 19465 6512 19499
rect 6460 19456 6512 19465
rect 9772 19456 9824 19508
rect 15660 19456 15712 19508
rect 16764 19499 16816 19508
rect 16764 19465 16773 19499
rect 16773 19465 16807 19499
rect 16807 19465 16816 19499
rect 16764 19456 16816 19465
rect 3240 19388 3292 19440
rect 3148 19320 3200 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2136 19295 2188 19304
rect 2136 19261 2145 19295
rect 2145 19261 2179 19295
rect 2179 19261 2188 19295
rect 2136 19252 2188 19261
rect 2412 19252 2464 19304
rect 2504 19252 2556 19304
rect 2596 19184 2648 19236
rect 3056 19295 3108 19304
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 3332 19252 3384 19304
rect 4252 19320 4304 19372
rect 4896 19320 4948 19372
rect 3608 19227 3660 19236
rect 3608 19193 3617 19227
rect 3617 19193 3651 19227
rect 3651 19193 3660 19227
rect 3608 19184 3660 19193
rect 4068 19252 4120 19304
rect 15568 19388 15620 19440
rect 16488 19388 16540 19440
rect 17224 19456 17276 19508
rect 5816 19295 5868 19304
rect 5816 19261 5825 19295
rect 5825 19261 5859 19295
rect 5859 19261 5868 19295
rect 5816 19252 5868 19261
rect 6368 19252 6420 19304
rect 6460 19252 6512 19304
rect 16120 19320 16172 19372
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 18052 19456 18104 19508
rect 18236 19456 18288 19508
rect 21180 19456 21232 19508
rect 22836 19456 22888 19508
rect 23204 19456 23256 19508
rect 28080 19456 28132 19508
rect 29828 19456 29880 19508
rect 20260 19388 20312 19440
rect 20536 19388 20588 19440
rect 6920 19252 6972 19304
rect 8208 19252 8260 19304
rect 10232 19252 10284 19304
rect 11060 19252 11112 19304
rect 14556 19295 14608 19304
rect 14556 19261 14565 19295
rect 14565 19261 14599 19295
rect 14599 19261 14608 19295
rect 14556 19252 14608 19261
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 14832 19252 14884 19304
rect 3516 19116 3568 19168
rect 4712 19184 4764 19236
rect 5080 19184 5132 19236
rect 6184 19227 6236 19236
rect 6184 19193 6193 19227
rect 6193 19193 6227 19227
rect 6227 19193 6236 19227
rect 6184 19184 6236 19193
rect 6644 19227 6696 19236
rect 6644 19193 6653 19227
rect 6653 19193 6687 19227
rect 6687 19193 6696 19227
rect 6644 19184 6696 19193
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 15752 19295 15804 19304
rect 15752 19261 15761 19295
rect 15761 19261 15795 19295
rect 15795 19261 15804 19295
rect 15752 19252 15804 19261
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 16764 19252 16816 19304
rect 16856 19295 16908 19304
rect 16856 19261 16865 19295
rect 16865 19261 16899 19295
rect 16899 19261 16908 19295
rect 16856 19252 16908 19261
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 16396 19184 16448 19236
rect 16948 19184 17000 19236
rect 17040 19184 17092 19236
rect 17592 19252 17644 19304
rect 17868 19295 17920 19304
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 19708 19320 19760 19372
rect 21088 19320 21140 19372
rect 22376 19320 22428 19372
rect 18972 19252 19024 19261
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 19616 19252 19668 19304
rect 21824 19295 21876 19304
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 22652 19252 22704 19304
rect 22744 19295 22796 19304
rect 22744 19261 22753 19295
rect 22753 19261 22787 19295
rect 22787 19261 22796 19295
rect 22744 19252 22796 19261
rect 23020 19252 23072 19304
rect 25780 19320 25832 19372
rect 25872 19363 25924 19372
rect 25872 19329 25881 19363
rect 25881 19329 25915 19363
rect 25915 19329 25924 19363
rect 25872 19320 25924 19329
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 25504 19295 25556 19304
rect 25504 19261 25522 19295
rect 25522 19261 25556 19295
rect 25504 19252 25556 19261
rect 25596 19295 25648 19304
rect 25596 19261 25605 19295
rect 25605 19261 25639 19295
rect 25639 19261 25648 19295
rect 25596 19252 25648 19261
rect 19800 19184 19852 19236
rect 4160 19116 4212 19168
rect 6276 19116 6328 19168
rect 11428 19116 11480 19168
rect 15752 19116 15804 19168
rect 20996 19159 21048 19168
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 22376 19184 22428 19236
rect 21364 19159 21416 19168
rect 21364 19125 21373 19159
rect 21373 19125 21407 19159
rect 21407 19125 21416 19159
rect 26700 19295 26752 19304
rect 26700 19261 26709 19295
rect 26709 19261 26743 19295
rect 26743 19261 26752 19295
rect 26700 19252 26752 19261
rect 26884 19295 26936 19304
rect 26884 19261 26893 19295
rect 26893 19261 26927 19295
rect 26927 19261 26936 19295
rect 26884 19252 26936 19261
rect 26976 19295 27028 19304
rect 26976 19261 26985 19295
rect 26985 19261 27019 19295
rect 27019 19261 27028 19295
rect 26976 19252 27028 19261
rect 26792 19184 26844 19236
rect 21364 19116 21416 19125
rect 23020 19159 23072 19168
rect 23020 19125 23029 19159
rect 23029 19125 23063 19159
rect 23063 19125 23072 19159
rect 23020 19116 23072 19125
rect 24584 19116 24636 19168
rect 24676 19159 24728 19168
rect 24676 19125 24685 19159
rect 24685 19125 24719 19159
rect 24719 19125 24728 19159
rect 24676 19116 24728 19125
rect 25044 19116 25096 19168
rect 25504 19116 25556 19168
rect 27436 19295 27488 19304
rect 27436 19261 27445 19295
rect 27445 19261 27479 19295
rect 27479 19261 27488 19295
rect 27436 19252 27488 19261
rect 29460 19388 29512 19440
rect 29920 19388 29972 19440
rect 28816 19320 28868 19372
rect 29092 19295 29144 19304
rect 29092 19261 29101 19295
rect 29101 19261 29135 19295
rect 29135 19261 29144 19295
rect 29092 19252 29144 19261
rect 29368 19295 29420 19304
rect 29368 19261 29377 19295
rect 29377 19261 29411 19295
rect 29411 19261 29420 19295
rect 29368 19252 29420 19261
rect 29460 19295 29512 19304
rect 29460 19261 29469 19295
rect 29469 19261 29503 19295
rect 29503 19261 29512 19295
rect 29460 19252 29512 19261
rect 29828 19252 29880 19304
rect 30196 19252 30248 19304
rect 30288 19295 30340 19304
rect 30288 19261 30297 19295
rect 30297 19261 30331 19295
rect 30331 19261 30340 19295
rect 30288 19252 30340 19261
rect 30380 19295 30432 19304
rect 30380 19261 30389 19295
rect 30389 19261 30423 19295
rect 30423 19261 30432 19295
rect 30380 19252 30432 19261
rect 29920 19184 29972 19236
rect 29368 19116 29420 19168
rect 29736 19116 29788 19168
rect 30656 19159 30708 19168
rect 30656 19125 30665 19159
rect 30665 19125 30699 19159
rect 30699 19125 30708 19159
rect 30656 19116 30708 19125
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 12096 19014 12148 19066
rect 12160 19014 12212 19066
rect 12224 19014 12276 19066
rect 12288 19014 12340 19066
rect 12352 19014 12404 19066
rect 19870 19014 19922 19066
rect 19934 19014 19986 19066
rect 19998 19014 20050 19066
rect 20062 19014 20114 19066
rect 20126 19014 20178 19066
rect 27644 19014 27696 19066
rect 27708 19014 27760 19066
rect 27772 19014 27824 19066
rect 27836 19014 27888 19066
rect 27900 19014 27952 19066
rect 2136 18912 2188 18964
rect 5080 18955 5132 18964
rect 5080 18921 5089 18955
rect 5089 18921 5123 18955
rect 5123 18921 5132 18955
rect 5080 18912 5132 18921
rect 5172 18912 5224 18964
rect 6184 18912 6236 18964
rect 6552 18912 6604 18964
rect 7196 18955 7248 18964
rect 7196 18921 7205 18955
rect 7205 18921 7239 18955
rect 7239 18921 7248 18955
rect 7196 18912 7248 18921
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 13820 18912 13872 18964
rect 16488 18955 16540 18964
rect 16488 18921 16497 18955
rect 16497 18921 16531 18955
rect 16531 18921 16540 18955
rect 16488 18912 16540 18921
rect 17316 18912 17368 18964
rect 17592 18912 17644 18964
rect 17776 18912 17828 18964
rect 2964 18844 3016 18896
rect 5816 18844 5868 18896
rect 6092 18844 6144 18896
rect 2412 18819 2464 18828
rect 2412 18785 2421 18819
rect 2421 18785 2455 18819
rect 2455 18785 2464 18819
rect 2412 18776 2464 18785
rect 2596 18819 2648 18828
rect 2596 18785 2605 18819
rect 2605 18785 2639 18819
rect 2639 18785 2648 18819
rect 2596 18776 2648 18785
rect 2688 18819 2740 18828
rect 2688 18785 2697 18819
rect 2697 18785 2731 18819
rect 2731 18785 2740 18819
rect 2688 18776 2740 18785
rect 3424 18776 3476 18828
rect 2044 18708 2096 18760
rect 3608 18708 3660 18760
rect 2136 18572 2188 18624
rect 3516 18640 3568 18692
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 5172 18819 5224 18828
rect 5172 18785 5181 18819
rect 5181 18785 5215 18819
rect 5215 18785 5224 18819
rect 5172 18776 5224 18785
rect 6184 18819 6236 18828
rect 6184 18785 6193 18819
rect 6193 18785 6227 18819
rect 6227 18785 6236 18819
rect 6184 18776 6236 18785
rect 11428 18887 11480 18896
rect 11428 18853 11437 18887
rect 11437 18853 11471 18887
rect 11471 18853 11480 18887
rect 11428 18844 11480 18853
rect 6920 18776 6972 18828
rect 8116 18776 8168 18828
rect 11060 18776 11112 18828
rect 11796 18776 11848 18828
rect 15200 18844 15252 18896
rect 9404 18708 9456 18760
rect 10968 18708 11020 18760
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 15292 18776 15344 18828
rect 11336 18640 11388 18692
rect 15568 18776 15620 18828
rect 15752 18819 15804 18828
rect 15752 18785 15761 18819
rect 15761 18785 15795 18819
rect 15795 18785 15804 18819
rect 15752 18776 15804 18785
rect 16120 18819 16172 18828
rect 16120 18785 16129 18819
rect 16129 18785 16163 18819
rect 16163 18785 16172 18819
rect 16120 18776 16172 18785
rect 19708 18844 19760 18896
rect 16212 18708 16264 18760
rect 15844 18640 15896 18692
rect 16948 18819 17000 18828
rect 16948 18785 16957 18819
rect 16957 18785 16991 18819
rect 16991 18785 17000 18819
rect 16948 18776 17000 18785
rect 17040 18776 17092 18828
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 17684 18776 17736 18828
rect 18052 18776 18104 18828
rect 18788 18776 18840 18828
rect 20260 18819 20312 18828
rect 20260 18785 20269 18819
rect 20269 18785 20303 18819
rect 20303 18785 20312 18819
rect 20260 18776 20312 18785
rect 20904 18912 20956 18964
rect 22284 18912 22336 18964
rect 22376 18912 22428 18964
rect 21548 18887 21600 18896
rect 21548 18853 21582 18887
rect 21582 18853 21600 18887
rect 21548 18844 21600 18853
rect 21824 18844 21876 18896
rect 20536 18776 20588 18828
rect 20628 18819 20680 18828
rect 20628 18785 20637 18819
rect 20637 18785 20671 18819
rect 20671 18785 20680 18819
rect 20628 18776 20680 18785
rect 20720 18819 20772 18828
rect 20720 18785 20729 18819
rect 20729 18785 20763 18819
rect 20763 18785 20772 18819
rect 20720 18776 20772 18785
rect 17500 18708 17552 18760
rect 18972 18708 19024 18760
rect 19616 18708 19668 18760
rect 20996 18776 21048 18828
rect 21272 18819 21324 18828
rect 21272 18785 21281 18819
rect 21281 18785 21315 18819
rect 21315 18785 21324 18819
rect 21272 18776 21324 18785
rect 22928 18819 22980 18828
rect 22928 18785 22937 18819
rect 22937 18785 22971 18819
rect 22971 18785 22980 18819
rect 22928 18776 22980 18785
rect 24032 18819 24084 18828
rect 24032 18785 24041 18819
rect 24041 18785 24075 18819
rect 24075 18785 24084 18819
rect 24032 18776 24084 18785
rect 24124 18819 24176 18828
rect 24124 18785 24133 18819
rect 24133 18785 24167 18819
rect 24167 18785 24176 18819
rect 24124 18776 24176 18785
rect 25136 18912 25188 18964
rect 25596 18912 25648 18964
rect 26056 18912 26108 18964
rect 26884 18912 26936 18964
rect 27436 18912 27488 18964
rect 27988 18844 28040 18896
rect 24584 18819 24636 18828
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 26700 18776 26752 18828
rect 26792 18819 26844 18828
rect 26792 18785 26801 18819
rect 26801 18785 26835 18819
rect 26835 18785 26844 18819
rect 26792 18776 26844 18785
rect 17316 18640 17368 18692
rect 17684 18640 17736 18692
rect 20904 18640 20956 18692
rect 27528 18819 27580 18828
rect 27528 18785 27537 18819
rect 27537 18785 27571 18819
rect 27571 18785 27580 18819
rect 27528 18776 27580 18785
rect 27712 18819 27764 18828
rect 27712 18785 27721 18819
rect 27721 18785 27755 18819
rect 27755 18785 27764 18819
rect 27712 18776 27764 18785
rect 27804 18819 27856 18828
rect 27804 18785 27813 18819
rect 27813 18785 27847 18819
rect 27847 18785 27856 18819
rect 27804 18776 27856 18785
rect 28080 18776 28132 18828
rect 29368 18955 29420 18964
rect 29368 18921 29377 18955
rect 29377 18921 29411 18955
rect 29411 18921 29420 18955
rect 29368 18912 29420 18921
rect 29460 18955 29512 18964
rect 29460 18921 29469 18955
rect 29469 18921 29503 18955
rect 29503 18921 29512 18955
rect 29460 18912 29512 18921
rect 29552 18912 29604 18964
rect 29736 18912 29788 18964
rect 29828 18955 29880 18964
rect 29828 18921 29837 18955
rect 29837 18921 29871 18955
rect 29871 18921 29880 18955
rect 29828 18912 29880 18921
rect 29920 18955 29972 18964
rect 29920 18921 29929 18955
rect 29929 18921 29963 18955
rect 29963 18921 29972 18955
rect 29920 18912 29972 18921
rect 30380 18912 30432 18964
rect 30288 18844 30340 18896
rect 28632 18819 28684 18828
rect 28632 18785 28641 18819
rect 28641 18785 28675 18819
rect 28675 18785 28684 18819
rect 28632 18776 28684 18785
rect 29460 18776 29512 18828
rect 30104 18819 30156 18828
rect 30104 18785 30113 18819
rect 30113 18785 30147 18819
rect 30147 18785 30156 18819
rect 30104 18776 30156 18785
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 29184 18751 29236 18760
rect 4344 18572 4396 18624
rect 7104 18572 7156 18624
rect 8208 18572 8260 18624
rect 15384 18572 15436 18624
rect 16028 18572 16080 18624
rect 16488 18572 16540 18624
rect 16672 18572 16724 18624
rect 17408 18572 17460 18624
rect 17868 18572 17920 18624
rect 20996 18572 21048 18624
rect 21548 18572 21600 18624
rect 22836 18615 22888 18624
rect 22836 18581 22845 18615
rect 22845 18581 22879 18615
rect 22879 18581 22888 18615
rect 22836 18572 22888 18581
rect 25504 18572 25556 18624
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 29552 18708 29604 18760
rect 29092 18640 29144 18692
rect 30472 18640 30524 18692
rect 30656 18640 30708 18692
rect 27804 18572 27856 18624
rect 28816 18572 28868 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 11436 18470 11488 18522
rect 11500 18470 11552 18522
rect 11564 18470 11616 18522
rect 11628 18470 11680 18522
rect 11692 18470 11744 18522
rect 19210 18470 19262 18522
rect 19274 18470 19326 18522
rect 19338 18470 19390 18522
rect 19402 18470 19454 18522
rect 19466 18470 19518 18522
rect 26984 18470 27036 18522
rect 27048 18470 27100 18522
rect 27112 18470 27164 18522
rect 27176 18470 27228 18522
rect 27240 18470 27292 18522
rect 2596 18368 2648 18420
rect 5908 18368 5960 18420
rect 10508 18368 10560 18420
rect 10968 18411 11020 18420
rect 10968 18377 10977 18411
rect 10977 18377 11011 18411
rect 11011 18377 11020 18411
rect 10968 18368 11020 18377
rect 15292 18411 15344 18420
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15292 18368 15344 18377
rect 6920 18343 6972 18352
rect 6920 18309 6929 18343
rect 6929 18309 6963 18343
rect 6963 18309 6972 18343
rect 6920 18300 6972 18309
rect 2228 18164 2280 18216
rect 2688 18164 2740 18216
rect 1308 18071 1360 18080
rect 1308 18037 1317 18071
rect 1317 18037 1351 18071
rect 1351 18037 1360 18071
rect 1308 18028 1360 18037
rect 1860 18139 1912 18148
rect 1860 18105 1869 18139
rect 1869 18105 1903 18139
rect 1903 18105 1912 18139
rect 1860 18096 1912 18105
rect 2044 18096 2096 18148
rect 2136 18139 2188 18148
rect 2136 18105 2145 18139
rect 2145 18105 2179 18139
rect 2179 18105 2188 18139
rect 2136 18096 2188 18105
rect 2872 18096 2924 18148
rect 6276 18164 6328 18216
rect 7656 18164 7708 18216
rect 7748 18207 7800 18216
rect 7748 18173 7757 18207
rect 7757 18173 7791 18207
rect 7791 18173 7800 18207
rect 7748 18164 7800 18173
rect 4252 18096 4304 18148
rect 4344 18139 4396 18148
rect 4344 18105 4362 18139
rect 4362 18105 4396 18139
rect 4344 18096 4396 18105
rect 6644 18096 6696 18148
rect 3792 18028 3844 18080
rect 4160 18028 4212 18080
rect 7380 18096 7432 18148
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 7564 18028 7616 18080
rect 8208 18164 8260 18216
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 9496 18096 9548 18148
rect 10508 18207 10560 18216
rect 10508 18173 10517 18207
rect 10517 18173 10551 18207
rect 10551 18173 10560 18207
rect 10508 18164 10560 18173
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 13636 18207 13688 18216
rect 12624 18164 12676 18173
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 14188 18207 14240 18216
rect 14188 18173 14197 18207
rect 14197 18173 14231 18207
rect 14231 18173 14240 18207
rect 14188 18164 14240 18173
rect 15844 18207 15896 18216
rect 15844 18173 15853 18207
rect 15853 18173 15887 18207
rect 15887 18173 15896 18207
rect 15844 18164 15896 18173
rect 17408 18368 17460 18420
rect 16856 18300 16908 18352
rect 17868 18368 17920 18420
rect 20260 18368 20312 18420
rect 20720 18368 20772 18420
rect 16396 18232 16448 18284
rect 16212 18207 16264 18216
rect 16212 18173 16221 18207
rect 16221 18173 16255 18207
rect 16255 18173 16264 18207
rect 16212 18164 16264 18173
rect 10876 18096 10928 18148
rect 11612 18096 11664 18148
rect 15200 18096 15252 18148
rect 10048 18028 10100 18080
rect 15292 18028 15344 18080
rect 16304 18096 16356 18148
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 17500 18275 17552 18284
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 18236 18232 18288 18284
rect 22192 18368 22244 18420
rect 22836 18368 22888 18420
rect 24032 18368 24084 18420
rect 27712 18368 27764 18420
rect 28080 18411 28132 18420
rect 28080 18377 28089 18411
rect 28089 18377 28123 18411
rect 28123 18377 28132 18411
rect 28080 18368 28132 18377
rect 29552 18368 29604 18420
rect 30104 18368 30156 18420
rect 23296 18300 23348 18352
rect 17132 18164 17184 18216
rect 15936 18028 15988 18080
rect 16488 18028 16540 18080
rect 17868 18096 17920 18148
rect 19800 18164 19852 18216
rect 20076 18207 20128 18216
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20444 18207 20496 18216
rect 20444 18173 20453 18207
rect 20453 18173 20487 18207
rect 20487 18173 20496 18207
rect 20444 18164 20496 18173
rect 20996 18275 21048 18284
rect 20996 18241 21005 18275
rect 21005 18241 21039 18275
rect 21039 18241 21048 18275
rect 20996 18232 21048 18241
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 21180 18275 21232 18284
rect 21180 18241 21189 18275
rect 21189 18241 21223 18275
rect 21223 18241 21232 18275
rect 21180 18232 21232 18241
rect 18880 18096 18932 18148
rect 21364 18164 21416 18216
rect 23020 18164 23072 18216
rect 23296 18139 23348 18148
rect 23296 18105 23305 18139
rect 23305 18105 23339 18139
rect 23339 18105 23348 18139
rect 23296 18096 23348 18105
rect 24492 18164 24544 18216
rect 25228 18232 25280 18284
rect 25044 18164 25096 18216
rect 25136 18164 25188 18216
rect 27620 18300 27672 18352
rect 28356 18300 28408 18352
rect 29092 18300 29144 18352
rect 29184 18300 29236 18352
rect 26056 18207 26108 18216
rect 26056 18173 26065 18207
rect 26065 18173 26099 18207
rect 26099 18173 26108 18207
rect 26056 18164 26108 18173
rect 19616 18028 19668 18080
rect 20904 18028 20956 18080
rect 24584 18028 24636 18080
rect 24952 18028 25004 18080
rect 25320 18028 25372 18080
rect 26148 18096 26200 18148
rect 26608 18207 26660 18216
rect 26608 18173 26617 18207
rect 26617 18173 26651 18207
rect 26651 18173 26660 18207
rect 26608 18164 26660 18173
rect 26792 18164 26844 18216
rect 27436 18096 27488 18148
rect 27620 18096 27672 18148
rect 29552 18275 29604 18284
rect 29552 18241 29561 18275
rect 29561 18241 29595 18275
rect 29595 18241 29604 18275
rect 29552 18232 29604 18241
rect 29644 18232 29696 18284
rect 28356 18207 28408 18216
rect 28356 18173 28365 18207
rect 28365 18173 28399 18207
rect 28399 18173 28408 18207
rect 28356 18164 28408 18173
rect 29460 18164 29512 18216
rect 28632 18096 28684 18148
rect 28908 18096 28960 18148
rect 29644 18096 29696 18148
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 12096 17926 12148 17978
rect 12160 17926 12212 17978
rect 12224 17926 12276 17978
rect 12288 17926 12340 17978
rect 12352 17926 12404 17978
rect 19870 17926 19922 17978
rect 19934 17926 19986 17978
rect 19998 17926 20050 17978
rect 20062 17926 20114 17978
rect 20126 17926 20178 17978
rect 27644 17926 27696 17978
rect 27708 17926 27760 17978
rect 27772 17926 27824 17978
rect 27836 17926 27888 17978
rect 27900 17926 27952 17978
rect 3516 17824 3568 17876
rect 4252 17867 4304 17876
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 2688 17756 2740 17808
rect 1308 17688 1360 17740
rect 2228 17731 2280 17740
rect 2228 17697 2262 17731
rect 2262 17697 2280 17731
rect 2228 17688 2280 17697
rect 3516 17688 3568 17740
rect 3792 17731 3844 17740
rect 3792 17697 3801 17731
rect 3801 17697 3835 17731
rect 3835 17697 3844 17731
rect 3792 17688 3844 17697
rect 5816 17799 5868 17808
rect 5816 17765 5825 17799
rect 5825 17765 5859 17799
rect 5859 17765 5868 17799
rect 5816 17756 5868 17765
rect 4252 17688 4304 17740
rect 5172 17688 5224 17740
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 4436 17620 4488 17672
rect 6644 17731 6696 17740
rect 6644 17697 6653 17731
rect 6653 17697 6687 17731
rect 6687 17697 6696 17731
rect 6644 17688 6696 17697
rect 7840 17824 7892 17876
rect 9496 17867 9548 17876
rect 9496 17833 9505 17867
rect 9505 17833 9539 17867
rect 9539 17833 9548 17867
rect 9496 17824 9548 17833
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10140 17824 10192 17833
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 11612 17867 11664 17876
rect 11612 17833 11621 17867
rect 11621 17833 11655 17867
rect 11655 17833 11664 17867
rect 11612 17824 11664 17833
rect 13268 17867 13320 17876
rect 13268 17833 13277 17867
rect 13277 17833 13311 17867
rect 13311 17833 13320 17867
rect 13268 17824 13320 17833
rect 14188 17824 14240 17876
rect 15752 17824 15804 17876
rect 16304 17824 16356 17876
rect 17868 17824 17920 17876
rect 25228 17867 25280 17876
rect 25228 17833 25237 17867
rect 25237 17833 25271 17867
rect 25271 17833 25280 17867
rect 25228 17824 25280 17833
rect 28172 17824 28224 17876
rect 29000 17824 29052 17876
rect 29276 17824 29328 17876
rect 29368 17867 29420 17876
rect 29368 17833 29377 17867
rect 29377 17833 29411 17867
rect 29411 17833 29420 17867
rect 29368 17824 29420 17833
rect 7380 17756 7432 17808
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 7564 17731 7616 17740
rect 7564 17697 7598 17731
rect 7598 17697 7616 17731
rect 7564 17688 7616 17697
rect 6920 17620 6972 17672
rect 9496 17620 9548 17672
rect 10876 17756 10928 17808
rect 10508 17731 10560 17740
rect 10508 17697 10517 17731
rect 10517 17697 10551 17731
rect 10551 17697 10560 17731
rect 10508 17688 10560 17697
rect 4712 17552 4764 17604
rect 3976 17484 4028 17536
rect 4160 17484 4212 17536
rect 6092 17527 6144 17536
rect 6092 17493 6101 17527
rect 6101 17493 6135 17527
rect 6135 17493 6144 17527
rect 6092 17484 6144 17493
rect 8392 17484 8444 17536
rect 8668 17527 8720 17536
rect 8668 17493 8677 17527
rect 8677 17493 8711 17527
rect 8711 17493 8720 17527
rect 8668 17484 8720 17493
rect 9680 17484 9732 17536
rect 10416 17484 10468 17536
rect 11060 17620 11112 17672
rect 11336 17731 11388 17740
rect 11336 17697 11345 17731
rect 11345 17697 11379 17731
rect 11379 17697 11388 17731
rect 11336 17688 11388 17697
rect 13636 17756 13688 17808
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 11152 17552 11204 17604
rect 12808 17663 12860 17672
rect 12808 17629 12817 17663
rect 12817 17629 12851 17663
rect 12851 17629 12860 17663
rect 13820 17731 13872 17740
rect 13820 17697 13829 17731
rect 13829 17697 13863 17731
rect 13863 17697 13872 17731
rect 13820 17688 13872 17697
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 12808 17620 12860 17629
rect 14832 17620 14884 17672
rect 15200 17688 15252 17740
rect 15384 17688 15436 17740
rect 16396 17731 16448 17740
rect 16396 17697 16405 17731
rect 16405 17697 16439 17731
rect 16439 17697 16448 17731
rect 16396 17688 16448 17697
rect 16672 17756 16724 17808
rect 16580 17731 16632 17740
rect 16580 17697 16589 17731
rect 16589 17697 16623 17731
rect 16623 17697 16632 17731
rect 16580 17688 16632 17697
rect 16764 17731 16816 17740
rect 16764 17697 16773 17731
rect 16773 17697 16807 17731
rect 16807 17697 16816 17731
rect 16764 17688 16816 17697
rect 17316 17688 17368 17740
rect 20536 17731 20588 17740
rect 20536 17697 20545 17731
rect 20545 17697 20579 17731
rect 20579 17697 20588 17731
rect 20536 17688 20588 17697
rect 20628 17731 20680 17740
rect 20628 17697 20637 17731
rect 20637 17697 20671 17731
rect 20671 17697 20680 17731
rect 20628 17688 20680 17697
rect 16212 17620 16264 17672
rect 16856 17620 16908 17672
rect 17592 17620 17644 17672
rect 20904 17731 20956 17740
rect 20904 17697 20913 17731
rect 20913 17697 20947 17731
rect 20947 17697 20956 17731
rect 20904 17688 20956 17697
rect 21916 17731 21968 17740
rect 21916 17697 21925 17731
rect 21925 17697 21959 17731
rect 21959 17697 21968 17731
rect 21916 17688 21968 17697
rect 22192 17731 22244 17740
rect 22192 17697 22201 17731
rect 22201 17697 22235 17731
rect 22235 17697 22244 17731
rect 22192 17688 22244 17697
rect 23296 17688 23348 17740
rect 12532 17484 12584 17536
rect 15568 17552 15620 17604
rect 16488 17552 16540 17604
rect 16764 17552 16816 17604
rect 21548 17620 21600 17672
rect 21272 17595 21324 17604
rect 21272 17561 21281 17595
rect 21281 17561 21315 17595
rect 21315 17561 21324 17595
rect 21272 17552 21324 17561
rect 21456 17552 21508 17604
rect 22468 17595 22520 17604
rect 22468 17561 22477 17595
rect 22477 17561 22511 17595
rect 22511 17561 22520 17595
rect 22468 17552 22520 17561
rect 23020 17620 23072 17672
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 23480 17688 23532 17740
rect 24216 17688 24268 17740
rect 24584 17731 24636 17740
rect 24584 17697 24593 17731
rect 24593 17697 24627 17731
rect 24627 17697 24636 17731
rect 24584 17688 24636 17697
rect 24768 17731 24820 17740
rect 24768 17697 24777 17731
rect 24777 17697 24811 17731
rect 24811 17697 24820 17731
rect 24768 17688 24820 17697
rect 26332 17756 26384 17808
rect 26608 17756 26660 17808
rect 24952 17731 25004 17740
rect 24952 17697 24961 17731
rect 24961 17697 24995 17731
rect 24995 17697 25004 17731
rect 24952 17688 25004 17697
rect 28540 17756 28592 17808
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 15660 17484 15712 17493
rect 20444 17484 20496 17536
rect 22376 17484 22428 17536
rect 23388 17484 23440 17536
rect 27528 17620 27580 17672
rect 28632 17620 28684 17672
rect 24860 17552 24912 17604
rect 28356 17552 28408 17604
rect 29552 17688 29604 17740
rect 29644 17620 29696 17672
rect 29552 17552 29604 17604
rect 23572 17527 23624 17536
rect 23572 17493 23581 17527
rect 23581 17493 23615 17527
rect 23615 17493 23624 17527
rect 23572 17484 23624 17493
rect 23664 17484 23716 17536
rect 24768 17484 24820 17536
rect 26240 17484 26292 17536
rect 27988 17484 28040 17536
rect 29000 17484 29052 17536
rect 30656 17484 30708 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 11436 17382 11488 17434
rect 11500 17382 11552 17434
rect 11564 17382 11616 17434
rect 11628 17382 11680 17434
rect 11692 17382 11744 17434
rect 19210 17382 19262 17434
rect 19274 17382 19326 17434
rect 19338 17382 19390 17434
rect 19402 17382 19454 17434
rect 19466 17382 19518 17434
rect 26984 17382 27036 17434
rect 27048 17382 27100 17434
rect 27112 17382 27164 17434
rect 27176 17382 27228 17434
rect 27240 17382 27292 17434
rect 2228 17280 2280 17332
rect 2964 17280 3016 17332
rect 6644 17280 6696 17332
rect 6920 17280 6972 17332
rect 7748 17280 7800 17332
rect 3056 17212 3108 17264
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 2872 17119 2924 17128
rect 2872 17085 2881 17119
rect 2881 17085 2915 17119
rect 2915 17085 2924 17119
rect 2872 17076 2924 17085
rect 6828 17212 6880 17264
rect 3148 17076 3200 17128
rect 3240 17051 3292 17060
rect 3240 17017 3249 17051
rect 3249 17017 3283 17051
rect 3283 17017 3292 17051
rect 3240 17008 3292 17017
rect 3332 17008 3384 17060
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 4436 17144 4488 17196
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 8668 17280 8720 17332
rect 10140 17280 10192 17332
rect 10508 17280 10560 17332
rect 11336 17280 11388 17332
rect 11980 17280 12032 17332
rect 12624 17280 12676 17332
rect 8208 17076 8260 17128
rect 8576 17076 8628 17128
rect 9588 17076 9640 17128
rect 10968 17212 11020 17264
rect 11796 17144 11848 17196
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 11060 17076 11112 17128
rect 12532 17119 12584 17128
rect 12532 17085 12541 17119
rect 12541 17085 12575 17119
rect 12575 17085 12584 17119
rect 12532 17076 12584 17085
rect 12624 17119 12676 17128
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 13176 17144 13228 17196
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 13636 17144 13688 17153
rect 15292 17212 15344 17264
rect 16672 17280 16724 17332
rect 16948 17280 17000 17332
rect 18052 17212 18104 17264
rect 19248 17212 19300 17264
rect 19800 17212 19852 17264
rect 20444 17212 20496 17264
rect 20536 17212 20588 17264
rect 21548 17212 21600 17264
rect 15108 17119 15160 17128
rect 15108 17085 15117 17119
rect 15117 17085 15151 17119
rect 15151 17085 15160 17119
rect 15108 17076 15160 17085
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 15660 17144 15712 17196
rect 17408 17144 17460 17196
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 16948 17076 17000 17128
rect 19800 17076 19852 17128
rect 7380 17051 7432 17060
rect 7380 17017 7389 17051
rect 7389 17017 7423 17051
rect 7423 17017 7432 17051
rect 7380 17008 7432 17017
rect 3424 16940 3476 16992
rect 7656 16983 7708 16992
rect 7656 16949 7683 16983
rect 7683 16949 7708 16983
rect 7656 16940 7708 16949
rect 7840 17051 7892 17060
rect 7840 17017 7849 17051
rect 7849 17017 7883 17051
rect 7883 17017 7892 17051
rect 7840 17008 7892 17017
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 21640 17144 21692 17196
rect 22652 17187 22704 17196
rect 22652 17153 22661 17187
rect 22661 17153 22695 17187
rect 22695 17153 22704 17187
rect 22652 17144 22704 17153
rect 24124 17280 24176 17332
rect 24400 17280 24452 17332
rect 25136 17280 25188 17332
rect 27436 17280 27488 17332
rect 28172 17280 28224 17332
rect 28540 17280 28592 17332
rect 23112 17212 23164 17264
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 12532 16940 12584 16992
rect 12992 16940 13044 16992
rect 15476 16940 15528 16992
rect 16580 16940 16632 16992
rect 17224 16983 17276 16992
rect 17224 16949 17233 16983
rect 17233 16949 17267 16983
rect 17267 16949 17276 16983
rect 17224 16940 17276 16949
rect 17592 16983 17644 16992
rect 17592 16949 17601 16983
rect 17601 16949 17635 16983
rect 17635 16949 17644 16983
rect 17592 16940 17644 16949
rect 19616 16940 19668 16992
rect 21824 17076 21876 17128
rect 22928 17119 22980 17128
rect 22928 17085 22937 17119
rect 22937 17085 22971 17119
rect 22971 17085 22980 17119
rect 22928 17076 22980 17085
rect 23204 17144 23256 17196
rect 24400 17187 24452 17196
rect 24400 17153 24409 17187
rect 24409 17153 24443 17187
rect 24443 17153 24452 17187
rect 24400 17144 24452 17153
rect 23480 17076 23532 17128
rect 24860 17076 24912 17128
rect 27620 17212 27672 17264
rect 28264 17212 28316 17264
rect 28908 17212 28960 17264
rect 29460 17280 29512 17332
rect 30748 17280 30800 17332
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 25596 17144 25648 17196
rect 21732 16940 21784 16992
rect 24584 17008 24636 17060
rect 26240 17119 26292 17128
rect 26240 17085 26249 17119
rect 26249 17085 26283 17119
rect 26283 17085 26292 17119
rect 26240 17076 26292 17085
rect 26332 17119 26384 17128
rect 26332 17085 26341 17119
rect 26341 17085 26375 17119
rect 26375 17085 26384 17119
rect 26332 17076 26384 17085
rect 29368 17144 29420 17196
rect 30656 17187 30708 17196
rect 30656 17153 30665 17187
rect 30665 17153 30699 17187
rect 30699 17153 30708 17187
rect 30656 17144 30708 17153
rect 28172 17119 28224 17128
rect 28172 17085 28181 17119
rect 28181 17085 28215 17119
rect 28215 17085 28224 17119
rect 28172 17076 28224 17085
rect 28356 17119 28408 17128
rect 28356 17085 28365 17119
rect 28365 17085 28399 17119
rect 28399 17085 28408 17119
rect 28356 17076 28408 17085
rect 25504 17051 25556 17060
rect 25504 17017 25513 17051
rect 25513 17017 25547 17051
rect 25547 17017 25556 17051
rect 25504 17008 25556 17017
rect 25596 17051 25648 17060
rect 25596 17017 25605 17051
rect 25605 17017 25639 17051
rect 25639 17017 25648 17051
rect 25596 17008 25648 17017
rect 25872 17008 25924 17060
rect 27620 17008 27672 17060
rect 29000 17076 29052 17128
rect 31024 17076 31076 17128
rect 22560 16940 22612 16992
rect 22652 16940 22704 16992
rect 23204 16940 23256 16992
rect 23480 16940 23532 16992
rect 23940 16940 23992 16992
rect 25228 16940 25280 16992
rect 26056 16940 26108 16992
rect 26884 16940 26936 16992
rect 28172 16940 28224 16992
rect 29092 16983 29144 16992
rect 29092 16949 29101 16983
rect 29101 16949 29135 16983
rect 29135 16949 29144 16983
rect 29092 16940 29144 16949
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 12096 16838 12148 16890
rect 12160 16838 12212 16890
rect 12224 16838 12276 16890
rect 12288 16838 12340 16890
rect 12352 16838 12404 16890
rect 19870 16838 19922 16890
rect 19934 16838 19986 16890
rect 19998 16838 20050 16890
rect 20062 16838 20114 16890
rect 20126 16838 20178 16890
rect 27644 16838 27696 16890
rect 27708 16838 27760 16890
rect 27772 16838 27824 16890
rect 27836 16838 27888 16890
rect 27900 16838 27952 16890
rect 3148 16736 3200 16788
rect 6184 16736 6236 16788
rect 7656 16736 7708 16788
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 15200 16736 15252 16788
rect 1860 16711 1912 16720
rect 1860 16677 1869 16711
rect 1869 16677 1903 16711
rect 1903 16677 1912 16711
rect 1860 16668 1912 16677
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 7380 16668 7432 16720
rect 9956 16668 10008 16720
rect 10048 16668 10100 16720
rect 3056 16643 3108 16652
rect 3056 16609 3065 16643
rect 3065 16609 3099 16643
rect 3099 16609 3108 16643
rect 3056 16600 3108 16609
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 6184 16600 6236 16652
rect 7840 16600 7892 16652
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 8484 16643 8536 16652
rect 8484 16609 8493 16643
rect 8493 16609 8527 16643
rect 8527 16609 8536 16643
rect 8484 16600 8536 16609
rect 9036 16600 9088 16652
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 10324 16600 10376 16652
rect 10692 16600 10744 16652
rect 14648 16668 14700 16720
rect 15108 16668 15160 16720
rect 16304 16736 16356 16788
rect 17224 16736 17276 16788
rect 17408 16779 17460 16788
rect 17408 16745 17417 16779
rect 17417 16745 17451 16779
rect 17451 16745 17460 16779
rect 17408 16736 17460 16745
rect 17592 16736 17644 16788
rect 12992 16600 13044 16652
rect 2412 16532 2464 16584
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 3332 16532 3384 16584
rect 4068 16575 4120 16584
rect 4068 16541 4102 16575
rect 4102 16541 4120 16575
rect 4068 16532 4120 16541
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 7748 16464 7800 16516
rect 8392 16532 8444 16584
rect 10048 16532 10100 16584
rect 11060 16532 11112 16584
rect 8208 16464 8260 16516
rect 10508 16464 10560 16516
rect 15660 16532 15712 16584
rect 16212 16600 16264 16652
rect 16948 16668 17000 16720
rect 18144 16668 18196 16720
rect 18696 16668 18748 16720
rect 19064 16668 19116 16720
rect 23020 16736 23072 16788
rect 23204 16736 23256 16788
rect 23940 16736 23992 16788
rect 25504 16736 25556 16788
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 17040 16532 17092 16584
rect 12900 16464 12952 16516
rect 17500 16600 17552 16652
rect 18788 16643 18840 16652
rect 18788 16609 18797 16643
rect 18797 16609 18831 16643
rect 18831 16609 18840 16643
rect 18788 16600 18840 16609
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 18972 16532 19024 16584
rect 21272 16643 21324 16652
rect 21272 16609 21281 16643
rect 21281 16609 21315 16643
rect 21315 16609 21324 16643
rect 21272 16600 21324 16609
rect 24860 16668 24912 16720
rect 25044 16668 25096 16720
rect 30288 16736 30340 16788
rect 23204 16600 23256 16652
rect 23388 16643 23440 16652
rect 23388 16609 23397 16643
rect 23397 16609 23431 16643
rect 23431 16609 23440 16643
rect 23388 16600 23440 16609
rect 19524 16532 19576 16584
rect 19800 16532 19852 16584
rect 19892 16507 19944 16516
rect 19892 16473 19901 16507
rect 19901 16473 19935 16507
rect 19935 16473 19944 16507
rect 19892 16464 19944 16473
rect 5816 16396 5868 16448
rect 9772 16439 9824 16448
rect 9772 16405 9781 16439
rect 9781 16405 9815 16439
rect 9815 16405 9824 16439
rect 9772 16396 9824 16405
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 12808 16396 12860 16448
rect 16304 16396 16356 16448
rect 16856 16396 16908 16448
rect 17132 16396 17184 16448
rect 20352 16532 20404 16584
rect 20628 16532 20680 16584
rect 23020 16532 23072 16584
rect 23572 16600 23624 16652
rect 24216 16643 24268 16652
rect 24216 16609 24225 16643
rect 24225 16609 24259 16643
rect 24259 16609 24268 16643
rect 24216 16600 24268 16609
rect 24492 16643 24544 16652
rect 24492 16609 24526 16643
rect 24526 16609 24544 16643
rect 24492 16600 24544 16609
rect 25688 16643 25740 16652
rect 25688 16609 25697 16643
rect 25697 16609 25731 16643
rect 25731 16609 25740 16643
rect 25688 16600 25740 16609
rect 25872 16600 25924 16652
rect 25964 16643 26016 16652
rect 25964 16609 25973 16643
rect 25973 16609 26007 16643
rect 26007 16609 26016 16643
rect 25964 16600 26016 16609
rect 26056 16643 26108 16652
rect 26056 16609 26065 16643
rect 26065 16609 26099 16643
rect 26099 16609 26108 16643
rect 26056 16600 26108 16609
rect 26148 16600 26200 16652
rect 26792 16643 26844 16652
rect 26792 16609 26801 16643
rect 26801 16609 26835 16643
rect 26835 16609 26844 16643
rect 26792 16600 26844 16609
rect 25228 16532 25280 16584
rect 27436 16643 27488 16652
rect 27436 16609 27445 16643
rect 27445 16609 27479 16643
rect 27479 16609 27488 16643
rect 27436 16600 27488 16609
rect 27988 16600 28040 16652
rect 29092 16668 29144 16720
rect 29460 16668 29512 16720
rect 29920 16711 29972 16720
rect 29920 16677 29929 16711
rect 29929 16677 29963 16711
rect 29963 16677 29972 16711
rect 29920 16668 29972 16677
rect 29368 16600 29420 16652
rect 29644 16532 29696 16584
rect 23664 16464 23716 16516
rect 30564 16643 30616 16652
rect 30564 16609 30573 16643
rect 30573 16609 30607 16643
rect 30607 16609 30616 16643
rect 30564 16600 30616 16609
rect 30748 16643 30800 16652
rect 30748 16609 30757 16643
rect 30757 16609 30791 16643
rect 30791 16609 30800 16643
rect 30748 16600 30800 16609
rect 30288 16532 30340 16584
rect 20996 16396 21048 16448
rect 23204 16396 23256 16448
rect 24952 16396 25004 16448
rect 25688 16396 25740 16448
rect 27528 16396 27580 16448
rect 27988 16396 28040 16448
rect 29552 16439 29604 16448
rect 29552 16405 29561 16439
rect 29561 16405 29595 16439
rect 29595 16405 29604 16439
rect 29552 16396 29604 16405
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 11436 16294 11488 16346
rect 11500 16294 11552 16346
rect 11564 16294 11616 16346
rect 11628 16294 11680 16346
rect 11692 16294 11744 16346
rect 19210 16294 19262 16346
rect 19274 16294 19326 16346
rect 19338 16294 19390 16346
rect 19402 16294 19454 16346
rect 19466 16294 19518 16346
rect 26984 16294 27036 16346
rect 27048 16294 27100 16346
rect 27112 16294 27164 16346
rect 27176 16294 27228 16346
rect 27240 16294 27292 16346
rect 2964 16192 3016 16244
rect 4068 16192 4120 16244
rect 8116 16235 8168 16244
rect 8116 16201 8125 16235
rect 8125 16201 8159 16235
rect 8159 16201 8168 16235
rect 8116 16192 8168 16201
rect 2688 16124 2740 16176
rect 2872 16124 2924 16176
rect 3332 16124 3384 16176
rect 7012 16124 7064 16176
rect 7748 16124 7800 16176
rect 8484 16124 8536 16176
rect 9496 16235 9548 16244
rect 9496 16201 9505 16235
rect 9505 16201 9539 16235
rect 9539 16201 9548 16235
rect 9496 16192 9548 16201
rect 9772 16192 9824 16244
rect 1584 16056 1636 16108
rect 9680 16124 9732 16176
rect 2412 15988 2464 16040
rect 3332 16031 3384 16040
rect 3332 15997 3341 16031
rect 3341 15997 3375 16031
rect 3375 15997 3384 16031
rect 3332 15988 3384 15997
rect 4252 16031 4304 16040
rect 4252 15997 4261 16031
rect 4261 15997 4295 16031
rect 4295 15997 4304 16031
rect 4252 15988 4304 15997
rect 4160 15920 4212 15972
rect 2964 15852 3016 15904
rect 3884 15895 3936 15904
rect 3884 15861 3893 15895
rect 3893 15861 3927 15895
rect 3927 15861 3936 15895
rect 3884 15852 3936 15861
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 4068 15852 4120 15904
rect 5632 15988 5684 16040
rect 7748 16031 7800 16040
rect 7748 15997 7757 16031
rect 7757 15997 7791 16031
rect 7791 15997 7800 16031
rect 7748 15988 7800 15997
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 4712 15920 4764 15972
rect 6920 15920 6972 15972
rect 7564 15920 7616 15972
rect 8024 15988 8076 16040
rect 9036 15963 9088 15972
rect 9036 15929 9045 15963
rect 9045 15929 9079 15963
rect 9079 15929 9088 15963
rect 9036 15920 9088 15929
rect 9496 16056 9548 16108
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 10048 16235 10100 16244
rect 10048 16201 10057 16235
rect 10057 16201 10091 16235
rect 10091 16201 10100 16235
rect 10048 16192 10100 16201
rect 10416 16235 10468 16244
rect 10416 16201 10425 16235
rect 10425 16201 10459 16235
rect 10459 16201 10468 16235
rect 10416 16192 10468 16201
rect 10600 16192 10652 16244
rect 15568 16192 15620 16244
rect 10968 16124 11020 16176
rect 10324 15988 10376 16040
rect 10784 15988 10836 16040
rect 15292 16124 15344 16176
rect 16212 16235 16264 16244
rect 16212 16201 16221 16235
rect 16221 16201 16255 16235
rect 16255 16201 16264 16235
rect 16212 16192 16264 16201
rect 19708 16192 19760 16244
rect 11152 15988 11204 16040
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 10508 15920 10560 15972
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 11980 15920 12032 15972
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 13176 15988 13228 15997
rect 14096 15988 14148 16040
rect 15568 16031 15620 16040
rect 15568 15997 15577 16031
rect 15577 15997 15611 16031
rect 15611 15997 15620 16031
rect 15568 15988 15620 15997
rect 16120 16056 16172 16108
rect 16672 16099 16724 16108
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 16396 15988 16448 16040
rect 10968 15852 11020 15904
rect 11060 15852 11112 15904
rect 11520 15852 11572 15904
rect 15660 15852 15712 15904
rect 18236 15920 18288 15972
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 19616 15988 19668 16040
rect 21364 16099 21416 16108
rect 21364 16065 21373 16099
rect 21373 16065 21407 16099
rect 21407 16065 21416 16099
rect 21364 16056 21416 16065
rect 22928 16192 22980 16244
rect 23112 16124 23164 16176
rect 20260 15920 20312 15972
rect 20628 15988 20680 16040
rect 20812 16031 20864 16040
rect 20812 15997 20821 16031
rect 20821 15997 20855 16031
rect 20855 15997 20864 16031
rect 20812 15988 20864 15997
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 22100 15988 22152 15997
rect 22284 15988 22336 16040
rect 22376 16031 22428 16040
rect 22376 15997 22385 16031
rect 22385 15997 22419 16031
rect 22419 15997 22428 16031
rect 22376 15988 22428 15997
rect 22652 15988 22704 16040
rect 21088 15920 21140 15972
rect 21916 15920 21968 15972
rect 23204 16031 23256 16040
rect 23204 15997 23213 16031
rect 23213 15997 23247 16031
rect 23247 15997 23256 16031
rect 23204 15988 23256 15997
rect 23664 16056 23716 16108
rect 24492 16235 24544 16244
rect 24492 16201 24501 16235
rect 24501 16201 24535 16235
rect 24535 16201 24544 16235
rect 24492 16192 24544 16201
rect 26148 16235 26200 16244
rect 26148 16201 26157 16235
rect 26157 16201 26191 16235
rect 26191 16201 26200 16235
rect 26148 16192 26200 16201
rect 28632 16192 28684 16244
rect 30564 16192 30616 16244
rect 26792 16124 26844 16176
rect 23480 16031 23532 16040
rect 23480 15997 23489 16031
rect 23489 15997 23523 16031
rect 23523 15997 23532 16031
rect 23480 15988 23532 15997
rect 23848 16031 23900 16040
rect 23848 15997 23857 16031
rect 23857 15997 23891 16031
rect 23891 15997 23900 16031
rect 23848 15988 23900 15997
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 26056 16056 26108 16108
rect 26608 16056 26660 16108
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 25044 16031 25096 16040
rect 25044 15997 25078 16031
rect 25078 15997 25096 16031
rect 25044 15988 25096 15997
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 19524 15852 19576 15904
rect 19892 15852 19944 15904
rect 21456 15852 21508 15904
rect 22100 15852 22152 15904
rect 22928 15895 22980 15904
rect 22928 15861 22937 15895
rect 22937 15861 22971 15895
rect 22971 15861 22980 15895
rect 22928 15852 22980 15861
rect 23112 15852 23164 15904
rect 24952 15920 25004 15972
rect 26608 15963 26660 15972
rect 26608 15929 26617 15963
rect 26617 15929 26651 15963
rect 26651 15929 26660 15963
rect 26608 15920 26660 15929
rect 27344 15963 27396 15972
rect 27344 15929 27353 15963
rect 27353 15929 27387 15963
rect 27387 15929 27396 15963
rect 28172 16031 28224 16040
rect 28172 15997 28181 16031
rect 28181 15997 28215 16031
rect 28215 15997 28224 16031
rect 28172 15988 28224 15997
rect 29552 16056 29604 16108
rect 29092 15988 29144 16040
rect 29276 16031 29328 16040
rect 29276 15997 29285 16031
rect 29285 15997 29319 16031
rect 29319 15997 29328 16031
rect 29276 15988 29328 15997
rect 29368 16031 29420 16040
rect 29368 15997 29377 16031
rect 29377 15997 29411 16031
rect 29411 15997 29420 16031
rect 29368 15988 29420 15997
rect 29920 16031 29972 16040
rect 29920 15997 29929 16031
rect 29929 15997 29963 16031
rect 29963 15997 29972 16031
rect 29920 15988 29972 15997
rect 27344 15920 27396 15929
rect 24584 15852 24636 15904
rect 29920 15852 29972 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 12096 15750 12148 15802
rect 12160 15750 12212 15802
rect 12224 15750 12276 15802
rect 12288 15750 12340 15802
rect 12352 15750 12404 15802
rect 19870 15750 19922 15802
rect 19934 15750 19986 15802
rect 19998 15750 20050 15802
rect 20062 15750 20114 15802
rect 20126 15750 20178 15802
rect 27644 15750 27696 15802
rect 27708 15750 27760 15802
rect 27772 15750 27824 15802
rect 27836 15750 27888 15802
rect 27900 15750 27952 15802
rect 2964 15648 3016 15700
rect 3884 15648 3936 15700
rect 3976 15580 4028 15632
rect 4160 15623 4212 15632
rect 4160 15589 4169 15623
rect 4169 15589 4203 15623
rect 4203 15589 4212 15623
rect 4160 15580 4212 15589
rect 4712 15648 4764 15700
rect 6920 15648 6972 15700
rect 7840 15648 7892 15700
rect 7196 15580 7248 15632
rect 9588 15623 9640 15632
rect 1676 15512 1728 15564
rect 3700 15555 3752 15564
rect 3700 15521 3709 15555
rect 3709 15521 3743 15555
rect 3743 15521 3752 15555
rect 3700 15512 3752 15521
rect 3792 15555 3844 15564
rect 3792 15521 3801 15555
rect 3801 15521 3835 15555
rect 3835 15521 3844 15555
rect 3792 15512 3844 15521
rect 3148 15444 3200 15496
rect 2964 15376 3016 15428
rect 3424 15376 3476 15428
rect 5632 15512 5684 15564
rect 9588 15589 9597 15623
rect 9597 15589 9631 15623
rect 9631 15589 9640 15623
rect 9588 15580 9640 15589
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 6000 15444 6052 15496
rect 8484 15512 8536 15564
rect 4252 15376 4304 15428
rect 4804 15376 4856 15428
rect 9036 15444 9088 15496
rect 13636 15648 13688 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 10324 15580 10376 15632
rect 9956 15512 10008 15564
rect 10232 15512 10284 15564
rect 2872 15308 2924 15360
rect 3516 15308 3568 15360
rect 3792 15308 3844 15360
rect 4068 15308 4120 15360
rect 4988 15351 5040 15360
rect 4988 15317 4997 15351
rect 4997 15317 5031 15351
rect 5031 15317 5040 15351
rect 4988 15308 5040 15317
rect 6736 15308 6788 15360
rect 10600 15555 10652 15564
rect 10600 15521 10609 15555
rect 10609 15521 10643 15555
rect 10643 15521 10652 15555
rect 10600 15512 10652 15521
rect 10784 15512 10836 15564
rect 11520 15555 11572 15564
rect 11520 15521 11529 15555
rect 11529 15521 11563 15555
rect 11563 15521 11572 15555
rect 11520 15512 11572 15521
rect 10968 15444 11020 15496
rect 14648 15555 14700 15564
rect 14648 15521 14657 15555
rect 14657 15521 14691 15555
rect 14691 15521 14700 15555
rect 14648 15512 14700 15521
rect 16028 15512 16080 15564
rect 15384 15444 15436 15496
rect 9680 15376 9732 15428
rect 10140 15376 10192 15428
rect 10232 15419 10284 15428
rect 10232 15385 10241 15419
rect 10241 15385 10275 15419
rect 10275 15385 10284 15419
rect 10232 15376 10284 15385
rect 10508 15376 10560 15428
rect 10692 15376 10744 15428
rect 12624 15376 12676 15428
rect 14004 15376 14056 15428
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 7932 15308 7984 15360
rect 11060 15308 11112 15360
rect 11152 15308 11204 15360
rect 11980 15308 12032 15360
rect 15568 15308 15620 15360
rect 17960 15648 18012 15700
rect 18236 15691 18288 15700
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 19064 15691 19116 15700
rect 19064 15657 19073 15691
rect 19073 15657 19107 15691
rect 19107 15657 19116 15691
rect 19064 15648 19116 15657
rect 17500 15580 17552 15632
rect 18972 15580 19024 15632
rect 20720 15648 20772 15700
rect 21088 15648 21140 15700
rect 22468 15648 22520 15700
rect 22744 15648 22796 15700
rect 23112 15648 23164 15700
rect 23664 15648 23716 15700
rect 24676 15648 24728 15700
rect 24768 15648 24820 15700
rect 20812 15580 20864 15632
rect 21272 15580 21324 15632
rect 26608 15580 26660 15632
rect 28264 15648 28316 15700
rect 29092 15648 29144 15700
rect 29276 15648 29328 15700
rect 16856 15555 16908 15564
rect 16856 15521 16865 15555
rect 16865 15521 16899 15555
rect 16899 15521 16908 15555
rect 16856 15512 16908 15521
rect 16948 15512 17000 15564
rect 17960 15512 18012 15564
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 19524 15555 19576 15564
rect 19524 15521 19533 15555
rect 19533 15521 19567 15555
rect 19567 15521 19576 15555
rect 19524 15512 19576 15521
rect 19800 15555 19852 15564
rect 19800 15521 19809 15555
rect 19809 15521 19843 15555
rect 19843 15521 19852 15555
rect 19800 15512 19852 15521
rect 20536 15512 20588 15564
rect 20720 15555 20772 15564
rect 20720 15521 20729 15555
rect 20729 15521 20763 15555
rect 20763 15521 20772 15555
rect 20720 15512 20772 15521
rect 20996 15555 21048 15564
rect 20996 15521 21005 15555
rect 21005 15521 21039 15555
rect 21039 15521 21048 15555
rect 20996 15512 21048 15521
rect 21456 15555 21508 15564
rect 21456 15521 21465 15555
rect 21465 15521 21499 15555
rect 21499 15521 21508 15555
rect 21456 15512 21508 15521
rect 19616 15444 19668 15496
rect 21824 15555 21876 15564
rect 21824 15521 21833 15555
rect 21833 15521 21867 15555
rect 21867 15521 21876 15555
rect 21824 15512 21876 15521
rect 22100 15555 22152 15564
rect 22100 15521 22109 15555
rect 22109 15521 22143 15555
rect 22143 15521 22152 15555
rect 22100 15512 22152 15521
rect 23388 15512 23440 15564
rect 23296 15444 23348 15496
rect 24492 15512 24544 15564
rect 24860 15555 24912 15564
rect 24860 15521 24869 15555
rect 24869 15521 24903 15555
rect 24903 15521 24912 15555
rect 24860 15512 24912 15521
rect 24400 15444 24452 15496
rect 24676 15444 24728 15496
rect 25780 15512 25832 15564
rect 27988 15512 28040 15564
rect 28448 15555 28500 15564
rect 28448 15521 28457 15555
rect 28457 15521 28491 15555
rect 28491 15521 28500 15555
rect 28448 15512 28500 15521
rect 29000 15512 29052 15564
rect 29092 15555 29144 15564
rect 29092 15521 29101 15555
rect 29101 15521 29135 15555
rect 29135 15521 29144 15555
rect 29092 15512 29144 15521
rect 29184 15555 29236 15564
rect 29184 15521 29193 15555
rect 29193 15521 29227 15555
rect 29227 15521 29236 15555
rect 29184 15512 29236 15521
rect 29276 15555 29328 15564
rect 29276 15521 29290 15555
rect 29290 15521 29324 15555
rect 29324 15521 29328 15555
rect 29276 15512 29328 15521
rect 29460 15555 29512 15564
rect 29460 15521 29469 15555
rect 29469 15521 29503 15555
rect 29503 15521 29512 15555
rect 29460 15512 29512 15521
rect 19064 15376 19116 15428
rect 20628 15376 20680 15428
rect 21640 15376 21692 15428
rect 22744 15376 22796 15428
rect 29092 15376 29144 15428
rect 16672 15308 16724 15360
rect 20812 15308 20864 15360
rect 21456 15308 21508 15360
rect 24584 15308 24636 15360
rect 25412 15308 25464 15360
rect 25688 15308 25740 15360
rect 28540 15308 28592 15360
rect 30656 15308 30708 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 11436 15206 11488 15258
rect 11500 15206 11552 15258
rect 11564 15206 11616 15258
rect 11628 15206 11680 15258
rect 11692 15206 11744 15258
rect 19210 15206 19262 15258
rect 19274 15206 19326 15258
rect 19338 15206 19390 15258
rect 19402 15206 19454 15258
rect 19466 15206 19518 15258
rect 26984 15206 27036 15258
rect 27048 15206 27100 15258
rect 27112 15206 27164 15258
rect 27176 15206 27228 15258
rect 27240 15206 27292 15258
rect 4896 15104 4948 15156
rect 5540 15104 5592 15156
rect 5632 15104 5684 15156
rect 4712 15036 4764 15088
rect 1584 14900 1636 14952
rect 1952 14943 2004 14952
rect 1952 14909 1961 14943
rect 1961 14909 1995 14943
rect 1995 14909 2004 14943
rect 1952 14900 2004 14909
rect 4160 14968 4212 15020
rect 2596 14943 2648 14952
rect 2596 14909 2605 14943
rect 2605 14909 2639 14943
rect 2639 14909 2648 14943
rect 2596 14900 2648 14909
rect 2780 14900 2832 14952
rect 3056 14900 3108 14952
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 5540 14968 5592 15020
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 3424 14832 3476 14884
rect 7196 14900 7248 14952
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 9588 15104 9640 15156
rect 10324 15104 10376 15156
rect 10416 15104 10468 15156
rect 10048 15079 10100 15088
rect 10048 15045 10057 15079
rect 10057 15045 10091 15079
rect 10091 15045 10100 15079
rect 10048 15036 10100 15045
rect 13728 15104 13780 15156
rect 15292 15104 15344 15156
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 16396 15147 16448 15156
rect 16396 15113 16405 15147
rect 16405 15113 16439 15147
rect 16439 15113 16448 15147
rect 16396 15104 16448 15113
rect 16580 15104 16632 15156
rect 21272 15104 21324 15156
rect 25964 15104 26016 15156
rect 26700 15104 26752 15156
rect 29000 15104 29052 15156
rect 29460 15104 29512 15156
rect 9036 14968 9088 15020
rect 6184 14832 6236 14884
rect 1676 14764 1728 14816
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 3608 14764 3660 14816
rect 4252 14764 4304 14816
rect 6920 14832 6972 14884
rect 8300 14900 8352 14952
rect 9496 14943 9548 14952
rect 9496 14909 9505 14943
rect 9505 14909 9539 14943
rect 9539 14909 9548 14943
rect 9496 14900 9548 14909
rect 9864 14968 9916 15020
rect 10692 14968 10744 15020
rect 10140 14900 10192 14952
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 10876 14900 10928 14952
rect 10968 14943 11020 14952
rect 10968 14909 10977 14943
rect 10977 14909 11011 14943
rect 11011 14909 11020 14943
rect 10968 14900 11020 14909
rect 15844 15036 15896 15088
rect 16948 15036 17000 15088
rect 19616 15036 19668 15088
rect 20720 15036 20772 15088
rect 21916 15036 21968 15088
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 15384 14968 15436 15020
rect 13176 14900 13228 14952
rect 13636 14943 13688 14952
rect 13636 14909 13645 14943
rect 13645 14909 13679 14943
rect 13679 14909 13688 14943
rect 13636 14900 13688 14909
rect 15752 14943 15804 14952
rect 15752 14909 15761 14943
rect 15761 14909 15795 14943
rect 15795 14909 15804 14943
rect 15752 14900 15804 14909
rect 16488 14968 16540 15020
rect 10508 14832 10560 14884
rect 7012 14764 7064 14816
rect 7104 14764 7156 14816
rect 7380 14764 7432 14816
rect 11244 14764 11296 14816
rect 13544 14832 13596 14884
rect 14372 14832 14424 14884
rect 11888 14764 11940 14816
rect 14096 14764 14148 14816
rect 16856 14900 16908 14952
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 17224 14900 17276 14952
rect 16120 14832 16172 14884
rect 17592 14943 17644 14952
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 19340 14968 19392 15020
rect 22560 15036 22612 15088
rect 22928 15036 22980 15088
rect 23664 15036 23716 15088
rect 24124 15036 24176 15088
rect 26792 15036 26844 15088
rect 27160 15036 27212 15088
rect 27436 15036 27488 15088
rect 28356 15036 28408 15088
rect 29276 15036 29328 15088
rect 30564 15036 30616 15088
rect 17776 14832 17828 14884
rect 16948 14764 17000 14816
rect 17868 14764 17920 14816
rect 19616 14900 19668 14952
rect 21548 14900 21600 14952
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 22928 14943 22980 14952
rect 18880 14832 18932 14884
rect 20628 14832 20680 14884
rect 21456 14832 21508 14884
rect 22928 14909 22937 14943
rect 22937 14909 22971 14943
rect 22971 14909 22980 14943
rect 22928 14900 22980 14909
rect 24124 14900 24176 14952
rect 24492 14968 24544 15020
rect 26700 14968 26752 15020
rect 29000 14968 29052 15020
rect 29644 15011 29696 15020
rect 29644 14977 29653 15011
rect 29653 14977 29687 15011
rect 29687 14977 29696 15011
rect 29644 14968 29696 14977
rect 29736 14968 29788 15020
rect 24400 14943 24452 14952
rect 24400 14909 24409 14943
rect 24409 14909 24443 14943
rect 24443 14909 24452 14943
rect 24400 14900 24452 14909
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24952 14943 25004 14952
rect 24952 14909 24961 14943
rect 24961 14909 24995 14943
rect 24995 14909 25004 14943
rect 24952 14900 25004 14909
rect 25044 14943 25096 14952
rect 25044 14909 25053 14943
rect 25053 14909 25087 14943
rect 25087 14909 25096 14943
rect 25044 14900 25096 14909
rect 25228 14943 25280 14952
rect 25228 14909 25237 14943
rect 25237 14909 25271 14943
rect 25271 14909 25280 14943
rect 25228 14900 25280 14909
rect 25136 14832 25188 14884
rect 26884 14900 26936 14952
rect 25596 14832 25648 14884
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27436 14900 27488 14909
rect 27988 14900 28040 14952
rect 28632 14943 28684 14952
rect 28632 14909 28641 14943
rect 28641 14909 28675 14943
rect 28675 14909 28684 14943
rect 28632 14900 28684 14909
rect 29552 14943 29604 14952
rect 29552 14909 29561 14943
rect 29561 14909 29595 14943
rect 29595 14909 29604 14943
rect 29552 14900 29604 14909
rect 30472 14943 30524 14952
rect 30472 14909 30481 14943
rect 30481 14909 30515 14943
rect 30515 14909 30524 14943
rect 30472 14900 30524 14909
rect 30656 14943 30708 14952
rect 30656 14909 30665 14943
rect 30665 14909 30699 14943
rect 30699 14909 30708 14943
rect 30656 14900 30708 14909
rect 28448 14832 28500 14884
rect 29920 14875 29972 14884
rect 29920 14841 29929 14875
rect 29929 14841 29963 14875
rect 29963 14841 29972 14875
rect 29920 14832 29972 14841
rect 30196 14832 30248 14884
rect 30840 14943 30892 14952
rect 30840 14909 30849 14943
rect 30849 14909 30883 14943
rect 30883 14909 30892 14943
rect 30840 14900 30892 14909
rect 20996 14764 21048 14816
rect 22652 14764 22704 14816
rect 23388 14807 23440 14816
rect 23388 14773 23397 14807
rect 23397 14773 23431 14807
rect 23431 14773 23440 14807
rect 23388 14764 23440 14773
rect 24216 14764 24268 14816
rect 25504 14807 25556 14816
rect 25504 14773 25513 14807
rect 25513 14773 25547 14807
rect 25547 14773 25556 14807
rect 25504 14764 25556 14773
rect 25872 14764 25924 14816
rect 27252 14764 27304 14816
rect 27528 14764 27580 14816
rect 29092 14764 29144 14816
rect 29276 14764 29328 14816
rect 29828 14764 29880 14816
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 12096 14662 12148 14714
rect 12160 14662 12212 14714
rect 12224 14662 12276 14714
rect 12288 14662 12340 14714
rect 12352 14662 12404 14714
rect 19870 14662 19922 14714
rect 19934 14662 19986 14714
rect 19998 14662 20050 14714
rect 20062 14662 20114 14714
rect 20126 14662 20178 14714
rect 27644 14662 27696 14714
rect 27708 14662 27760 14714
rect 27772 14662 27824 14714
rect 27836 14662 27888 14714
rect 27900 14662 27952 14714
rect 3424 14560 3476 14612
rect 5540 14603 5592 14612
rect 5540 14569 5549 14603
rect 5549 14569 5583 14603
rect 5583 14569 5592 14603
rect 5540 14560 5592 14569
rect 7104 14603 7156 14612
rect 7104 14569 7113 14603
rect 7113 14569 7147 14603
rect 7147 14569 7156 14603
rect 7104 14560 7156 14569
rect 7564 14560 7616 14612
rect 10416 14560 10468 14612
rect 10600 14560 10652 14612
rect 12716 14560 12768 14612
rect 13268 14603 13320 14612
rect 13268 14569 13277 14603
rect 13277 14569 13311 14603
rect 13311 14569 13320 14603
rect 13268 14560 13320 14569
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 2228 14492 2280 14544
rect 1676 14467 1728 14476
rect 1676 14433 1685 14467
rect 1685 14433 1719 14467
rect 1719 14433 1728 14467
rect 1676 14424 1728 14433
rect 3240 14288 3292 14340
rect 3148 14263 3200 14272
rect 3148 14229 3157 14263
rect 3157 14229 3191 14263
rect 3191 14229 3200 14263
rect 3148 14220 3200 14229
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 3608 14467 3660 14476
rect 3608 14433 3617 14467
rect 3617 14433 3651 14467
rect 3651 14433 3660 14467
rect 3608 14424 3660 14433
rect 4988 14492 5040 14544
rect 5908 14492 5960 14544
rect 4252 14424 4304 14476
rect 6000 14467 6052 14476
rect 6000 14433 6009 14467
rect 6009 14433 6043 14467
rect 6043 14433 6052 14467
rect 6000 14424 6052 14433
rect 9036 14492 9088 14544
rect 10140 14492 10192 14544
rect 10692 14492 10744 14544
rect 11888 14535 11940 14544
rect 11888 14501 11897 14535
rect 11897 14501 11931 14535
rect 11931 14501 11940 14535
rect 11888 14492 11940 14501
rect 11980 14492 12032 14544
rect 13544 14492 13596 14544
rect 15200 14492 15252 14544
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 6920 14356 6972 14408
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 10508 14424 10560 14476
rect 10876 14424 10928 14476
rect 11244 14467 11296 14476
rect 11244 14433 11253 14467
rect 11253 14433 11287 14467
rect 11287 14433 11296 14467
rect 11244 14424 11296 14433
rect 11152 14356 11204 14408
rect 6644 14263 6696 14272
rect 6644 14229 6653 14263
rect 6653 14229 6687 14263
rect 6687 14229 6696 14263
rect 6644 14220 6696 14229
rect 9588 14288 9640 14340
rect 11612 14424 11664 14476
rect 17316 14560 17368 14612
rect 19064 14603 19116 14612
rect 19064 14569 19073 14603
rect 19073 14569 19107 14603
rect 19107 14569 19116 14603
rect 19064 14560 19116 14569
rect 21364 14560 21416 14612
rect 22376 14560 22428 14612
rect 23572 14560 23624 14612
rect 24492 14603 24544 14612
rect 24492 14569 24501 14603
rect 24501 14569 24535 14603
rect 24535 14569 24544 14603
rect 24492 14560 24544 14569
rect 25044 14560 25096 14612
rect 26332 14560 26384 14612
rect 18420 14492 18472 14544
rect 12808 14424 12860 14476
rect 13728 14467 13780 14476
rect 13728 14433 13737 14467
rect 13737 14433 13771 14467
rect 13771 14433 13780 14467
rect 13728 14424 13780 14433
rect 7196 14220 7248 14272
rect 7472 14263 7524 14272
rect 7472 14229 7481 14263
rect 7481 14229 7515 14263
rect 7515 14229 7524 14263
rect 7472 14220 7524 14229
rect 9956 14220 10008 14272
rect 13820 14356 13872 14408
rect 14004 14467 14056 14476
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 14556 14424 14608 14476
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 16304 14424 16356 14476
rect 17868 14424 17920 14476
rect 18328 14467 18380 14476
rect 18328 14433 18341 14467
rect 18341 14433 18380 14467
rect 21272 14492 21324 14544
rect 18328 14424 18380 14433
rect 18972 14467 19024 14476
rect 18972 14433 18981 14467
rect 18981 14433 19015 14467
rect 19015 14433 19024 14467
rect 18972 14424 19024 14433
rect 16764 14356 16816 14408
rect 16856 14356 16908 14408
rect 19616 14424 19668 14476
rect 19340 14399 19392 14408
rect 19340 14365 19349 14399
rect 19349 14365 19383 14399
rect 19383 14365 19392 14399
rect 19340 14356 19392 14365
rect 19892 14356 19944 14408
rect 20812 14467 20864 14476
rect 20812 14433 20821 14467
rect 20821 14433 20855 14467
rect 20855 14433 20864 14467
rect 20812 14424 20864 14433
rect 21640 14424 21692 14476
rect 21916 14424 21968 14476
rect 22836 14424 22888 14476
rect 25504 14492 25556 14544
rect 23664 14467 23716 14476
rect 23664 14433 23673 14467
rect 23673 14433 23707 14467
rect 23707 14433 23716 14467
rect 23664 14424 23716 14433
rect 23756 14467 23808 14476
rect 23756 14433 23765 14467
rect 23765 14433 23799 14467
rect 23799 14433 23808 14467
rect 23756 14424 23808 14433
rect 23848 14424 23900 14476
rect 24308 14424 24360 14476
rect 21548 14356 21600 14408
rect 22008 14356 22060 14408
rect 23204 14356 23256 14408
rect 24124 14356 24176 14408
rect 24584 14424 24636 14476
rect 24768 14424 24820 14476
rect 25228 14424 25280 14476
rect 25872 14467 25924 14476
rect 25872 14433 25881 14467
rect 25881 14433 25915 14467
rect 25915 14433 25924 14467
rect 25872 14424 25924 14433
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 26148 14424 26200 14476
rect 27160 14560 27212 14612
rect 27436 14560 27488 14612
rect 29368 14603 29420 14612
rect 29368 14569 29377 14603
rect 29377 14569 29411 14603
rect 29411 14569 29420 14603
rect 29368 14560 29420 14569
rect 30932 14560 30984 14612
rect 26608 14492 26660 14544
rect 24676 14399 24728 14408
rect 24676 14365 24685 14399
rect 24685 14365 24719 14399
rect 24719 14365 24728 14399
rect 24676 14356 24728 14365
rect 26792 14467 26844 14476
rect 26792 14433 26801 14467
rect 26801 14433 26835 14467
rect 26835 14433 26844 14467
rect 26792 14424 26844 14433
rect 26976 14424 27028 14476
rect 11612 14288 11664 14340
rect 15752 14288 15804 14340
rect 16948 14288 17000 14340
rect 17408 14288 17460 14340
rect 12716 14220 12768 14272
rect 14188 14220 14240 14272
rect 16212 14220 16264 14272
rect 17500 14220 17552 14272
rect 22100 14288 22152 14340
rect 18328 14220 18380 14272
rect 19064 14263 19116 14272
rect 19064 14229 19073 14263
rect 19073 14229 19107 14263
rect 19107 14229 19116 14263
rect 19064 14220 19116 14229
rect 22468 14263 22520 14272
rect 22468 14229 22477 14263
rect 22477 14229 22511 14263
rect 22511 14229 22520 14263
rect 22468 14220 22520 14229
rect 25228 14288 25280 14340
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 23940 14220 23992 14272
rect 24308 14220 24360 14272
rect 26148 14288 26200 14340
rect 26332 14288 26384 14340
rect 26792 14288 26844 14340
rect 27160 14467 27212 14476
rect 27160 14433 27169 14467
rect 27169 14433 27203 14467
rect 27203 14433 27212 14467
rect 27160 14424 27212 14433
rect 27252 14424 27304 14476
rect 29184 14492 29236 14544
rect 27528 14467 27580 14476
rect 27528 14433 27537 14467
rect 27537 14433 27571 14467
rect 27571 14433 27580 14467
rect 27528 14424 27580 14433
rect 27804 14424 27856 14476
rect 28264 14467 28316 14476
rect 28264 14433 28273 14467
rect 28273 14433 28307 14467
rect 28307 14433 28316 14467
rect 28264 14424 28316 14433
rect 28356 14467 28408 14476
rect 28356 14433 28365 14467
rect 28365 14433 28399 14467
rect 28399 14433 28408 14467
rect 28356 14424 28408 14433
rect 28540 14467 28592 14476
rect 28540 14433 28549 14467
rect 28549 14433 28583 14467
rect 28583 14433 28592 14467
rect 28540 14424 28592 14433
rect 28632 14424 28684 14476
rect 27896 14356 27948 14408
rect 27988 14288 28040 14340
rect 25596 14263 25648 14272
rect 25596 14229 25605 14263
rect 25605 14229 25639 14263
rect 25639 14229 25648 14263
rect 25596 14220 25648 14229
rect 25688 14220 25740 14272
rect 27712 14220 27764 14272
rect 29000 14356 29052 14408
rect 29184 14356 29236 14408
rect 29644 14356 29696 14408
rect 30472 14467 30524 14476
rect 30472 14433 30481 14467
rect 30481 14433 30515 14467
rect 30515 14433 30524 14467
rect 30472 14424 30524 14433
rect 30564 14424 30616 14476
rect 29276 14288 29328 14340
rect 29000 14220 29052 14272
rect 29092 14220 29144 14272
rect 30104 14220 30156 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 11436 14118 11488 14170
rect 11500 14118 11552 14170
rect 11564 14118 11616 14170
rect 11628 14118 11680 14170
rect 11692 14118 11744 14170
rect 19210 14118 19262 14170
rect 19274 14118 19326 14170
rect 19338 14118 19390 14170
rect 19402 14118 19454 14170
rect 19466 14118 19518 14170
rect 26984 14118 27036 14170
rect 27048 14118 27100 14170
rect 27112 14118 27164 14170
rect 27176 14118 27228 14170
rect 27240 14118 27292 14170
rect 1952 14016 2004 14068
rect 3056 14059 3108 14068
rect 3056 14025 3065 14059
rect 3065 14025 3099 14059
rect 3099 14025 3108 14059
rect 3056 14016 3108 14025
rect 5540 14016 5592 14068
rect 6000 14016 6052 14068
rect 10600 14016 10652 14068
rect 11244 14016 11296 14068
rect 3240 13880 3292 13932
rect 11980 13948 12032 14000
rect 3148 13812 3200 13864
rect 6184 13855 6236 13864
rect 6184 13821 6193 13855
rect 6193 13821 6227 13855
rect 6227 13821 6236 13855
rect 6184 13812 6236 13821
rect 7472 13812 7524 13864
rect 11888 13812 11940 13864
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 12900 13812 12952 13864
rect 14004 13948 14056 14000
rect 16304 14016 16356 14068
rect 18972 14016 19024 14068
rect 19248 14016 19300 14068
rect 13452 13812 13504 13864
rect 13728 13812 13780 13864
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 17776 13948 17828 14000
rect 17960 13948 18012 14000
rect 17500 13880 17552 13932
rect 4712 13744 4764 13796
rect 10048 13744 10100 13796
rect 12716 13744 12768 13796
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 15752 13812 15804 13864
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 17040 13812 17092 13864
rect 17960 13855 18012 13864
rect 17960 13821 17969 13855
rect 17969 13821 18003 13855
rect 18003 13821 18012 13855
rect 17960 13812 18012 13821
rect 18420 13880 18472 13932
rect 19248 13880 19300 13932
rect 19800 13812 19852 13864
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 21640 14016 21692 14068
rect 22836 14016 22888 14068
rect 24584 14016 24636 14068
rect 25228 14059 25280 14068
rect 25228 14025 25237 14059
rect 25237 14025 25271 14059
rect 25271 14025 25280 14059
rect 25228 14016 25280 14025
rect 26700 14059 26752 14068
rect 26700 14025 26709 14059
rect 26709 14025 26743 14059
rect 26743 14025 26752 14059
rect 26700 14016 26752 14025
rect 26884 14016 26936 14068
rect 20720 13880 20772 13932
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 6092 13719 6144 13728
rect 6092 13685 6101 13719
rect 6101 13685 6135 13719
rect 6135 13685 6144 13719
rect 6092 13676 6144 13685
rect 7472 13676 7524 13728
rect 7932 13676 7984 13728
rect 11796 13676 11848 13728
rect 15200 13744 15252 13796
rect 16120 13744 16172 13796
rect 15476 13676 15528 13728
rect 15936 13676 15988 13728
rect 16396 13719 16448 13728
rect 16396 13685 16405 13719
rect 16405 13685 16439 13719
rect 16439 13685 16448 13719
rect 16396 13676 16448 13685
rect 16856 13744 16908 13796
rect 20996 13812 21048 13864
rect 22284 13812 22336 13864
rect 22744 13855 22796 13864
rect 22744 13821 22753 13855
rect 22753 13821 22787 13855
rect 22787 13821 22796 13855
rect 22744 13812 22796 13821
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 23204 13880 23256 13932
rect 23296 13880 23348 13932
rect 29276 14016 29328 14068
rect 30472 14016 30524 14068
rect 30932 14059 30984 14068
rect 30932 14025 30941 14059
rect 30941 14025 30975 14059
rect 30975 14025 30984 14059
rect 30932 14016 30984 14025
rect 23572 13812 23624 13864
rect 21088 13744 21140 13796
rect 21732 13744 21784 13796
rect 22192 13744 22244 13796
rect 24860 13812 24912 13864
rect 25320 13855 25372 13864
rect 25320 13821 25329 13855
rect 25329 13821 25363 13855
rect 25363 13821 25372 13855
rect 25320 13812 25372 13821
rect 25596 13855 25648 13864
rect 25596 13821 25630 13855
rect 25630 13821 25648 13855
rect 25596 13812 25648 13821
rect 26332 13812 26384 13864
rect 27344 13812 27396 13864
rect 27712 13923 27764 13932
rect 27712 13889 27721 13923
rect 27721 13889 27755 13923
rect 27755 13889 27764 13923
rect 27712 13880 27764 13889
rect 27804 13812 27856 13864
rect 27896 13812 27948 13864
rect 28264 13812 28316 13864
rect 29184 13948 29236 14000
rect 29460 13880 29512 13932
rect 29092 13812 29144 13864
rect 29368 13812 29420 13864
rect 29552 13855 29604 13864
rect 29552 13821 29561 13855
rect 29561 13821 29595 13855
rect 29595 13821 29604 13855
rect 29552 13812 29604 13821
rect 29828 13855 29880 13864
rect 29828 13821 29862 13855
rect 29862 13821 29880 13855
rect 29828 13812 29880 13821
rect 31024 13855 31076 13864
rect 31024 13821 31033 13855
rect 31033 13821 31067 13855
rect 31067 13821 31076 13855
rect 31024 13812 31076 13821
rect 22928 13676 22980 13728
rect 23388 13676 23440 13728
rect 26976 13719 27028 13728
rect 26976 13685 26985 13719
rect 26985 13685 27019 13719
rect 27019 13685 27028 13719
rect 26976 13676 27028 13685
rect 29920 13744 29972 13796
rect 28816 13676 28868 13728
rect 31116 13719 31168 13728
rect 31116 13685 31125 13719
rect 31125 13685 31159 13719
rect 31159 13685 31168 13719
rect 31116 13676 31168 13685
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 12096 13574 12148 13626
rect 12160 13574 12212 13626
rect 12224 13574 12276 13626
rect 12288 13574 12340 13626
rect 12352 13574 12404 13626
rect 19870 13574 19922 13626
rect 19934 13574 19986 13626
rect 19998 13574 20050 13626
rect 20062 13574 20114 13626
rect 20126 13574 20178 13626
rect 27644 13574 27696 13626
rect 27708 13574 27760 13626
rect 27772 13574 27824 13626
rect 27836 13574 27888 13626
rect 27900 13574 27952 13626
rect 2780 13472 2832 13524
rect 3240 13404 3292 13456
rect 4160 13472 4212 13524
rect 7196 13472 7248 13524
rect 6644 13404 6696 13456
rect 6920 13404 6972 13456
rect 5724 13268 5776 13320
rect 3516 13132 3568 13184
rect 6092 13336 6144 13388
rect 7104 13336 7156 13388
rect 7840 13379 7892 13388
rect 7840 13345 7849 13379
rect 7849 13345 7883 13379
rect 7883 13345 7892 13379
rect 7840 13336 7892 13345
rect 7472 13268 7524 13320
rect 8208 13268 8260 13320
rect 9588 13404 9640 13456
rect 12900 13472 12952 13524
rect 13268 13472 13320 13524
rect 13912 13472 13964 13524
rect 14004 13472 14056 13524
rect 15568 13472 15620 13524
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 16856 13515 16908 13524
rect 16856 13481 16865 13515
rect 16865 13481 16899 13515
rect 16899 13481 16908 13515
rect 16856 13472 16908 13481
rect 17040 13515 17092 13524
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 18880 13472 18932 13524
rect 20076 13472 20128 13524
rect 20536 13472 20588 13524
rect 21732 13515 21784 13524
rect 21732 13481 21741 13515
rect 21741 13481 21775 13515
rect 21775 13481 21784 13515
rect 21732 13472 21784 13481
rect 22192 13472 22244 13524
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 23756 13515 23808 13524
rect 23756 13481 23765 13515
rect 23765 13481 23799 13515
rect 23799 13481 23808 13515
rect 23756 13472 23808 13481
rect 24400 13472 24452 13524
rect 24860 13515 24912 13524
rect 24860 13481 24869 13515
rect 24869 13481 24903 13515
rect 24903 13481 24912 13515
rect 24860 13472 24912 13481
rect 25136 13515 25188 13524
rect 25136 13481 25145 13515
rect 25145 13481 25179 13515
rect 25179 13481 25188 13515
rect 25136 13472 25188 13481
rect 25320 13472 25372 13524
rect 26792 13515 26844 13524
rect 26792 13481 26801 13515
rect 26801 13481 26835 13515
rect 26835 13481 26844 13515
rect 26792 13472 26844 13481
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 9956 13336 10008 13388
rect 15200 13447 15252 13456
rect 15200 13413 15209 13447
rect 15209 13413 15243 13447
rect 15243 13413 15252 13447
rect 15200 13404 15252 13413
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 10416 13336 10468 13388
rect 13268 13336 13320 13388
rect 9772 13268 9824 13320
rect 11244 13268 11296 13320
rect 11888 13268 11940 13320
rect 14648 13336 14700 13388
rect 14924 13336 14976 13388
rect 15936 13404 15988 13456
rect 17224 13404 17276 13456
rect 7104 13132 7156 13184
rect 12992 13200 13044 13252
rect 9036 13132 9088 13184
rect 10140 13132 10192 13184
rect 10232 13132 10284 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 12808 13132 12860 13184
rect 13912 13268 13964 13320
rect 16396 13379 16448 13388
rect 16396 13345 16405 13379
rect 16405 13345 16439 13379
rect 16439 13345 16448 13379
rect 16396 13336 16448 13345
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 16764 13336 16816 13388
rect 17868 13336 17920 13388
rect 22100 13447 22152 13456
rect 22100 13413 22109 13447
rect 22109 13413 22143 13447
rect 22143 13413 22152 13447
rect 22100 13404 22152 13413
rect 17040 13268 17092 13320
rect 16028 13200 16080 13252
rect 19708 13336 19760 13388
rect 20076 13379 20128 13388
rect 20076 13345 20085 13379
rect 20085 13345 20119 13379
rect 20119 13345 20128 13379
rect 20076 13336 20128 13345
rect 20444 13268 20496 13320
rect 20720 13243 20772 13252
rect 20720 13209 20729 13243
rect 20729 13209 20763 13243
rect 20763 13209 20772 13243
rect 20720 13200 20772 13209
rect 21640 13379 21692 13388
rect 21640 13345 21649 13379
rect 21649 13345 21683 13379
rect 21683 13345 21692 13379
rect 21640 13336 21692 13345
rect 21916 13336 21968 13388
rect 20996 13268 21048 13320
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 23940 13379 23992 13388
rect 23940 13345 23949 13379
rect 23949 13345 23983 13379
rect 23983 13345 23992 13379
rect 23940 13336 23992 13345
rect 24584 13404 24636 13456
rect 24216 13379 24268 13388
rect 24216 13345 24225 13379
rect 24225 13345 24259 13379
rect 24259 13345 24268 13379
rect 24216 13336 24268 13345
rect 25228 13404 25280 13456
rect 28632 13472 28684 13524
rect 29552 13472 29604 13524
rect 30840 13472 30892 13524
rect 27988 13404 28040 13456
rect 29460 13404 29512 13456
rect 22008 13268 22060 13320
rect 21732 13200 21784 13252
rect 24400 13268 24452 13320
rect 26056 13336 26108 13388
rect 26332 13336 26384 13388
rect 25688 13311 25740 13320
rect 25688 13277 25697 13311
rect 25697 13277 25731 13311
rect 25731 13277 25740 13311
rect 25688 13268 25740 13277
rect 26976 13336 27028 13388
rect 28172 13336 28224 13388
rect 28908 13379 28960 13388
rect 28908 13345 28917 13379
rect 28917 13345 28951 13379
rect 28951 13345 28960 13379
rect 28908 13336 28960 13345
rect 31116 13336 31168 13388
rect 30932 13268 30984 13320
rect 24952 13200 25004 13252
rect 29276 13200 29328 13252
rect 13544 13132 13596 13184
rect 14740 13175 14792 13184
rect 14740 13141 14749 13175
rect 14749 13141 14783 13175
rect 14783 13141 14792 13175
rect 14740 13132 14792 13141
rect 16672 13132 16724 13184
rect 17684 13132 17736 13184
rect 18880 13132 18932 13184
rect 19708 13132 19760 13184
rect 19800 13175 19852 13184
rect 19800 13141 19809 13175
rect 19809 13141 19843 13175
rect 19843 13141 19852 13175
rect 19800 13132 19852 13141
rect 20996 13132 21048 13184
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 22468 13132 22520 13184
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 11436 13030 11488 13082
rect 11500 13030 11552 13082
rect 11564 13030 11616 13082
rect 11628 13030 11680 13082
rect 11692 13030 11744 13082
rect 19210 13030 19262 13082
rect 19274 13030 19326 13082
rect 19338 13030 19390 13082
rect 19402 13030 19454 13082
rect 19466 13030 19518 13082
rect 26984 13030 27036 13082
rect 27048 13030 27100 13082
rect 27112 13030 27164 13082
rect 27176 13030 27228 13082
rect 27240 13030 27292 13082
rect 10416 12928 10468 12980
rect 5080 12860 5132 12912
rect 9404 12860 9456 12912
rect 10600 12860 10652 12912
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 5908 12792 5960 12844
rect 6092 12835 6144 12844
rect 6092 12801 6101 12835
rect 6101 12801 6135 12835
rect 6135 12801 6144 12835
rect 6092 12792 6144 12801
rect 2044 12724 2096 12776
rect 1860 12656 1912 12708
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 7472 12724 7524 12776
rect 7748 12724 7800 12776
rect 3516 12656 3568 12708
rect 7104 12656 7156 12708
rect 8208 12724 8260 12776
rect 9036 12724 9088 12776
rect 9772 12724 9824 12776
rect 11520 12724 11572 12776
rect 11888 12767 11940 12776
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 14556 12928 14608 12980
rect 14924 12971 14976 12980
rect 14924 12937 14933 12971
rect 14933 12937 14967 12971
rect 14967 12937 14976 12971
rect 14924 12928 14976 12937
rect 15476 12928 15528 12980
rect 16488 12928 16540 12980
rect 19064 12928 19116 12980
rect 19616 12971 19668 12980
rect 19616 12937 19625 12971
rect 19625 12937 19659 12971
rect 19659 12937 19668 12971
rect 19616 12928 19668 12937
rect 21640 12971 21692 12980
rect 21640 12937 21649 12971
rect 21649 12937 21683 12971
rect 21683 12937 21692 12971
rect 21640 12928 21692 12937
rect 29184 12928 29236 12980
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 15384 12792 15436 12844
rect 11888 12724 11940 12733
rect 14096 12724 14148 12776
rect 15844 12724 15896 12776
rect 16396 12724 16448 12776
rect 16488 12767 16540 12776
rect 16488 12733 16497 12767
rect 16497 12733 16531 12767
rect 16531 12733 16540 12767
rect 16488 12724 16540 12733
rect 16672 12724 16724 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 11060 12656 11112 12708
rect 12992 12656 13044 12708
rect 1952 12588 2004 12640
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 6920 12588 6972 12640
rect 7656 12631 7708 12640
rect 7656 12597 7665 12631
rect 7665 12597 7699 12631
rect 7699 12597 7708 12631
rect 7656 12588 7708 12597
rect 10968 12588 11020 12640
rect 12440 12588 12492 12640
rect 13452 12588 13504 12640
rect 13820 12699 13872 12708
rect 13820 12665 13854 12699
rect 13854 12665 13872 12699
rect 13820 12656 13872 12665
rect 14648 12588 14700 12640
rect 15384 12588 15436 12640
rect 18144 12656 18196 12708
rect 20076 12860 20128 12912
rect 19708 12767 19760 12776
rect 19708 12733 19717 12767
rect 19717 12733 19751 12767
rect 19751 12733 19760 12767
rect 19708 12724 19760 12733
rect 19984 12767 20036 12776
rect 19984 12733 19993 12767
rect 19993 12733 20027 12767
rect 20027 12733 20036 12767
rect 19984 12724 20036 12733
rect 19800 12656 19852 12708
rect 20536 12724 20588 12776
rect 20904 12792 20956 12844
rect 23756 12792 23808 12844
rect 24400 12792 24452 12844
rect 28448 12792 28500 12844
rect 21088 12724 21140 12776
rect 20628 12699 20680 12708
rect 20628 12665 20637 12699
rect 20637 12665 20671 12699
rect 20671 12665 20680 12699
rect 20628 12656 20680 12665
rect 21732 12724 21784 12776
rect 23112 12724 23164 12776
rect 29000 12724 29052 12776
rect 30104 12792 30156 12844
rect 28816 12656 28868 12708
rect 16672 12588 16724 12640
rect 19064 12631 19116 12640
rect 19064 12597 19073 12631
rect 19073 12597 19107 12631
rect 19107 12597 19116 12631
rect 19064 12588 19116 12597
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 21364 12588 21416 12640
rect 21640 12588 21692 12640
rect 22008 12588 22060 12640
rect 23756 12588 23808 12640
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 12096 12486 12148 12538
rect 12160 12486 12212 12538
rect 12224 12486 12276 12538
rect 12288 12486 12340 12538
rect 12352 12486 12404 12538
rect 19870 12486 19922 12538
rect 19934 12486 19986 12538
rect 19998 12486 20050 12538
rect 20062 12486 20114 12538
rect 20126 12486 20178 12538
rect 27644 12486 27696 12538
rect 27708 12486 27760 12538
rect 27772 12486 27824 12538
rect 27836 12486 27888 12538
rect 27900 12486 27952 12538
rect 1952 12291 2004 12300
rect 1952 12257 1961 12291
rect 1961 12257 1995 12291
rect 1995 12257 2004 12291
rect 1952 12248 2004 12257
rect 2780 12248 2832 12300
rect 3424 12248 3476 12300
rect 5172 12384 5224 12436
rect 6920 12384 6972 12436
rect 7748 12384 7800 12436
rect 4068 12316 4120 12368
rect 9036 12384 9088 12436
rect 9588 12384 9640 12436
rect 11060 12384 11112 12436
rect 13728 12384 13780 12436
rect 4436 12248 4488 12300
rect 6920 12291 6972 12300
rect 6920 12257 6929 12291
rect 6929 12257 6963 12291
rect 6963 12257 6972 12291
rect 6920 12248 6972 12257
rect 7104 12291 7156 12300
rect 7104 12257 7113 12291
rect 7113 12257 7147 12291
rect 7147 12257 7156 12291
rect 7104 12248 7156 12257
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 4804 12180 4856 12232
rect 7012 12155 7064 12164
rect 7012 12121 7021 12155
rect 7021 12121 7055 12155
rect 7055 12121 7064 12155
rect 7012 12112 7064 12121
rect 7104 12112 7156 12164
rect 7380 12112 7432 12164
rect 8392 12248 8444 12300
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 8668 12291 8720 12300
rect 8668 12257 8677 12291
rect 8677 12257 8711 12291
rect 8711 12257 8720 12291
rect 8668 12248 8720 12257
rect 9496 12248 9548 12300
rect 14740 12384 14792 12436
rect 18144 12384 18196 12436
rect 19064 12384 19116 12436
rect 14188 12316 14240 12368
rect 8116 12180 8168 12232
rect 8484 12044 8536 12096
rect 9496 12044 9548 12096
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 10232 12291 10284 12300
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 11152 12248 11204 12300
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 14280 12291 14332 12300
rect 14280 12257 14289 12291
rect 14289 12257 14323 12291
rect 14323 12257 14332 12291
rect 14280 12248 14332 12257
rect 11244 12112 11296 12164
rect 11888 12180 11940 12232
rect 13452 12180 13504 12232
rect 15292 12248 15344 12300
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 12440 12112 12492 12164
rect 14648 12180 14700 12232
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 17868 12316 17920 12368
rect 20996 12384 21048 12436
rect 19616 12316 19668 12368
rect 19984 12316 20036 12368
rect 21364 12316 21416 12368
rect 21824 12316 21876 12368
rect 16672 12248 16724 12300
rect 16856 12291 16908 12300
rect 16856 12257 16890 12291
rect 16890 12257 16908 12291
rect 16856 12248 16908 12257
rect 18696 12291 18748 12300
rect 18696 12257 18705 12291
rect 18705 12257 18739 12291
rect 18739 12257 18748 12291
rect 18696 12248 18748 12257
rect 18880 12291 18932 12300
rect 18880 12257 18889 12291
rect 18889 12257 18923 12291
rect 18923 12257 18932 12291
rect 18880 12248 18932 12257
rect 17960 12180 18012 12232
rect 20168 12248 20220 12300
rect 20628 12248 20680 12300
rect 22836 12291 22888 12300
rect 22836 12257 22845 12291
rect 22845 12257 22879 12291
rect 22879 12257 22888 12291
rect 22836 12248 22888 12257
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 27344 12316 27396 12368
rect 23756 12291 23808 12300
rect 23756 12257 23765 12291
rect 23765 12257 23799 12291
rect 23799 12257 23808 12291
rect 23756 12248 23808 12257
rect 28908 12248 28960 12300
rect 28816 12180 28868 12232
rect 29552 12291 29604 12300
rect 29552 12257 29561 12291
rect 29561 12257 29595 12291
rect 29595 12257 29604 12291
rect 29552 12248 29604 12257
rect 31024 12248 31076 12300
rect 30932 12223 30984 12232
rect 30932 12189 30941 12223
rect 30941 12189 30975 12223
rect 30975 12189 30984 12223
rect 30932 12180 30984 12189
rect 16488 12112 16540 12164
rect 21456 12112 21508 12164
rect 10324 12044 10376 12096
rect 10600 12044 10652 12096
rect 13912 12044 13964 12096
rect 14004 12044 14056 12096
rect 15752 12044 15804 12096
rect 16120 12044 16172 12096
rect 16396 12044 16448 12096
rect 18512 12044 18564 12096
rect 18696 12044 18748 12096
rect 20352 12044 20404 12096
rect 26424 12112 26476 12164
rect 21732 12044 21784 12096
rect 21916 12044 21968 12096
rect 23480 12087 23532 12096
rect 23480 12053 23489 12087
rect 23489 12053 23523 12087
rect 23523 12053 23532 12087
rect 23480 12044 23532 12053
rect 23572 12044 23624 12096
rect 23848 12044 23900 12096
rect 28172 12087 28224 12096
rect 28172 12053 28181 12087
rect 28181 12053 28215 12087
rect 28215 12053 28224 12087
rect 28172 12044 28224 12053
rect 29184 12044 29236 12096
rect 29736 12087 29788 12096
rect 29736 12053 29745 12087
rect 29745 12053 29779 12087
rect 29779 12053 29788 12087
rect 29736 12044 29788 12053
rect 29920 12087 29972 12096
rect 29920 12053 29929 12087
rect 29929 12053 29963 12087
rect 29963 12053 29972 12087
rect 29920 12044 29972 12053
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 11436 11942 11488 11994
rect 11500 11942 11552 11994
rect 11564 11942 11616 11994
rect 11628 11942 11680 11994
rect 11692 11942 11744 11994
rect 19210 11942 19262 11994
rect 19274 11942 19326 11994
rect 19338 11942 19390 11994
rect 19402 11942 19454 11994
rect 19466 11942 19518 11994
rect 26984 11942 27036 11994
rect 27048 11942 27100 11994
rect 27112 11942 27164 11994
rect 27176 11942 27228 11994
rect 27240 11942 27292 11994
rect 3516 11840 3568 11892
rect 7748 11840 7800 11892
rect 3424 11772 3476 11824
rect 10048 11883 10100 11892
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 12440 11840 12492 11892
rect 3884 11747 3936 11756
rect 2504 11636 2556 11688
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 13636 11772 13688 11824
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14280 11840 14332 11892
rect 15660 11840 15712 11892
rect 16856 11840 16908 11892
rect 18052 11840 18104 11892
rect 28080 11840 28132 11892
rect 28816 11883 28868 11892
rect 28816 11849 28825 11883
rect 28825 11849 28859 11883
rect 28859 11849 28868 11883
rect 28816 11840 28868 11849
rect 17960 11772 18012 11824
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 3792 11636 3844 11688
rect 3976 11636 4028 11688
rect 4160 11704 4212 11756
rect 4344 11704 4396 11756
rect 4896 11704 4948 11756
rect 6276 11704 6328 11756
rect 7380 11704 7432 11756
rect 1952 11611 2004 11620
rect 1952 11577 1986 11611
rect 1986 11577 2004 11611
rect 1952 11568 2004 11577
rect 2044 11568 2096 11620
rect 2780 11568 2832 11620
rect 3516 11611 3568 11620
rect 3516 11577 3525 11611
rect 3525 11577 3559 11611
rect 3559 11577 3568 11611
rect 3516 11568 3568 11577
rect 3608 11611 3660 11620
rect 3608 11577 3617 11611
rect 3617 11577 3651 11611
rect 3651 11577 3660 11611
rect 4436 11636 4488 11688
rect 5540 11636 5592 11688
rect 7196 11636 7248 11688
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 3608 11568 3660 11577
rect 5724 11568 5776 11620
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 8484 11636 8536 11688
rect 9956 11636 10008 11688
rect 10784 11636 10836 11688
rect 9036 11568 9088 11620
rect 10324 11568 10376 11620
rect 11796 11636 11848 11688
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 12992 11636 13044 11645
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 15200 11704 15252 11756
rect 15476 11704 15528 11756
rect 14096 11679 14148 11688
rect 14096 11645 14105 11679
rect 14105 11645 14139 11679
rect 14139 11645 14148 11679
rect 14096 11636 14148 11645
rect 4896 11500 4948 11552
rect 5816 11500 5868 11552
rect 7564 11500 7616 11552
rect 8392 11500 8444 11552
rect 9312 11500 9364 11552
rect 14004 11543 14056 11552
rect 14004 11509 14013 11543
rect 14013 11509 14047 11543
rect 14047 11509 14056 11543
rect 14004 11500 14056 11509
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 15752 11679 15804 11688
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 15936 11679 15988 11688
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 16580 11636 16632 11688
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 18604 11704 18656 11756
rect 19248 11704 19300 11756
rect 17684 11568 17736 11620
rect 18512 11636 18564 11688
rect 20628 11704 20680 11756
rect 19800 11636 19852 11688
rect 19984 11679 20036 11688
rect 19984 11645 19993 11679
rect 19993 11645 20027 11679
rect 20027 11645 20036 11679
rect 19984 11636 20036 11645
rect 20168 11679 20220 11688
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 21732 11772 21784 11824
rect 23020 11772 23072 11824
rect 23480 11772 23532 11824
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 21180 11636 21232 11645
rect 21456 11704 21508 11756
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 21548 11636 21600 11688
rect 21732 11679 21784 11688
rect 21732 11645 21741 11679
rect 21741 11645 21775 11679
rect 21775 11645 21784 11679
rect 21732 11636 21784 11645
rect 26424 11815 26476 11824
rect 26424 11781 26433 11815
rect 26433 11781 26467 11815
rect 26467 11781 26476 11815
rect 26424 11772 26476 11781
rect 23848 11747 23900 11756
rect 23848 11713 23857 11747
rect 23857 11713 23891 11747
rect 23891 11713 23900 11747
rect 23848 11704 23900 11713
rect 25320 11679 25372 11688
rect 18420 11500 18472 11552
rect 20720 11568 20772 11620
rect 23480 11611 23532 11620
rect 23480 11577 23489 11611
rect 23489 11577 23523 11611
rect 23523 11577 23532 11611
rect 23480 11568 23532 11577
rect 24216 11568 24268 11620
rect 19248 11500 19300 11552
rect 19708 11500 19760 11552
rect 19800 11543 19852 11552
rect 19800 11509 19809 11543
rect 19809 11509 19843 11543
rect 19843 11509 19852 11543
rect 19800 11500 19852 11509
rect 19892 11500 19944 11552
rect 21272 11500 21324 11552
rect 23296 11500 23348 11552
rect 25320 11645 25329 11679
rect 25329 11645 25363 11679
rect 25363 11645 25372 11679
rect 25320 11636 25372 11645
rect 25596 11636 25648 11688
rect 25780 11679 25832 11688
rect 25780 11645 25789 11679
rect 25789 11645 25823 11679
rect 25823 11645 25832 11679
rect 25780 11636 25832 11645
rect 25872 11679 25924 11688
rect 25872 11645 25882 11679
rect 25882 11645 25916 11679
rect 25916 11645 25924 11679
rect 25872 11636 25924 11645
rect 26792 11679 26844 11688
rect 26792 11645 26801 11679
rect 26801 11645 26835 11679
rect 26835 11645 26844 11679
rect 26792 11636 26844 11645
rect 26884 11679 26936 11688
rect 26884 11645 26893 11679
rect 26893 11645 26927 11679
rect 26927 11645 26936 11679
rect 26884 11636 26936 11645
rect 27344 11704 27396 11756
rect 29184 11747 29236 11756
rect 29184 11713 29193 11747
rect 29193 11713 29227 11747
rect 29227 11713 29236 11747
rect 29184 11704 29236 11713
rect 28172 11636 28224 11688
rect 29736 11636 29788 11688
rect 31116 11636 31168 11688
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 27068 11611 27120 11620
rect 27068 11577 27077 11611
rect 27077 11577 27111 11611
rect 27111 11577 27120 11611
rect 27068 11568 27120 11577
rect 27528 11568 27580 11620
rect 29092 11568 29144 11620
rect 25228 11500 25280 11509
rect 28540 11500 28592 11552
rect 30748 11500 30800 11552
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 12096 11398 12148 11450
rect 12160 11398 12212 11450
rect 12224 11398 12276 11450
rect 12288 11398 12340 11450
rect 12352 11398 12404 11450
rect 19870 11398 19922 11450
rect 19934 11398 19986 11450
rect 19998 11398 20050 11450
rect 20062 11398 20114 11450
rect 20126 11398 20178 11450
rect 27644 11398 27696 11450
rect 27708 11398 27760 11450
rect 27772 11398 27824 11450
rect 27836 11398 27888 11450
rect 27900 11398 27952 11450
rect 3516 11296 3568 11348
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 2596 11203 2648 11212
rect 2596 11169 2630 11203
rect 2630 11169 2648 11203
rect 2596 11160 2648 11169
rect 5172 11296 5224 11348
rect 6552 11296 6604 11348
rect 5908 11228 5960 11280
rect 6092 11271 6144 11280
rect 6092 11237 6126 11271
rect 6126 11237 6144 11271
rect 6092 11228 6144 11237
rect 6184 11228 6236 11280
rect 7564 11296 7616 11348
rect 7656 11228 7708 11280
rect 8576 11296 8628 11348
rect 13636 11296 13688 11348
rect 19616 11296 19668 11348
rect 19800 11296 19852 11348
rect 20536 11296 20588 11348
rect 21732 11296 21784 11348
rect 23480 11296 23532 11348
rect 25228 11296 25280 11348
rect 25780 11296 25832 11348
rect 26792 11296 26844 11348
rect 28816 11296 28868 11348
rect 5356 11203 5408 11212
rect 5356 11169 5365 11203
rect 5365 11169 5399 11203
rect 5399 11169 5408 11203
rect 5356 11160 5408 11169
rect 5724 11160 5776 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 5264 11092 5316 11144
rect 8300 11160 8352 11212
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 8760 11203 8812 11212
rect 8760 11169 8769 11203
rect 8769 11169 8803 11203
rect 8803 11169 8812 11203
rect 8760 11160 8812 11169
rect 9956 11271 10008 11280
rect 9956 11237 9965 11271
rect 9965 11237 9999 11271
rect 9999 11237 10008 11271
rect 9956 11228 10008 11237
rect 10048 11228 10100 11280
rect 9312 11203 9364 11212
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 9312 11160 9364 11169
rect 9864 11160 9916 11212
rect 10600 11203 10652 11212
rect 10600 11169 10609 11203
rect 10609 11169 10643 11203
rect 10643 11169 10652 11203
rect 10600 11160 10652 11169
rect 11060 11228 11112 11280
rect 15384 11160 15436 11212
rect 15844 11203 15896 11212
rect 15844 11169 15853 11203
rect 15853 11169 15887 11203
rect 15887 11169 15896 11203
rect 15844 11160 15896 11169
rect 16120 11203 16172 11212
rect 16120 11169 16129 11203
rect 16129 11169 16163 11203
rect 16163 11169 16172 11203
rect 16120 11160 16172 11169
rect 20352 11228 20404 11280
rect 21180 11228 21232 11280
rect 8484 11024 8536 11076
rect 9036 11024 9088 11076
rect 10324 11067 10376 11076
rect 10324 11033 10333 11067
rect 10333 11033 10367 11067
rect 10367 11033 10376 11067
rect 10324 11024 10376 11033
rect 5264 10956 5316 11008
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 8944 10956 8996 11008
rect 10416 10956 10468 11008
rect 12716 11092 12768 11144
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 18236 11092 18288 11144
rect 11888 11024 11940 11076
rect 12808 11024 12860 11076
rect 13176 11024 13228 11076
rect 13544 11024 13596 11076
rect 16028 11024 16080 11076
rect 18788 11024 18840 11076
rect 20260 11092 20312 11144
rect 19708 11024 19760 11076
rect 22008 11203 22060 11212
rect 22008 11169 22017 11203
rect 22017 11169 22051 11203
rect 22051 11169 22060 11203
rect 22008 11160 22060 11169
rect 24216 11228 24268 11280
rect 25596 11228 25648 11280
rect 22100 11092 22152 11144
rect 23296 11203 23348 11212
rect 23296 11169 23305 11203
rect 23305 11169 23339 11203
rect 23339 11169 23348 11203
rect 23296 11160 23348 11169
rect 23572 11160 23624 11212
rect 23756 11203 23808 11212
rect 23756 11169 23790 11203
rect 23790 11169 23808 11203
rect 23756 11160 23808 11169
rect 28172 11160 28224 11212
rect 28908 11160 28960 11212
rect 29092 11203 29144 11212
rect 29092 11169 29101 11203
rect 29101 11169 29135 11203
rect 29135 11169 29144 11203
rect 29092 11160 29144 11169
rect 25320 11024 25372 11076
rect 27620 11024 27672 11076
rect 11336 10956 11388 11008
rect 12992 10956 13044 11008
rect 16764 10956 16816 11008
rect 21732 10956 21784 11008
rect 24860 10999 24912 11008
rect 24860 10965 24869 10999
rect 24869 10965 24903 10999
rect 24903 10965 24912 10999
rect 24860 10956 24912 10965
rect 26148 10956 26200 11008
rect 31116 11296 31168 11348
rect 29920 11228 29972 11280
rect 30012 11160 30064 11212
rect 30748 11203 30800 11212
rect 30748 11169 30757 11203
rect 30757 11169 30791 11203
rect 30791 11169 30800 11203
rect 30748 11160 30800 11169
rect 29552 11024 29604 11076
rect 28540 10999 28592 11008
rect 28540 10965 28549 10999
rect 28549 10965 28583 10999
rect 28583 10965 28592 10999
rect 28540 10956 28592 10965
rect 29000 10999 29052 11008
rect 29000 10965 29009 10999
rect 29009 10965 29043 10999
rect 29043 10965 29052 10999
rect 29000 10956 29052 10965
rect 31300 10999 31352 11008
rect 31300 10965 31309 10999
rect 31309 10965 31343 10999
rect 31343 10965 31352 10999
rect 31300 10956 31352 10965
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 11436 10854 11488 10906
rect 11500 10854 11552 10906
rect 11564 10854 11616 10906
rect 11628 10854 11680 10906
rect 11692 10854 11744 10906
rect 19210 10854 19262 10906
rect 19274 10854 19326 10906
rect 19338 10854 19390 10906
rect 19402 10854 19454 10906
rect 19466 10854 19518 10906
rect 26984 10854 27036 10906
rect 27048 10854 27100 10906
rect 27112 10854 27164 10906
rect 27176 10854 27228 10906
rect 27240 10854 27292 10906
rect 2596 10752 2648 10804
rect 3056 10752 3108 10804
rect 5172 10752 5224 10804
rect 6092 10752 6144 10804
rect 6736 10752 6788 10804
rect 8760 10795 8812 10804
rect 8760 10761 8769 10795
rect 8769 10761 8803 10795
rect 8803 10761 8812 10795
rect 8760 10752 8812 10761
rect 12624 10752 12676 10804
rect 15844 10795 15896 10804
rect 15844 10761 15853 10795
rect 15853 10761 15887 10795
rect 15887 10761 15896 10795
rect 15844 10752 15896 10761
rect 18236 10752 18288 10804
rect 20444 10752 20496 10804
rect 20720 10752 20772 10804
rect 22100 10795 22152 10804
rect 22100 10761 22109 10795
rect 22109 10761 22143 10795
rect 22143 10761 22152 10795
rect 22100 10752 22152 10761
rect 23756 10752 23808 10804
rect 25872 10795 25924 10804
rect 25872 10761 25881 10795
rect 25881 10761 25915 10795
rect 25915 10761 25924 10795
rect 25872 10752 25924 10761
rect 30012 10752 30064 10804
rect 7196 10727 7248 10736
rect 7196 10693 7205 10727
rect 7205 10693 7239 10727
rect 7239 10693 7248 10727
rect 7196 10684 7248 10693
rect 8852 10684 8904 10736
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 2044 10548 2096 10600
rect 2780 10548 2832 10600
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 8944 10616 8996 10668
rect 4160 10480 4212 10532
rect 4804 10480 4856 10532
rect 5908 10480 5960 10532
rect 6276 10480 6328 10532
rect 6460 10480 6512 10532
rect 8024 10548 8076 10600
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 10232 10591 10284 10600
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 11796 10548 11848 10600
rect 12164 10548 12216 10600
rect 18696 10684 18748 10736
rect 15384 10659 15436 10668
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 15936 10616 15988 10668
rect 12532 10591 12584 10600
rect 12532 10557 12541 10591
rect 12541 10557 12575 10591
rect 12575 10557 12584 10591
rect 12532 10548 12584 10557
rect 12808 10591 12860 10600
rect 12808 10557 12843 10591
rect 12843 10557 12860 10591
rect 12808 10548 12860 10557
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 1952 10412 2004 10464
rect 5540 10412 5592 10464
rect 11980 10480 12032 10532
rect 12440 10480 12492 10532
rect 12716 10523 12768 10532
rect 12716 10489 12725 10523
rect 12725 10489 12759 10523
rect 12759 10489 12768 10523
rect 12716 10480 12768 10489
rect 14004 10548 14056 10600
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 9772 10412 9824 10464
rect 10048 10412 10100 10464
rect 10416 10412 10468 10464
rect 11704 10412 11756 10464
rect 12164 10412 12216 10464
rect 13728 10480 13780 10532
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15200 10548 15252 10557
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 16396 10616 16448 10668
rect 16488 10659 16540 10668
rect 16488 10625 16497 10659
rect 16497 10625 16531 10659
rect 16531 10625 16540 10659
rect 16488 10616 16540 10625
rect 16764 10591 16816 10600
rect 16764 10557 16773 10591
rect 16773 10557 16807 10591
rect 16807 10557 16816 10591
rect 16764 10548 16816 10557
rect 18236 10591 18288 10600
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 14556 10412 14608 10464
rect 15016 10455 15068 10464
rect 15016 10421 15025 10455
rect 15025 10421 15059 10455
rect 15059 10421 15068 10455
rect 15016 10412 15068 10421
rect 16304 10523 16356 10532
rect 16304 10489 16339 10523
rect 16339 10489 16356 10523
rect 16304 10480 16356 10489
rect 18328 10480 18380 10532
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 18788 10548 18840 10600
rect 20444 10591 20496 10600
rect 20444 10557 20453 10591
rect 20453 10557 20487 10591
rect 20487 10557 20496 10591
rect 20444 10548 20496 10557
rect 22836 10548 22888 10600
rect 19064 10480 19116 10532
rect 21272 10480 21324 10532
rect 21456 10480 21508 10532
rect 22008 10480 22060 10532
rect 23112 10591 23164 10600
rect 23112 10557 23121 10591
rect 23121 10557 23155 10591
rect 23155 10557 23164 10591
rect 23112 10548 23164 10557
rect 24860 10548 24912 10600
rect 24216 10523 24268 10532
rect 24216 10489 24225 10523
rect 24225 10489 24259 10523
rect 24259 10489 24268 10523
rect 24216 10480 24268 10489
rect 16764 10412 16816 10464
rect 17960 10412 18012 10464
rect 18972 10412 19024 10464
rect 20260 10412 20312 10464
rect 25872 10616 25924 10668
rect 29552 10684 29604 10736
rect 30932 10752 30984 10804
rect 29000 10616 29052 10668
rect 26148 10548 26200 10600
rect 26332 10591 26384 10600
rect 26332 10557 26341 10591
rect 26341 10557 26375 10591
rect 26375 10557 26384 10591
rect 26332 10548 26384 10557
rect 28908 10548 28960 10600
rect 30104 10659 30156 10668
rect 30104 10625 30113 10659
rect 30113 10625 30147 10659
rect 30147 10625 30156 10659
rect 30104 10616 30156 10625
rect 31116 10548 31168 10600
rect 31300 10548 31352 10600
rect 30748 10480 30800 10532
rect 28632 10412 28684 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 12096 10310 12148 10362
rect 12160 10310 12212 10362
rect 12224 10310 12276 10362
rect 12288 10310 12340 10362
rect 12352 10310 12404 10362
rect 19870 10310 19922 10362
rect 19934 10310 19986 10362
rect 19998 10310 20050 10362
rect 20062 10310 20114 10362
rect 20126 10310 20178 10362
rect 27644 10310 27696 10362
rect 27708 10310 27760 10362
rect 27772 10310 27824 10362
rect 27836 10310 27888 10362
rect 27900 10310 27952 10362
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 2044 10140 2096 10192
rect 3516 10140 3568 10192
rect 4436 10140 4488 10192
rect 4712 10140 4764 10192
rect 5356 10140 5408 10192
rect 6460 10140 6512 10192
rect 7196 10208 7248 10260
rect 9312 10208 9364 10260
rect 6828 10183 6880 10192
rect 6828 10149 6863 10183
rect 6863 10149 6880 10183
rect 6828 10140 6880 10149
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 1584 10004 1636 10056
rect 2964 10072 3016 10124
rect 3700 10115 3752 10124
rect 3700 10081 3709 10115
rect 3709 10081 3743 10115
rect 3743 10081 3752 10115
rect 3700 10072 3752 10081
rect 3792 10115 3844 10124
rect 3792 10081 3801 10115
rect 3801 10081 3835 10115
rect 3835 10081 3844 10115
rect 3792 10072 3844 10081
rect 4252 10072 4304 10124
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 7748 10140 7800 10192
rect 8668 10140 8720 10192
rect 7288 10072 7340 10124
rect 8392 10072 8444 10124
rect 9772 10115 9824 10124
rect 9772 10081 9790 10115
rect 9790 10081 9824 10115
rect 9772 10072 9824 10081
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 4344 10004 4396 10056
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 3792 9936 3844 9988
rect 10968 10140 11020 10192
rect 12072 10140 12124 10192
rect 13544 10208 13596 10260
rect 13636 10208 13688 10260
rect 14004 10251 14056 10260
rect 14004 10217 14013 10251
rect 14013 10217 14047 10251
rect 14047 10217 14056 10251
rect 14004 10208 14056 10217
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11704 10072 11756 10124
rect 12440 10140 12492 10192
rect 11336 10004 11388 10056
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 3240 9868 3292 9920
rect 3516 9868 3568 9920
rect 3700 9868 3752 9920
rect 5724 9868 5776 9920
rect 6828 9868 6880 9920
rect 8484 9868 8536 9920
rect 8760 9868 8812 9920
rect 10784 9868 10836 9920
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 12624 10115 12676 10124
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 15016 10140 15068 10192
rect 18420 10208 18472 10260
rect 18696 10208 18748 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 18328 10140 18380 10192
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 16028 10072 16080 10124
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 18052 10115 18104 10124
rect 18052 10081 18061 10115
rect 18061 10081 18095 10115
rect 18095 10081 18104 10115
rect 18052 10072 18104 10081
rect 18880 10072 18932 10124
rect 20444 10140 20496 10192
rect 21548 10115 21600 10124
rect 21548 10081 21557 10115
rect 21557 10081 21591 10115
rect 21591 10081 21600 10115
rect 21548 10072 21600 10081
rect 21364 10004 21416 10056
rect 21732 10115 21784 10124
rect 21732 10081 21741 10115
rect 21741 10081 21775 10115
rect 21775 10081 21784 10115
rect 21732 10072 21784 10081
rect 21916 10115 21968 10124
rect 21916 10081 21925 10115
rect 21925 10081 21959 10115
rect 21959 10081 21968 10115
rect 21916 10072 21968 10081
rect 22376 10140 22428 10192
rect 24216 10140 24268 10192
rect 24860 10140 24912 10192
rect 25872 10208 25924 10260
rect 26332 10208 26384 10260
rect 30104 10208 30156 10260
rect 30288 10208 30340 10260
rect 23480 10072 23532 10124
rect 25044 10072 25096 10124
rect 22008 10004 22060 10056
rect 12440 9868 12492 9920
rect 15476 9868 15528 9920
rect 16212 9868 16264 9920
rect 16856 9868 16908 9920
rect 22100 9868 22152 9920
rect 22928 9868 22980 9920
rect 25136 9868 25188 9920
rect 25780 10115 25832 10124
rect 25780 10081 25789 10115
rect 25789 10081 25823 10115
rect 25823 10081 25832 10115
rect 25780 10072 25832 10081
rect 25872 10115 25924 10124
rect 25872 10081 25881 10115
rect 25881 10081 25915 10115
rect 25915 10081 25924 10115
rect 25872 10072 25924 10081
rect 26792 10072 26844 10124
rect 28632 10115 28684 10124
rect 28632 10081 28641 10115
rect 28641 10081 28675 10115
rect 28675 10081 28684 10115
rect 28632 10072 28684 10081
rect 28816 10115 28868 10124
rect 28816 10081 28825 10115
rect 28825 10081 28859 10115
rect 28859 10081 28868 10115
rect 28816 10072 28868 10081
rect 30196 10072 30248 10124
rect 31024 10115 31076 10124
rect 31024 10081 31033 10115
rect 31033 10081 31067 10115
rect 31067 10081 31076 10115
rect 31024 10072 31076 10081
rect 28908 10047 28960 10056
rect 26332 9936 26384 9988
rect 28908 10013 28917 10047
rect 28917 10013 28951 10047
rect 28951 10013 28960 10047
rect 28908 10004 28960 10013
rect 30104 9868 30156 9920
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 11436 9766 11488 9818
rect 11500 9766 11552 9818
rect 11564 9766 11616 9818
rect 11628 9766 11680 9818
rect 11692 9766 11744 9818
rect 19210 9766 19262 9818
rect 19274 9766 19326 9818
rect 19338 9766 19390 9818
rect 19402 9766 19454 9818
rect 19466 9766 19518 9818
rect 26984 9766 27036 9818
rect 27048 9766 27100 9818
rect 27112 9766 27164 9818
rect 27176 9766 27228 9818
rect 27240 9766 27292 9818
rect 1584 9707 1636 9716
rect 1584 9673 1593 9707
rect 1593 9673 1627 9707
rect 1627 9673 1636 9707
rect 1584 9664 1636 9673
rect 2044 9664 2096 9716
rect 2964 9664 3016 9716
rect 3746 9664 3798 9716
rect 3976 9664 4028 9716
rect 4436 9664 4488 9716
rect 4896 9664 4948 9716
rect 7196 9664 7248 9716
rect 8300 9664 8352 9716
rect 10140 9664 10192 9716
rect 11244 9664 11296 9716
rect 12348 9664 12400 9716
rect 12716 9664 12768 9716
rect 15200 9664 15252 9716
rect 3516 9596 3568 9648
rect 5172 9596 5224 9648
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 4896 9528 4948 9580
rect 5540 9596 5592 9648
rect 8852 9596 8904 9648
rect 2872 9460 2924 9512
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 4344 9503 4396 9512
rect 4344 9469 4353 9503
rect 4353 9469 4387 9503
rect 4387 9469 4396 9503
rect 4344 9460 4396 9469
rect 7012 9528 7064 9580
rect 7748 9528 7800 9580
rect 8576 9528 8628 9580
rect 9680 9596 9732 9648
rect 2320 9392 2372 9444
rect 3148 9392 3200 9444
rect 3516 9435 3568 9444
rect 3516 9401 3525 9435
rect 3525 9401 3559 9435
rect 3559 9401 3568 9435
rect 3516 9392 3568 9401
rect 4252 9392 4304 9444
rect 7012 9392 7064 9444
rect 2964 9324 3016 9376
rect 3240 9324 3292 9376
rect 6368 9324 6420 9376
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9312 9460 9364 9512
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 10784 9503 10836 9512
rect 10784 9469 10818 9503
rect 10818 9469 10836 9503
rect 10784 9460 10836 9469
rect 11980 9503 12032 9512
rect 11980 9469 11989 9503
rect 11989 9469 12023 9503
rect 12023 9469 12032 9503
rect 11980 9460 12032 9469
rect 12072 9460 12124 9512
rect 14280 9528 14332 9580
rect 16672 9596 16724 9648
rect 21916 9664 21968 9716
rect 25136 9707 25188 9716
rect 25136 9673 25145 9707
rect 25145 9673 25179 9707
rect 25179 9673 25188 9707
rect 25136 9664 25188 9673
rect 25780 9664 25832 9716
rect 8484 9392 8536 9444
rect 8944 9392 8996 9444
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8392 9324 8444 9376
rect 11796 9392 11848 9444
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 16212 9503 16264 9512
rect 16212 9469 16221 9503
rect 16221 9469 16255 9503
rect 16255 9469 16264 9503
rect 16212 9460 16264 9469
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 18420 9528 18472 9580
rect 23480 9639 23532 9648
rect 23480 9605 23489 9639
rect 23489 9605 23523 9639
rect 23523 9605 23532 9639
rect 23480 9596 23532 9605
rect 18696 9460 18748 9512
rect 18880 9503 18932 9512
rect 18880 9469 18889 9503
rect 18889 9469 18923 9503
rect 18923 9469 18932 9503
rect 18880 9460 18932 9469
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 14372 9392 14424 9444
rect 15936 9392 15988 9444
rect 16396 9435 16448 9444
rect 16396 9401 16431 9435
rect 16431 9401 16448 9435
rect 16396 9392 16448 9401
rect 17500 9392 17552 9444
rect 20352 9460 20404 9512
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 22100 9571 22152 9580
rect 22100 9537 22109 9571
rect 22109 9537 22143 9571
rect 22143 9537 22152 9571
rect 22100 9528 22152 9537
rect 23112 9528 23164 9580
rect 26700 9664 26752 9716
rect 28172 9664 28224 9716
rect 25964 9596 26016 9648
rect 26608 9596 26660 9648
rect 26884 9596 26936 9648
rect 27068 9596 27120 9648
rect 28080 9596 28132 9648
rect 29000 9596 29052 9648
rect 22008 9460 22060 9512
rect 21088 9392 21140 9444
rect 22468 9392 22520 9444
rect 24860 9460 24912 9512
rect 24492 9392 24544 9444
rect 25044 9503 25096 9512
rect 25044 9469 25053 9503
rect 25053 9469 25087 9503
rect 25087 9469 25096 9503
rect 25044 9460 25096 9469
rect 25228 9460 25280 9512
rect 25412 9503 25464 9512
rect 25412 9469 25421 9503
rect 25421 9469 25455 9503
rect 25455 9469 25464 9503
rect 25412 9460 25464 9469
rect 26332 9528 26384 9580
rect 27344 9528 27396 9580
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 26700 9503 26752 9512
rect 26700 9469 26709 9503
rect 26709 9469 26743 9503
rect 26743 9469 26752 9503
rect 26700 9460 26752 9469
rect 26884 9460 26936 9512
rect 26148 9392 26200 9444
rect 26240 9435 26292 9444
rect 26240 9401 26249 9435
rect 26249 9401 26283 9435
rect 26283 9401 26292 9435
rect 26240 9392 26292 9401
rect 27068 9392 27120 9444
rect 10048 9324 10100 9376
rect 11612 9324 11664 9376
rect 13544 9324 13596 9376
rect 14832 9324 14884 9376
rect 15844 9367 15896 9376
rect 15844 9333 15853 9367
rect 15853 9333 15887 9367
rect 15887 9333 15896 9367
rect 15844 9324 15896 9333
rect 17960 9324 18012 9376
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 20076 9324 20128 9376
rect 21272 9324 21324 9376
rect 22284 9324 22336 9376
rect 24952 9324 25004 9376
rect 25964 9367 26016 9376
rect 25964 9333 25973 9367
rect 25973 9333 26007 9367
rect 26007 9333 26016 9367
rect 25964 9324 26016 9333
rect 26424 9324 26476 9376
rect 26608 9324 26660 9376
rect 28080 9503 28132 9512
rect 28080 9469 28089 9503
rect 28089 9469 28123 9503
rect 28123 9469 28132 9503
rect 28080 9460 28132 9469
rect 28172 9503 28224 9512
rect 28172 9469 28181 9503
rect 28181 9469 28215 9503
rect 28215 9469 28224 9503
rect 28172 9460 28224 9469
rect 30196 9571 30248 9580
rect 30196 9537 30205 9571
rect 30205 9537 30239 9571
rect 30239 9537 30248 9571
rect 30196 9528 30248 9537
rect 28448 9435 28500 9444
rect 28448 9401 28457 9435
rect 28457 9401 28491 9435
rect 28491 9401 28500 9435
rect 28448 9392 28500 9401
rect 29920 9503 29972 9512
rect 29920 9469 29929 9503
rect 29929 9469 29963 9503
rect 29963 9469 29972 9503
rect 29920 9460 29972 9469
rect 30104 9503 30156 9512
rect 30104 9469 30113 9503
rect 30113 9469 30147 9503
rect 30147 9469 30156 9503
rect 30104 9460 30156 9469
rect 30288 9503 30340 9512
rect 30288 9469 30297 9503
rect 30297 9469 30331 9503
rect 30331 9469 30340 9503
rect 30288 9460 30340 9469
rect 28080 9324 28132 9376
rect 28816 9367 28868 9376
rect 28816 9333 28825 9367
rect 28825 9333 28859 9367
rect 28859 9333 28868 9367
rect 28816 9324 28868 9333
rect 29092 9367 29144 9376
rect 29092 9333 29101 9367
rect 29101 9333 29135 9367
rect 29135 9333 29144 9367
rect 29092 9324 29144 9333
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 12096 9222 12148 9274
rect 12160 9222 12212 9274
rect 12224 9222 12276 9274
rect 12288 9222 12340 9274
rect 12352 9222 12404 9274
rect 19870 9222 19922 9274
rect 19934 9222 19986 9274
rect 19998 9222 20050 9274
rect 20062 9222 20114 9274
rect 20126 9222 20178 9274
rect 27644 9222 27696 9274
rect 27708 9222 27760 9274
rect 27772 9222 27824 9274
rect 27836 9222 27888 9274
rect 27900 9222 27952 9274
rect 1676 9120 1728 9172
rect 2964 9120 3016 9172
rect 2044 9052 2096 9104
rect 3056 9052 3108 9104
rect 3332 9052 3384 9104
rect 3976 9052 4028 9104
rect 6828 9120 6880 9172
rect 7012 9163 7064 9172
rect 7012 9129 7021 9163
rect 7021 9129 7055 9163
rect 7055 9129 7064 9163
rect 7012 9120 7064 9129
rect 4896 9095 4948 9104
rect 4896 9061 4905 9095
rect 4905 9061 4939 9095
rect 4939 9061 4948 9095
rect 4896 9052 4948 9061
rect 7840 9120 7892 9172
rect 7564 9052 7616 9104
rect 3240 8984 3292 9036
rect 3516 8984 3568 9036
rect 3700 9027 3752 9036
rect 3700 8993 3709 9027
rect 3709 8993 3743 9027
rect 3743 8993 3752 9027
rect 3700 8984 3752 8993
rect 1768 8916 1820 8968
rect 3332 8916 3384 8968
rect 3608 8916 3660 8968
rect 4160 9027 4212 9036
rect 4160 8993 4169 9027
rect 4169 8993 4203 9027
rect 4203 8993 4212 9027
rect 4160 8984 4212 8993
rect 4988 8916 5040 8968
rect 4620 8848 4672 8900
rect 4252 8780 4304 8832
rect 4712 8780 4764 8832
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 7748 8984 7800 9036
rect 9312 9027 9364 9036
rect 9312 8993 9321 9027
rect 9321 8993 9355 9027
rect 9355 8993 9364 9027
rect 9312 8984 9364 8993
rect 9680 8984 9732 9036
rect 8668 8848 8720 8900
rect 9772 8780 9824 8832
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 11060 9120 11112 9172
rect 11980 9120 12032 9172
rect 11612 9095 11664 9104
rect 9956 8959 10008 8968
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 11244 8984 11296 9036
rect 11612 9061 11621 9095
rect 11621 9061 11655 9095
rect 11655 9061 11664 9095
rect 11612 9052 11664 9061
rect 11888 9052 11940 9104
rect 13084 9120 13136 9172
rect 14464 9120 14516 9172
rect 11152 8916 11204 8968
rect 11704 9027 11756 9036
rect 11704 8993 11713 9027
rect 11713 8993 11747 9027
rect 11747 8993 11756 9027
rect 11704 8984 11756 8993
rect 14372 9095 14424 9104
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 12072 8984 12124 9036
rect 13728 9027 13780 9036
rect 13728 8993 13737 9027
rect 13737 8993 13771 9027
rect 13771 8993 13780 9027
rect 13728 8984 13780 8993
rect 12532 8916 12584 8968
rect 14648 8984 14700 9036
rect 16120 9120 16172 9172
rect 17132 9120 17184 9172
rect 14832 9095 14884 9104
rect 14832 9061 14841 9095
rect 14841 9061 14875 9095
rect 14875 9061 14884 9095
rect 14832 9052 14884 9061
rect 16396 9052 16448 9104
rect 15200 9027 15252 9036
rect 15200 8993 15209 9027
rect 15209 8993 15243 9027
rect 15243 8993 15252 9027
rect 15200 8984 15252 8993
rect 15476 8984 15528 9036
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 18880 9120 18932 9172
rect 20628 9120 20680 9172
rect 21272 9163 21324 9172
rect 21272 9129 21281 9163
rect 21281 9129 21315 9163
rect 21315 9129 21324 9163
rect 21272 9120 21324 9129
rect 18788 9052 18840 9104
rect 20352 9052 20404 9104
rect 21088 9052 21140 9104
rect 18236 9027 18288 9036
rect 18236 8993 18270 9027
rect 18270 8993 18288 9027
rect 18236 8984 18288 8993
rect 20444 8984 20496 9036
rect 22376 9120 22428 9172
rect 22468 9163 22520 9172
rect 22468 9129 22477 9163
rect 22477 9129 22511 9163
rect 22511 9129 22520 9163
rect 22468 9120 22520 9129
rect 21916 9052 21968 9104
rect 22100 8984 22152 9036
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 22928 9027 22980 9036
rect 22928 8993 22937 9027
rect 22937 8993 22971 9027
rect 22971 8993 22980 9027
rect 22928 8984 22980 8993
rect 12716 8848 12768 8900
rect 15936 8916 15988 8968
rect 22284 8916 22336 8968
rect 15384 8848 15436 8900
rect 16028 8848 16080 8900
rect 22008 8848 22060 8900
rect 22836 8848 22888 8900
rect 10600 8780 10652 8832
rect 11152 8780 11204 8832
rect 11704 8780 11756 8832
rect 15476 8780 15528 8832
rect 18144 8780 18196 8832
rect 18972 8780 19024 8832
rect 20260 8780 20312 8832
rect 24492 8984 24544 9036
rect 24952 9095 25004 9104
rect 24952 9061 24961 9095
rect 24961 9061 24995 9095
rect 24995 9061 25004 9095
rect 24952 9052 25004 9061
rect 25872 9120 25924 9172
rect 25964 9052 26016 9104
rect 26240 9095 26292 9104
rect 26240 9061 26249 9095
rect 26249 9061 26283 9095
rect 26283 9061 26292 9095
rect 26240 9052 26292 9061
rect 26700 9120 26752 9172
rect 28448 9120 28500 9172
rect 29920 9120 29972 9172
rect 26516 9052 26568 9104
rect 29092 9052 29144 9104
rect 24584 8916 24636 8968
rect 25412 8984 25464 9036
rect 26332 8984 26384 9036
rect 28172 8984 28224 9036
rect 30012 9027 30064 9036
rect 30012 8993 30030 9027
rect 30030 8993 30064 9027
rect 30012 8984 30064 8993
rect 25228 8848 25280 8900
rect 26424 8848 26476 8900
rect 24032 8780 24084 8832
rect 25596 8823 25648 8832
rect 25596 8789 25605 8823
rect 25605 8789 25639 8823
rect 25639 8789 25648 8823
rect 25596 8780 25648 8789
rect 25780 8823 25832 8832
rect 25780 8789 25789 8823
rect 25789 8789 25823 8823
rect 25823 8789 25832 8823
rect 25780 8780 25832 8789
rect 26792 8780 26844 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 11436 8678 11488 8730
rect 11500 8678 11552 8730
rect 11564 8678 11616 8730
rect 11628 8678 11680 8730
rect 11692 8678 11744 8730
rect 19210 8678 19262 8730
rect 19274 8678 19326 8730
rect 19338 8678 19390 8730
rect 19402 8678 19454 8730
rect 19466 8678 19518 8730
rect 26984 8678 27036 8730
rect 27048 8678 27100 8730
rect 27112 8678 27164 8730
rect 27176 8678 27228 8730
rect 27240 8678 27292 8730
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 9312 8576 9364 8628
rect 9772 8576 9824 8628
rect 11612 8576 11664 8628
rect 14556 8576 14608 8628
rect 18236 8576 18288 8628
rect 3424 8440 3476 8492
rect 7288 8508 7340 8560
rect 2872 8372 2924 8424
rect 3056 8372 3108 8424
rect 4252 8372 4304 8424
rect 5172 8372 5224 8424
rect 4988 8304 5040 8356
rect 6276 8415 6328 8424
rect 6276 8381 6285 8415
rect 6285 8381 6319 8415
rect 6319 8381 6328 8415
rect 6276 8372 6328 8381
rect 6920 8440 6972 8492
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 7472 8440 7524 8492
rect 15476 8508 15528 8560
rect 15936 8508 15988 8560
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 8760 8372 8812 8424
rect 9956 8372 10008 8424
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 16212 8372 16264 8424
rect 18420 8415 18472 8424
rect 18420 8381 18429 8415
rect 18429 8381 18463 8415
rect 18463 8381 18472 8415
rect 18420 8372 18472 8381
rect 18880 8415 18932 8424
rect 18880 8381 18889 8415
rect 18889 8381 18923 8415
rect 18923 8381 18932 8415
rect 18880 8372 18932 8381
rect 21548 8440 21600 8492
rect 19156 8415 19208 8424
rect 19156 8381 19191 8415
rect 19191 8381 19208 8415
rect 19156 8372 19208 8381
rect 9588 8304 9640 8356
rect 10600 8304 10652 8356
rect 16672 8304 16724 8356
rect 18972 8347 19024 8356
rect 18972 8313 18981 8347
rect 18981 8313 19015 8347
rect 19015 8313 19024 8347
rect 18972 8304 19024 8313
rect 4896 8236 4948 8288
rect 8484 8236 8536 8288
rect 8576 8236 8628 8288
rect 10968 8236 11020 8288
rect 14832 8236 14884 8288
rect 15292 8236 15344 8288
rect 18788 8236 18840 8288
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 20444 8372 20496 8424
rect 23112 8576 23164 8628
rect 23204 8576 23256 8628
rect 22836 8440 22888 8492
rect 22652 8415 22704 8424
rect 22652 8381 22661 8415
rect 22661 8381 22695 8415
rect 22695 8381 22704 8415
rect 22652 8372 22704 8381
rect 23112 8372 23164 8424
rect 23204 8415 23256 8424
rect 23204 8381 23213 8415
rect 23213 8381 23247 8415
rect 23247 8381 23256 8415
rect 23204 8372 23256 8381
rect 24308 8440 24360 8492
rect 24492 8619 24544 8628
rect 24492 8585 24501 8619
rect 24501 8585 24535 8619
rect 24535 8585 24544 8619
rect 24492 8576 24544 8585
rect 26148 8576 26200 8628
rect 28172 8576 28224 8628
rect 30012 8576 30064 8628
rect 24584 8551 24636 8560
rect 24584 8517 24593 8551
rect 24593 8517 24627 8551
rect 24627 8517 24636 8551
rect 24584 8508 24636 8517
rect 25596 8440 25648 8492
rect 29000 8483 29052 8492
rect 29000 8449 29009 8483
rect 29009 8449 29043 8483
rect 29043 8449 29052 8483
rect 29000 8440 29052 8449
rect 23388 8415 23440 8424
rect 23388 8381 23397 8415
rect 23397 8381 23431 8415
rect 23431 8381 23440 8415
rect 23388 8372 23440 8381
rect 22744 8304 22796 8356
rect 26332 8372 26384 8424
rect 27344 8372 27396 8424
rect 27988 8372 28040 8424
rect 28816 8372 28868 8424
rect 24032 8347 24084 8356
rect 24032 8313 24041 8347
rect 24041 8313 24075 8347
rect 24075 8313 24084 8347
rect 24032 8304 24084 8313
rect 24216 8347 24268 8356
rect 24216 8313 24225 8347
rect 24225 8313 24259 8347
rect 24259 8313 24268 8347
rect 24216 8304 24268 8313
rect 24860 8304 24912 8356
rect 19800 8279 19852 8288
rect 19800 8245 19809 8279
rect 19809 8245 19843 8279
rect 19843 8245 19852 8279
rect 19800 8236 19852 8245
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 22100 8279 22152 8288
rect 22100 8245 22109 8279
rect 22109 8245 22143 8279
rect 22143 8245 22152 8279
rect 22100 8236 22152 8245
rect 23020 8236 23072 8288
rect 25228 8347 25280 8356
rect 25228 8313 25237 8347
rect 25237 8313 25271 8347
rect 25271 8313 25280 8347
rect 25228 8304 25280 8313
rect 25780 8304 25832 8356
rect 27528 8304 27580 8356
rect 25596 8279 25648 8288
rect 25596 8245 25605 8279
rect 25605 8245 25639 8279
rect 25639 8245 25648 8279
rect 25596 8236 25648 8245
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 12096 8134 12148 8186
rect 12160 8134 12212 8186
rect 12224 8134 12276 8186
rect 12288 8134 12340 8186
rect 12352 8134 12404 8186
rect 19870 8134 19922 8186
rect 19934 8134 19986 8186
rect 19998 8134 20050 8186
rect 20062 8134 20114 8186
rect 20126 8134 20178 8186
rect 27644 8134 27696 8186
rect 27708 8134 27760 8186
rect 27772 8134 27824 8186
rect 27836 8134 27888 8186
rect 27900 8134 27952 8186
rect 6828 8032 6880 8084
rect 6920 8075 6972 8084
rect 6920 8041 6929 8075
rect 6929 8041 6963 8075
rect 6963 8041 6972 8075
rect 6920 8032 6972 8041
rect 7012 8032 7064 8084
rect 7196 8032 7248 8084
rect 9772 8032 9824 8084
rect 9864 8032 9916 8084
rect 14556 8032 14608 8084
rect 18604 8032 18656 8084
rect 18696 8032 18748 8084
rect 18880 8032 18932 8084
rect 1400 7964 1452 8016
rect 4988 7964 5040 8016
rect 6092 7964 6144 8016
rect 6736 7964 6788 8016
rect 4896 7896 4948 7948
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 6184 7896 6236 7948
rect 6552 7939 6604 7948
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6552 7896 6604 7905
rect 2320 7760 2372 7812
rect 3240 7828 3292 7880
rect 4252 7828 4304 7880
rect 6368 7828 6420 7880
rect 7012 7896 7064 7948
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 7656 7939 7708 7948
rect 7656 7905 7665 7939
rect 7665 7905 7699 7939
rect 7699 7905 7708 7939
rect 7656 7896 7708 7905
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 9496 7964 9548 8016
rect 8852 7896 8904 7948
rect 9128 7896 9180 7948
rect 9680 7896 9732 7948
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 10968 7896 11020 7948
rect 8300 7828 8352 7880
rect 8668 7828 8720 7880
rect 8852 7803 8904 7812
rect 8852 7769 8861 7803
rect 8861 7769 8895 7803
rect 8895 7769 8904 7803
rect 8852 7760 8904 7769
rect 9312 7760 9364 7812
rect 9496 7803 9548 7812
rect 9496 7769 9505 7803
rect 9505 7769 9539 7803
rect 9539 7769 9548 7803
rect 9496 7760 9548 7769
rect 9956 7828 10008 7880
rect 11336 7964 11388 8016
rect 11612 8007 11664 8016
rect 11612 7973 11621 8007
rect 11621 7973 11655 8007
rect 11655 7973 11664 8007
rect 11612 7964 11664 7973
rect 13268 7964 13320 8016
rect 1952 7692 2004 7744
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 7012 7692 7064 7744
rect 7564 7692 7616 7744
rect 8208 7692 8260 7744
rect 8484 7692 8536 7744
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 11980 7896 12032 7948
rect 12716 7939 12768 7948
rect 12716 7905 12725 7939
rect 12725 7905 12759 7939
rect 12759 7905 12768 7939
rect 12716 7896 12768 7905
rect 12900 7896 12952 7948
rect 13176 7939 13228 7948
rect 13176 7905 13186 7939
rect 13186 7905 13220 7939
rect 13220 7905 13228 7939
rect 13176 7896 13228 7905
rect 13452 7939 13504 7948
rect 13452 7905 13461 7939
rect 13461 7905 13495 7939
rect 13495 7905 13504 7939
rect 13452 7896 13504 7905
rect 13544 7939 13596 7948
rect 13544 7905 13558 7939
rect 13558 7905 13592 7939
rect 13592 7905 13596 7939
rect 13544 7896 13596 7905
rect 13268 7760 13320 7812
rect 14004 7828 14056 7880
rect 14464 7828 14516 7880
rect 15844 7964 15896 8016
rect 16396 7964 16448 8016
rect 15108 7939 15160 7948
rect 15108 7905 15117 7939
rect 15117 7905 15151 7939
rect 15151 7905 15160 7939
rect 15108 7896 15160 7905
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 15384 7828 15436 7880
rect 16672 7828 16724 7880
rect 17040 7828 17092 7880
rect 17408 7760 17460 7812
rect 12532 7692 12584 7744
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 13912 7692 13964 7744
rect 14740 7692 14792 7744
rect 15108 7692 15160 7744
rect 15476 7692 15528 7744
rect 15660 7692 15712 7744
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 18880 7896 18932 7948
rect 18512 7828 18564 7880
rect 19616 8032 19668 8084
rect 24584 8032 24636 8084
rect 27528 8032 27580 8084
rect 27988 8032 28040 8084
rect 19800 7964 19852 8016
rect 20720 7896 20772 7948
rect 20904 7896 20956 7948
rect 22100 7896 22152 7948
rect 23020 7939 23072 7948
rect 23020 7905 23054 7939
rect 23054 7905 23072 7939
rect 23020 7896 23072 7905
rect 25596 7964 25648 8016
rect 24308 7896 24360 7948
rect 26792 7939 26844 7948
rect 26792 7905 26801 7939
rect 26801 7905 26835 7939
rect 26835 7905 26844 7939
rect 26792 7896 26844 7905
rect 27344 7896 27396 7948
rect 26240 7828 26292 7880
rect 25228 7760 25280 7812
rect 20996 7692 21048 7744
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 11436 7590 11488 7642
rect 11500 7590 11552 7642
rect 11564 7590 11616 7642
rect 11628 7590 11680 7642
rect 11692 7590 11744 7642
rect 19210 7590 19262 7642
rect 19274 7590 19326 7642
rect 19338 7590 19390 7642
rect 19402 7590 19454 7642
rect 19466 7590 19518 7642
rect 26984 7590 27036 7642
rect 27048 7590 27100 7642
rect 27112 7590 27164 7642
rect 27176 7590 27228 7642
rect 27240 7590 27292 7642
rect 3240 7531 3292 7540
rect 3240 7497 3249 7531
rect 3249 7497 3283 7531
rect 3283 7497 3292 7531
rect 3240 7488 3292 7497
rect 7656 7488 7708 7540
rect 7748 7488 7800 7540
rect 8944 7531 8996 7540
rect 8944 7497 8953 7531
rect 8953 7497 8987 7531
rect 8987 7497 8996 7531
rect 8944 7488 8996 7497
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 1952 7327 2004 7336
rect 1952 7293 1986 7327
rect 1986 7293 2004 7327
rect 1952 7284 2004 7293
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 4712 7352 4764 7404
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6552 7420 6604 7472
rect 6736 7352 6788 7404
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 3332 7216 3384 7268
rect 1216 7191 1268 7200
rect 1216 7157 1225 7191
rect 1225 7157 1259 7191
rect 1259 7157 1268 7191
rect 1216 7148 1268 7157
rect 3148 7148 3200 7200
rect 4160 7148 4212 7200
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 6552 7284 6604 7336
rect 6644 7216 6696 7268
rect 6920 7420 6972 7472
rect 6920 7284 6972 7336
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 10324 7420 10376 7472
rect 10692 7420 10744 7472
rect 13268 7463 13320 7472
rect 13268 7429 13277 7463
rect 13277 7429 13311 7463
rect 13311 7429 13320 7463
rect 13268 7420 13320 7429
rect 7196 7216 7248 7268
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 9772 7352 9824 7404
rect 13728 7488 13780 7540
rect 14004 7531 14056 7540
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 14464 7488 14516 7540
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 15108 7420 15160 7472
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10324 7327 10376 7336
rect 10324 7293 10333 7327
rect 10333 7293 10367 7327
rect 10367 7293 10376 7327
rect 10324 7284 10376 7293
rect 10600 7327 10652 7336
rect 10600 7293 10639 7327
rect 10639 7293 10652 7327
rect 10600 7284 10652 7293
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11336 7284 11388 7336
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 11888 7327 11940 7336
rect 11888 7293 11897 7327
rect 11897 7293 11931 7327
rect 11931 7293 11940 7327
rect 11888 7284 11940 7293
rect 13636 7284 13688 7336
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 9772 7148 9824 7200
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 11060 7259 11112 7268
rect 11060 7225 11069 7259
rect 11069 7225 11103 7259
rect 11103 7225 11112 7259
rect 11060 7216 11112 7225
rect 11612 7216 11664 7268
rect 13452 7216 13504 7268
rect 13728 7216 13780 7268
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 14924 7327 14976 7336
rect 14924 7293 14933 7327
rect 14933 7293 14967 7327
rect 14967 7293 14976 7327
rect 14924 7284 14976 7293
rect 15016 7327 15068 7336
rect 15016 7293 15026 7327
rect 15026 7293 15060 7327
rect 15060 7293 15068 7327
rect 15016 7284 15068 7293
rect 15200 7327 15252 7336
rect 15200 7293 15209 7327
rect 15209 7293 15243 7327
rect 15243 7293 15252 7327
rect 15200 7284 15252 7293
rect 15568 7420 15620 7472
rect 15568 7284 15620 7336
rect 15660 7327 15712 7336
rect 15660 7293 15669 7327
rect 15669 7293 15703 7327
rect 15703 7293 15712 7327
rect 15660 7284 15712 7293
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 15844 7284 15896 7293
rect 16120 7284 16172 7336
rect 18880 7488 18932 7540
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 20444 7352 20496 7404
rect 21456 7352 21508 7404
rect 16764 7327 16816 7336
rect 16764 7293 16773 7327
rect 16773 7293 16807 7327
rect 16807 7293 16816 7327
rect 16764 7284 16816 7293
rect 17408 7327 17460 7336
rect 17408 7293 17417 7327
rect 17417 7293 17451 7327
rect 17451 7293 17460 7327
rect 17408 7284 17460 7293
rect 13820 7148 13872 7200
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 15660 7148 15712 7200
rect 15752 7148 15804 7200
rect 16488 7191 16540 7200
rect 16488 7157 16497 7191
rect 16497 7157 16531 7191
rect 16531 7157 16540 7191
rect 16488 7148 16540 7157
rect 16764 7148 16816 7200
rect 18788 7327 18840 7336
rect 18788 7293 18797 7327
rect 18797 7293 18831 7327
rect 18831 7293 18840 7327
rect 18788 7284 18840 7293
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 20720 7284 20772 7336
rect 22376 7352 22428 7404
rect 23388 7352 23440 7404
rect 22744 7284 22796 7336
rect 24860 7284 24912 7336
rect 27344 7284 27396 7336
rect 30380 7284 30432 7336
rect 22100 7259 22152 7268
rect 22100 7225 22135 7259
rect 22135 7225 22152 7259
rect 22100 7216 22152 7225
rect 27528 7216 27580 7268
rect 22284 7148 22336 7200
rect 26240 7191 26292 7200
rect 26240 7157 26249 7191
rect 26249 7157 26283 7191
rect 26283 7157 26292 7191
rect 26240 7148 26292 7157
rect 26424 7148 26476 7200
rect 29092 7191 29144 7200
rect 29092 7157 29101 7191
rect 29101 7157 29135 7191
rect 29135 7157 29144 7191
rect 29092 7148 29144 7157
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 12096 7046 12148 7098
rect 12160 7046 12212 7098
rect 12224 7046 12276 7098
rect 12288 7046 12340 7098
rect 12352 7046 12404 7098
rect 19870 7046 19922 7098
rect 19934 7046 19986 7098
rect 19998 7046 20050 7098
rect 20062 7046 20114 7098
rect 20126 7046 20178 7098
rect 27644 7046 27696 7098
rect 27708 7046 27760 7098
rect 27772 7046 27824 7098
rect 27836 7046 27888 7098
rect 27900 7046 27952 7098
rect 2780 6944 2832 6996
rect 4160 6944 4212 6996
rect 1216 6808 1268 6860
rect 1952 6808 2004 6860
rect 3332 6876 3384 6928
rect 7840 6944 7892 6996
rect 9680 6944 9732 6996
rect 10232 6944 10284 6996
rect 10784 6944 10836 6996
rect 11888 6944 11940 6996
rect 6736 6919 6788 6928
rect 6736 6885 6745 6919
rect 6745 6885 6779 6919
rect 6779 6885 6788 6919
rect 6736 6876 6788 6885
rect 7380 6876 7432 6928
rect 2872 6851 2924 6860
rect 2872 6817 2906 6851
rect 2906 6817 2924 6851
rect 2872 6808 2924 6817
rect 3424 6808 3476 6860
rect 5080 6808 5132 6860
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 2964 6604 3016 6656
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6368 6851 6420 6860
rect 6368 6817 6377 6851
rect 6377 6817 6411 6851
rect 6411 6817 6420 6851
rect 6368 6808 6420 6817
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 6460 6808 6512 6817
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 6276 6672 6328 6724
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 7012 6808 7064 6860
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 8024 6808 8076 6817
rect 8576 6876 8628 6928
rect 11612 6876 11664 6928
rect 13728 6944 13780 6996
rect 15384 6987 15436 6996
rect 15384 6953 15393 6987
rect 15393 6953 15427 6987
rect 15427 6953 15436 6987
rect 15384 6944 15436 6953
rect 15476 6987 15528 6996
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 18972 6944 19024 6996
rect 22100 6944 22152 6996
rect 8208 6851 8260 6860
rect 8208 6817 8222 6851
rect 8222 6817 8256 6851
rect 8256 6817 8260 6851
rect 8208 6808 8260 6817
rect 9312 6808 9364 6860
rect 7196 6740 7248 6792
rect 7564 6740 7616 6792
rect 9036 6740 9088 6792
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 10968 6808 11020 6860
rect 11060 6851 11112 6860
rect 11060 6817 11069 6851
rect 11069 6817 11103 6851
rect 11103 6817 11112 6851
rect 11060 6808 11112 6817
rect 11980 6808 12032 6860
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 12900 6808 12952 6860
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 13544 6876 13596 6928
rect 15568 6876 15620 6928
rect 16120 6876 16172 6928
rect 13636 6851 13688 6860
rect 13636 6817 13645 6851
rect 13645 6817 13679 6851
rect 13679 6817 13688 6851
rect 13636 6808 13688 6817
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 14280 6851 14332 6860
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 7472 6715 7524 6724
rect 7472 6681 7481 6715
rect 7481 6681 7515 6715
rect 7515 6681 7524 6715
rect 7472 6672 7524 6681
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 8668 6604 8720 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 11244 6672 11296 6724
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 15476 6808 15528 6860
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 16396 6851 16448 6860
rect 16396 6817 16405 6851
rect 16405 6817 16439 6851
rect 16439 6817 16448 6851
rect 16396 6808 16448 6817
rect 15752 6740 15804 6792
rect 13912 6672 13964 6724
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 20444 6808 20496 6860
rect 20720 6851 20772 6860
rect 20720 6817 20729 6851
rect 20729 6817 20763 6851
rect 20763 6817 20772 6851
rect 20720 6808 20772 6817
rect 18788 6740 18840 6792
rect 10324 6604 10376 6656
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 16488 6604 16540 6656
rect 20444 6672 20496 6724
rect 20996 6808 21048 6860
rect 21824 6808 21876 6860
rect 21916 6851 21968 6860
rect 21916 6817 21925 6851
rect 21925 6817 21959 6851
rect 21959 6817 21968 6851
rect 21916 6808 21968 6817
rect 22284 6808 22336 6860
rect 21824 6672 21876 6724
rect 26240 6808 26292 6860
rect 26424 6851 26476 6860
rect 26424 6817 26433 6851
rect 26433 6817 26467 6851
rect 26467 6817 26476 6851
rect 26424 6808 26476 6817
rect 26148 6740 26200 6792
rect 26976 6808 27028 6860
rect 28080 6851 28132 6860
rect 28080 6817 28089 6851
rect 28089 6817 28123 6851
rect 28123 6817 28132 6851
rect 28080 6808 28132 6817
rect 29092 6876 29144 6928
rect 28908 6851 28960 6860
rect 28908 6817 28942 6851
rect 28942 6817 28960 6851
rect 28908 6808 28960 6817
rect 29276 6808 29328 6860
rect 18972 6604 19024 6656
rect 20996 6604 21048 6656
rect 21548 6647 21600 6656
rect 21548 6613 21557 6647
rect 21557 6613 21591 6647
rect 21591 6613 21600 6647
rect 21548 6604 21600 6613
rect 22008 6604 22060 6656
rect 23388 6604 23440 6656
rect 26056 6647 26108 6656
rect 26056 6613 26065 6647
rect 26065 6613 26099 6647
rect 26099 6613 26108 6647
rect 26056 6604 26108 6613
rect 27528 6672 27580 6724
rect 28356 6715 28408 6724
rect 28356 6681 28365 6715
rect 28365 6681 28399 6715
rect 28399 6681 28408 6715
rect 28356 6672 28408 6681
rect 26332 6604 26384 6656
rect 27436 6604 27488 6656
rect 28908 6604 28960 6656
rect 30012 6647 30064 6656
rect 30012 6613 30021 6647
rect 30021 6613 30055 6647
rect 30055 6613 30064 6647
rect 30012 6604 30064 6613
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 11436 6502 11488 6554
rect 11500 6502 11552 6554
rect 11564 6502 11616 6554
rect 11628 6502 11680 6554
rect 11692 6502 11744 6554
rect 19210 6502 19262 6554
rect 19274 6502 19326 6554
rect 19338 6502 19390 6554
rect 19402 6502 19454 6554
rect 19466 6502 19518 6554
rect 26984 6502 27036 6554
rect 27048 6502 27100 6554
rect 27112 6502 27164 6554
rect 27176 6502 27228 6554
rect 27240 6502 27292 6554
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 8024 6400 8076 6452
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 3148 6332 3200 6384
rect 3240 6375 3292 6384
rect 3240 6341 3249 6375
rect 3249 6341 3283 6375
rect 3283 6341 3292 6375
rect 3240 6332 3292 6341
rect 6276 6332 6328 6384
rect 7564 6332 7616 6384
rect 8392 6332 8444 6384
rect 9864 6400 9916 6452
rect 10324 6400 10376 6452
rect 15476 6400 15528 6452
rect 17132 6400 17184 6452
rect 18236 6400 18288 6452
rect 18788 6400 18840 6452
rect 21824 6400 21876 6452
rect 21916 6400 21968 6452
rect 26148 6400 26200 6452
rect 26240 6400 26292 6452
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 6092 6264 6144 6316
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 3516 6239 3568 6248
rect 3516 6205 3525 6239
rect 3525 6205 3559 6239
rect 3559 6205 3568 6239
rect 3516 6196 3568 6205
rect 4068 6196 4120 6248
rect 6368 6196 6420 6248
rect 6460 6196 6512 6248
rect 8300 6264 8352 6316
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 9496 6264 9548 6316
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 11244 6264 11296 6316
rect 12900 6332 12952 6384
rect 20444 6332 20496 6384
rect 20996 6332 21048 6384
rect 24860 6332 24912 6384
rect 27252 6332 27304 6384
rect 27988 6332 28040 6384
rect 16304 6264 16356 6316
rect 18420 6264 18472 6316
rect 19708 6264 19760 6316
rect 6736 6239 6788 6248
rect 6736 6205 6745 6239
rect 6745 6205 6779 6239
rect 6779 6205 6788 6239
rect 6736 6196 6788 6205
rect 7472 6196 7524 6248
rect 2688 6171 2740 6180
rect 2688 6137 2697 6171
rect 2697 6137 2731 6171
rect 2731 6137 2740 6171
rect 2688 6128 2740 6137
rect 3332 6128 3384 6180
rect 4160 6128 4212 6180
rect 6828 6171 6880 6180
rect 6828 6137 6837 6171
rect 6837 6137 6871 6171
rect 6871 6137 6880 6171
rect 6828 6128 6880 6137
rect 11704 6196 11756 6248
rect 11980 6196 12032 6248
rect 14832 6196 14884 6248
rect 18328 6196 18380 6248
rect 18696 6196 18748 6248
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 8944 6128 8996 6180
rect 9128 6128 9180 6180
rect 10416 6128 10468 6180
rect 18512 6128 18564 6180
rect 19064 6171 19116 6180
rect 19064 6137 19073 6171
rect 19073 6137 19107 6171
rect 19107 6137 19116 6171
rect 19064 6128 19116 6137
rect 2228 6060 2280 6112
rect 2780 6060 2832 6112
rect 6552 6060 6604 6112
rect 11888 6060 11940 6112
rect 12808 6060 12860 6112
rect 13084 6060 13136 6112
rect 13728 6060 13780 6112
rect 18880 6060 18932 6112
rect 19616 6171 19668 6180
rect 19616 6137 19625 6171
rect 19625 6137 19659 6171
rect 19659 6137 19668 6171
rect 19616 6128 19668 6137
rect 20628 6196 20680 6248
rect 21088 6196 21140 6248
rect 21732 6239 21784 6248
rect 21732 6205 21749 6239
rect 21749 6205 21784 6239
rect 21732 6196 21784 6205
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22468 6196 22520 6248
rect 23664 6196 23716 6248
rect 21456 6128 21508 6180
rect 22284 6128 22336 6180
rect 23388 6128 23440 6180
rect 24952 6239 25004 6248
rect 24952 6205 24961 6239
rect 24961 6205 24995 6239
rect 24995 6205 25004 6239
rect 24952 6196 25004 6205
rect 27436 6264 27488 6316
rect 27528 6264 27580 6316
rect 26424 6196 26476 6248
rect 25596 6128 25648 6180
rect 27436 6171 27488 6180
rect 27436 6137 27445 6171
rect 27445 6137 27479 6171
rect 27479 6137 27488 6171
rect 27436 6128 27488 6137
rect 27988 6239 28040 6248
rect 27988 6205 27997 6239
rect 27997 6205 28031 6239
rect 28031 6205 28040 6239
rect 27988 6196 28040 6205
rect 28080 6239 28132 6248
rect 28080 6205 28089 6239
rect 28089 6205 28123 6239
rect 28123 6205 28132 6239
rect 28080 6196 28132 6205
rect 30472 6239 30524 6248
rect 30472 6205 30481 6239
rect 30481 6205 30515 6239
rect 30515 6205 30524 6239
rect 30472 6196 30524 6205
rect 29920 6128 29972 6180
rect 26332 6060 26384 6112
rect 26700 6060 26752 6112
rect 28080 6060 28132 6112
rect 30012 6060 30064 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 12096 5958 12148 6010
rect 12160 5958 12212 6010
rect 12224 5958 12276 6010
rect 12288 5958 12340 6010
rect 12352 5958 12404 6010
rect 19870 5958 19922 6010
rect 19934 5958 19986 6010
rect 19998 5958 20050 6010
rect 20062 5958 20114 6010
rect 20126 5958 20178 6010
rect 27644 5958 27696 6010
rect 27708 5958 27760 6010
rect 27772 5958 27824 6010
rect 27836 5958 27888 6010
rect 27900 5958 27952 6010
rect 2872 5856 2924 5908
rect 8944 5856 8996 5908
rect 11704 5856 11756 5908
rect 1400 5720 1452 5772
rect 2228 5763 2280 5772
rect 2228 5729 2237 5763
rect 2237 5729 2271 5763
rect 2271 5729 2280 5763
rect 2228 5720 2280 5729
rect 2320 5763 2372 5772
rect 2320 5729 2329 5763
rect 2329 5729 2363 5763
rect 2363 5729 2372 5763
rect 2320 5720 2372 5729
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 8300 5788 8352 5840
rect 9404 5788 9456 5840
rect 4160 5720 4212 5772
rect 8392 5763 8444 5772
rect 8392 5729 8401 5763
rect 8401 5729 8435 5763
rect 8435 5729 8444 5763
rect 8392 5720 8444 5729
rect 8484 5763 8536 5772
rect 8484 5729 8494 5763
rect 8494 5729 8528 5763
rect 8528 5729 8536 5763
rect 8484 5720 8536 5729
rect 9588 5763 9640 5772
rect 9588 5729 9597 5763
rect 9597 5729 9631 5763
rect 9631 5729 9640 5763
rect 9588 5720 9640 5729
rect 11796 5788 11848 5840
rect 2780 5584 2832 5636
rect 6184 5584 6236 5636
rect 8576 5584 8628 5636
rect 9956 5584 10008 5636
rect 1676 5516 1728 5568
rect 1952 5516 2004 5568
rect 3148 5516 3200 5568
rect 11152 5559 11204 5568
rect 11152 5525 11161 5559
rect 11161 5525 11195 5559
rect 11195 5525 11204 5559
rect 11152 5516 11204 5525
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11888 5720 11940 5772
rect 13268 5856 13320 5908
rect 11612 5584 11664 5636
rect 11888 5584 11940 5636
rect 12164 5720 12216 5772
rect 15660 5856 15712 5908
rect 15752 5856 15804 5908
rect 22376 5856 22428 5908
rect 23388 5856 23440 5908
rect 25596 5899 25648 5908
rect 25596 5865 25605 5899
rect 25605 5865 25639 5899
rect 25639 5865 25648 5899
rect 25596 5856 25648 5865
rect 26700 5856 26752 5908
rect 27988 5856 28040 5908
rect 13544 5763 13596 5772
rect 13544 5729 13553 5763
rect 13553 5729 13587 5763
rect 13587 5729 13596 5763
rect 13544 5720 13596 5729
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 17960 5788 18012 5840
rect 18696 5831 18748 5840
rect 18696 5797 18705 5831
rect 18705 5797 18739 5831
rect 18739 5797 18748 5831
rect 18696 5788 18748 5797
rect 19064 5788 19116 5840
rect 26424 5831 26476 5840
rect 26424 5797 26433 5831
rect 26433 5797 26467 5831
rect 26467 5797 26476 5831
rect 26424 5788 26476 5797
rect 14004 5763 14056 5772
rect 14004 5729 14013 5763
rect 14013 5729 14047 5763
rect 14047 5729 14056 5763
rect 14004 5720 14056 5729
rect 14096 5763 14148 5772
rect 14096 5729 14105 5763
rect 14105 5729 14139 5763
rect 14139 5729 14148 5763
rect 14096 5720 14148 5729
rect 12808 5584 12860 5636
rect 13820 5652 13872 5704
rect 14372 5763 14424 5772
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 14556 5763 14608 5772
rect 14556 5729 14570 5763
rect 14570 5729 14604 5763
rect 14604 5729 14608 5763
rect 14556 5720 14608 5729
rect 14832 5763 14884 5772
rect 14832 5729 14841 5763
rect 14841 5729 14875 5763
rect 14875 5729 14884 5763
rect 14832 5720 14884 5729
rect 16396 5720 16448 5772
rect 18328 5720 18380 5772
rect 18880 5763 18932 5772
rect 18880 5729 18915 5763
rect 18915 5729 18932 5763
rect 18880 5720 18932 5729
rect 19616 5720 19668 5772
rect 14648 5652 14700 5704
rect 21916 5720 21968 5772
rect 22652 5763 22704 5772
rect 22652 5729 22661 5763
rect 22661 5729 22695 5763
rect 22695 5729 22704 5763
rect 22652 5720 22704 5729
rect 22744 5720 22796 5772
rect 24952 5720 25004 5772
rect 27344 5788 27396 5840
rect 14096 5584 14148 5636
rect 21824 5652 21876 5704
rect 26332 5652 26384 5704
rect 27528 5652 27580 5704
rect 12900 5516 12952 5568
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 13452 5516 13504 5568
rect 19708 5584 19760 5636
rect 14924 5516 14976 5568
rect 18328 5516 18380 5568
rect 18512 5516 18564 5568
rect 18696 5516 18748 5568
rect 21272 5516 21324 5568
rect 22008 5516 22060 5568
rect 23112 5516 23164 5568
rect 23940 5516 23992 5568
rect 26056 5516 26108 5568
rect 26240 5584 26292 5636
rect 28080 5720 28132 5772
rect 29276 5788 29328 5840
rect 29920 5899 29972 5908
rect 29920 5865 29929 5899
rect 29929 5865 29963 5899
rect 29963 5865 29972 5899
rect 29920 5856 29972 5865
rect 30472 5899 30524 5908
rect 30472 5865 30481 5899
rect 30481 5865 30515 5899
rect 30515 5865 30524 5899
rect 30472 5856 30524 5865
rect 28356 5652 28408 5704
rect 29092 5652 29144 5704
rect 30380 5763 30432 5772
rect 30380 5729 30389 5763
rect 30389 5729 30423 5763
rect 30423 5729 30432 5763
rect 30380 5720 30432 5729
rect 30472 5652 30524 5704
rect 30656 5584 30708 5636
rect 28080 5516 28132 5568
rect 29644 5516 29696 5568
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 11436 5414 11488 5466
rect 11500 5414 11552 5466
rect 11564 5414 11616 5466
rect 11628 5414 11680 5466
rect 11692 5414 11744 5466
rect 19210 5414 19262 5466
rect 19274 5414 19326 5466
rect 19338 5414 19390 5466
rect 19402 5414 19454 5466
rect 19466 5414 19518 5466
rect 26984 5414 27036 5466
rect 27048 5414 27100 5466
rect 27112 5414 27164 5466
rect 27176 5414 27228 5466
rect 27240 5414 27292 5466
rect 2780 5312 2832 5364
rect 4068 5312 4120 5364
rect 5172 5312 5224 5364
rect 8300 5312 8352 5364
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 3608 5244 3660 5296
rect 8484 5244 8536 5296
rect 7380 5176 7432 5228
rect 8852 5219 8904 5228
rect 8852 5185 8861 5219
rect 8861 5185 8895 5219
rect 8895 5185 8904 5219
rect 8852 5176 8904 5185
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 1952 5151 2004 5160
rect 1952 5117 1986 5151
rect 1986 5117 2004 5151
rect 1952 5108 2004 5117
rect 6184 5108 6236 5160
rect 4252 5040 4304 5092
rect 7840 5040 7892 5092
rect 10048 5151 10100 5160
rect 10048 5117 10057 5151
rect 10057 5117 10091 5151
rect 10091 5117 10100 5151
rect 10048 5108 10100 5117
rect 11152 5312 11204 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 13636 5312 13688 5364
rect 15016 5312 15068 5364
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 18052 5312 18104 5364
rect 18512 5312 18564 5364
rect 21456 5312 21508 5364
rect 14372 5244 14424 5296
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 13268 5176 13320 5228
rect 13636 5176 13688 5228
rect 14556 5219 14608 5228
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 18696 5244 18748 5296
rect 13820 5108 13872 5160
rect 9864 5040 9916 5092
rect 3424 4972 3476 5024
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 5080 4972 5132 5024
rect 12808 5040 12860 5092
rect 14464 5108 14516 5160
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 14924 5151 14976 5160
rect 14924 5117 14933 5151
rect 14933 5117 14967 5151
rect 14967 5117 14976 5151
rect 14924 5108 14976 5117
rect 15016 5151 15068 5160
rect 15016 5117 15025 5151
rect 15025 5117 15059 5151
rect 15059 5117 15068 5151
rect 15016 5108 15068 5117
rect 15200 5108 15252 5160
rect 16120 5151 16172 5160
rect 16120 5117 16155 5151
rect 16155 5117 16172 5151
rect 16120 5108 16172 5117
rect 15936 5083 15988 5092
rect 15936 5049 15945 5083
rect 15945 5049 15979 5083
rect 15979 5049 15988 5083
rect 15936 5040 15988 5049
rect 13820 4972 13872 5024
rect 14924 4972 14976 5024
rect 15752 4972 15804 5024
rect 15844 4972 15896 5024
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 17132 5151 17184 5160
rect 17132 5117 17141 5151
rect 17141 5117 17175 5151
rect 17175 5117 17184 5151
rect 17132 5108 17184 5117
rect 17592 5108 17644 5160
rect 18420 5176 18472 5228
rect 21824 5244 21876 5296
rect 22008 5244 22060 5296
rect 22100 5244 22152 5296
rect 22652 5312 22704 5364
rect 18328 5151 18380 5160
rect 18328 5117 18337 5151
rect 18337 5117 18371 5151
rect 18371 5117 18380 5151
rect 18328 5108 18380 5117
rect 21548 5176 21600 5228
rect 21916 5219 21968 5228
rect 21916 5185 21925 5219
rect 21925 5185 21959 5219
rect 21959 5185 21968 5219
rect 21916 5176 21968 5185
rect 18512 5040 18564 5092
rect 21640 5151 21692 5160
rect 21640 5117 21649 5151
rect 21649 5117 21683 5151
rect 21683 5117 21692 5151
rect 21640 5108 21692 5117
rect 22008 5151 22060 5160
rect 22008 5117 22017 5151
rect 22017 5117 22051 5151
rect 22051 5117 22060 5151
rect 22008 5108 22060 5117
rect 22744 5176 22796 5228
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 30564 5244 30616 5296
rect 23388 5219 23440 5228
rect 23388 5185 23397 5219
rect 23397 5185 23431 5219
rect 23431 5185 23440 5219
rect 23388 5176 23440 5185
rect 25044 5176 25096 5228
rect 26240 5219 26292 5228
rect 26240 5185 26258 5219
rect 26258 5185 26292 5219
rect 26240 5176 26292 5185
rect 26332 5219 26384 5228
rect 26332 5185 26341 5219
rect 26341 5185 26375 5219
rect 26375 5185 26384 5219
rect 26332 5176 26384 5185
rect 26608 5219 26660 5228
rect 26608 5185 26617 5219
rect 26617 5185 26651 5219
rect 26651 5185 26660 5219
rect 26608 5176 26660 5185
rect 26884 5176 26936 5228
rect 27344 5176 27396 5228
rect 22468 5108 22520 5117
rect 23664 5151 23716 5160
rect 23664 5117 23673 5151
rect 23673 5117 23707 5151
rect 23707 5117 23716 5151
rect 23664 5108 23716 5117
rect 27436 5108 27488 5160
rect 29368 5151 29420 5160
rect 29368 5117 29377 5151
rect 29377 5117 29411 5151
rect 29411 5117 29420 5151
rect 29368 5108 29420 5117
rect 29460 5108 29512 5160
rect 29644 5151 29696 5160
rect 29644 5117 29653 5151
rect 29653 5117 29687 5151
rect 29687 5117 29696 5151
rect 29644 5108 29696 5117
rect 30472 5108 30524 5160
rect 21732 5083 21784 5092
rect 21732 5049 21767 5083
rect 21767 5049 21784 5083
rect 21732 5040 21784 5049
rect 19616 4972 19668 5024
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 21640 4972 21692 5024
rect 22376 5083 22428 5092
rect 22376 5049 22385 5083
rect 22385 5049 22419 5083
rect 22419 5049 22428 5083
rect 22376 5040 22428 5049
rect 23020 5083 23072 5092
rect 23020 5049 23029 5083
rect 23029 5049 23063 5083
rect 23063 5049 23072 5083
rect 23020 5040 23072 5049
rect 28908 5040 28960 5092
rect 30656 5151 30708 5160
rect 30656 5117 30665 5151
rect 30665 5117 30699 5151
rect 30699 5117 30708 5151
rect 30656 5108 30708 5117
rect 23572 5015 23624 5024
rect 23572 4981 23581 5015
rect 23581 4981 23615 5015
rect 23615 4981 23624 5015
rect 23572 4972 23624 4981
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 28724 5015 28776 5024
rect 28724 4981 28733 5015
rect 28733 4981 28767 5015
rect 28767 4981 28776 5015
rect 28724 4972 28776 4981
rect 29000 4972 29052 5024
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 12096 4870 12148 4922
rect 12160 4870 12212 4922
rect 12224 4870 12276 4922
rect 12288 4870 12340 4922
rect 12352 4870 12404 4922
rect 19870 4870 19922 4922
rect 19934 4870 19986 4922
rect 19998 4870 20050 4922
rect 20062 4870 20114 4922
rect 20126 4870 20178 4922
rect 27644 4870 27696 4922
rect 27708 4870 27760 4922
rect 27772 4870 27824 4922
rect 27836 4870 27888 4922
rect 27900 4870 27952 4922
rect 3516 4768 3568 4820
rect 5172 4768 5224 4820
rect 6644 4768 6696 4820
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 10416 4768 10468 4820
rect 11244 4768 11296 4820
rect 13728 4768 13780 4820
rect 14648 4768 14700 4820
rect 18512 4768 18564 4820
rect 3332 4700 3384 4752
rect 4896 4700 4948 4752
rect 6920 4700 6972 4752
rect 8208 4700 8260 4752
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 2504 4632 2556 4684
rect 3148 4675 3200 4684
rect 3148 4641 3157 4675
rect 3157 4641 3191 4675
rect 3191 4641 3200 4675
rect 3148 4632 3200 4641
rect 3424 4675 3476 4684
rect 3424 4641 3458 4675
rect 3458 4641 3476 4675
rect 3424 4632 3476 4641
rect 4252 4496 4304 4548
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 11060 4632 11112 4684
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 13360 4632 13412 4684
rect 14924 4675 14976 4684
rect 14924 4641 14933 4675
rect 14933 4641 14967 4675
rect 14967 4641 14976 4675
rect 14924 4632 14976 4641
rect 16028 4700 16080 4752
rect 7656 4564 7708 4616
rect 10048 4496 10100 4548
rect 6276 4471 6328 4480
rect 6276 4437 6285 4471
rect 6285 4437 6319 4471
rect 6319 4437 6328 4471
rect 6276 4428 6328 4437
rect 13544 4428 13596 4480
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16488 4700 16540 4752
rect 16672 4700 16724 4752
rect 18236 4632 18288 4684
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 18604 4743 18656 4752
rect 18604 4709 18613 4743
rect 18613 4709 18647 4743
rect 18647 4709 18656 4743
rect 18604 4700 18656 4709
rect 20628 4700 20680 4752
rect 19616 4632 19668 4684
rect 20720 4675 20772 4684
rect 20720 4641 20729 4675
rect 20729 4641 20763 4675
rect 20763 4641 20772 4675
rect 20720 4632 20772 4641
rect 21640 4768 21692 4820
rect 25412 4768 25464 4820
rect 28080 4768 28132 4820
rect 29000 4811 29052 4820
rect 29000 4777 29009 4811
rect 29009 4777 29043 4811
rect 29043 4777 29052 4811
rect 29000 4768 29052 4777
rect 21180 4700 21232 4752
rect 21088 4675 21140 4684
rect 21088 4641 21097 4675
rect 21097 4641 21131 4675
rect 21131 4641 21140 4675
rect 21088 4632 21140 4641
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 23572 4700 23624 4752
rect 28172 4700 28224 4752
rect 29368 4768 29420 4820
rect 23112 4632 23164 4684
rect 28080 4675 28132 4684
rect 28080 4641 28089 4675
rect 28089 4641 28123 4675
rect 28123 4641 28132 4675
rect 28080 4632 28132 4641
rect 20076 4564 20128 4616
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 15936 4428 15988 4480
rect 17960 4428 18012 4480
rect 21548 4428 21600 4480
rect 22652 4471 22704 4480
rect 22652 4437 22661 4471
rect 22661 4437 22695 4471
rect 22695 4437 22704 4471
rect 22652 4428 22704 4437
rect 23020 4428 23072 4480
rect 25688 4496 25740 4548
rect 27988 4564 28040 4616
rect 28724 4632 28776 4684
rect 29000 4564 29052 4616
rect 28264 4539 28316 4548
rect 28264 4505 28273 4539
rect 28273 4505 28307 4539
rect 28307 4505 28316 4539
rect 28264 4496 28316 4505
rect 29092 4496 29144 4548
rect 25320 4471 25372 4480
rect 25320 4437 25329 4471
rect 25329 4437 25363 4471
rect 25363 4437 25372 4471
rect 25320 4428 25372 4437
rect 28540 4471 28592 4480
rect 28540 4437 28549 4471
rect 28549 4437 28583 4471
rect 28583 4437 28592 4471
rect 28540 4428 28592 4437
rect 29184 4428 29236 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 11436 4326 11488 4378
rect 11500 4326 11552 4378
rect 11564 4326 11616 4378
rect 11628 4326 11680 4378
rect 11692 4326 11744 4378
rect 19210 4326 19262 4378
rect 19274 4326 19326 4378
rect 19338 4326 19390 4378
rect 19402 4326 19454 4378
rect 19466 4326 19518 4378
rect 26984 4326 27036 4378
rect 27048 4326 27100 4378
rect 27112 4326 27164 4378
rect 27176 4326 27228 4378
rect 27240 4326 27292 4378
rect 2504 4224 2556 4276
rect 4068 4224 4120 4276
rect 4712 4224 4764 4276
rect 5172 4224 5224 4276
rect 6828 4224 6880 4276
rect 7840 4224 7892 4276
rect 8760 4224 8812 4276
rect 13084 4224 13136 4276
rect 14740 4224 14792 4276
rect 17132 4224 17184 4276
rect 17776 4267 17828 4276
rect 17776 4233 17785 4267
rect 17785 4233 17819 4267
rect 17819 4233 17828 4267
rect 17776 4224 17828 4233
rect 18328 4224 18380 4276
rect 19616 4224 19668 4276
rect 20076 4267 20128 4276
rect 20076 4233 20085 4267
rect 20085 4233 20119 4267
rect 20119 4233 20128 4267
rect 20076 4224 20128 4233
rect 21548 4224 21600 4276
rect 15844 4156 15896 4208
rect 15936 4088 15988 4140
rect 17316 4088 17368 4140
rect 20720 4156 20772 4208
rect 25320 4224 25372 4276
rect 25780 4224 25832 4276
rect 26608 4224 26660 4276
rect 3332 4020 3384 4072
rect 3516 4020 3568 4072
rect 3792 4020 3844 4072
rect 5356 4063 5408 4072
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 6644 4020 6696 4072
rect 8668 4020 8720 4072
rect 11060 4020 11112 4072
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 13820 4063 13872 4072
rect 13820 4029 13854 4063
rect 13854 4029 13872 4063
rect 13820 4020 13872 4029
rect 14372 4020 14424 4072
rect 16580 4020 16632 4072
rect 18328 4063 18380 4072
rect 18328 4029 18337 4063
rect 18337 4029 18371 4063
rect 18371 4029 18380 4063
rect 18328 4020 18380 4029
rect 3976 3995 4028 4004
rect 3976 3961 4010 3995
rect 4010 3961 4028 3995
rect 3976 3952 4028 3961
rect 5816 3952 5868 4004
rect 3332 3884 3384 3936
rect 10048 3952 10100 4004
rect 14004 3952 14056 4004
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 10968 3884 11020 3936
rect 17868 3884 17920 3936
rect 20076 4020 20128 4072
rect 24860 4156 24912 4208
rect 29092 4224 29144 4276
rect 21640 4088 21692 4140
rect 22652 4131 22704 4140
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 25688 4088 25740 4140
rect 21548 4063 21600 4072
rect 21548 4029 21557 4063
rect 21557 4029 21591 4063
rect 21591 4029 21600 4063
rect 21548 4020 21600 4029
rect 21088 3952 21140 4004
rect 22192 4063 22244 4072
rect 22192 4029 22201 4063
rect 22201 4029 22235 4063
rect 22235 4029 22244 4063
rect 22192 4020 22244 4029
rect 23020 4020 23072 4072
rect 23940 4020 23992 4072
rect 25044 4020 25096 4072
rect 27252 4088 27304 4140
rect 28080 4156 28132 4208
rect 29368 4224 29420 4276
rect 29460 4267 29512 4276
rect 29460 4233 29469 4267
rect 29469 4233 29503 4267
rect 29503 4233 29512 4267
rect 29460 4224 29512 4233
rect 28172 4131 28224 4140
rect 28172 4097 28181 4131
rect 28181 4097 28215 4131
rect 28215 4097 28224 4131
rect 28172 4088 28224 4097
rect 28264 4088 28316 4140
rect 26976 4063 27028 4072
rect 26976 4029 26994 4063
rect 26994 4029 27028 4063
rect 26976 4020 27028 4029
rect 23664 3952 23716 4004
rect 25044 3884 25096 3936
rect 30564 4063 30616 4072
rect 30564 4029 30582 4063
rect 30582 4029 30616 4063
rect 30564 4020 30616 4029
rect 30932 4063 30984 4072
rect 30932 4029 30941 4063
rect 30941 4029 30975 4063
rect 30975 4029 30984 4063
rect 30932 4020 30984 4029
rect 28816 3927 28868 3936
rect 28816 3893 28825 3927
rect 28825 3893 28859 3927
rect 28859 3893 28868 3927
rect 28816 3884 28868 3893
rect 29644 3884 29696 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 12096 3782 12148 3834
rect 12160 3782 12212 3834
rect 12224 3782 12276 3834
rect 12288 3782 12340 3834
rect 12352 3782 12404 3834
rect 19870 3782 19922 3834
rect 19934 3782 19986 3834
rect 19998 3782 20050 3834
rect 20062 3782 20114 3834
rect 20126 3782 20178 3834
rect 27644 3782 27696 3834
rect 27708 3782 27760 3834
rect 27772 3782 27824 3834
rect 27836 3782 27888 3834
rect 27900 3782 27952 3834
rect 3332 3723 3384 3732
rect 3332 3689 3341 3723
rect 3341 3689 3375 3723
rect 3375 3689 3384 3723
rect 3332 3680 3384 3689
rect 3792 3723 3844 3732
rect 3792 3689 3801 3723
rect 3801 3689 3835 3723
rect 3835 3689 3844 3723
rect 3792 3680 3844 3689
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 4068 3680 4120 3732
rect 4620 3680 4672 3732
rect 3240 3544 3292 3596
rect 3516 3587 3568 3596
rect 3516 3553 3525 3587
rect 3525 3553 3559 3587
rect 3559 3553 3568 3587
rect 3516 3544 3568 3553
rect 4160 3612 4212 3664
rect 5356 3680 5408 3732
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 7380 3680 7432 3732
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 5080 3544 5132 3596
rect 5632 3587 5684 3596
rect 5632 3553 5641 3587
rect 5641 3553 5675 3587
rect 5675 3553 5684 3587
rect 5632 3544 5684 3553
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 8576 3680 8628 3732
rect 6920 3544 6972 3596
rect 7564 3587 7616 3596
rect 7564 3553 7573 3587
rect 7573 3553 7607 3587
rect 7607 3553 7616 3587
rect 7564 3544 7616 3553
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 8484 3587 8536 3596
rect 8484 3553 8493 3587
rect 8493 3553 8527 3587
rect 8527 3553 8536 3587
rect 8484 3544 8536 3553
rect 8668 3655 8720 3664
rect 8668 3621 8677 3655
rect 8677 3621 8711 3655
rect 8711 3621 8720 3655
rect 8668 3612 8720 3621
rect 8668 3476 8720 3528
rect 8208 3408 8260 3460
rect 4712 3340 4764 3392
rect 7104 3340 7156 3392
rect 7656 3340 7708 3392
rect 8484 3340 8536 3392
rect 9772 3544 9824 3596
rect 8944 3476 8996 3528
rect 9404 3476 9456 3528
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 11060 3680 11112 3732
rect 14372 3680 14424 3732
rect 26976 3680 27028 3732
rect 28172 3680 28224 3732
rect 29000 3723 29052 3732
rect 29000 3689 29009 3723
rect 29009 3689 29043 3723
rect 29043 3689 29052 3723
rect 29000 3680 29052 3689
rect 20996 3655 21048 3664
rect 20996 3621 21005 3655
rect 21005 3621 21039 3655
rect 21039 3621 21048 3655
rect 20996 3612 21048 3621
rect 28540 3612 28592 3664
rect 28816 3612 28868 3664
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 10232 3476 10284 3528
rect 16488 3587 16540 3596
rect 16488 3553 16497 3587
rect 16497 3553 16531 3587
rect 16531 3553 16540 3587
rect 16488 3544 16540 3553
rect 19800 3544 19852 3596
rect 20352 3544 20404 3596
rect 28908 3587 28960 3596
rect 28908 3553 28917 3587
rect 28917 3553 28951 3587
rect 28951 3553 28960 3587
rect 28908 3544 28960 3553
rect 29092 3544 29144 3596
rect 21916 3519 21968 3528
rect 21916 3485 21925 3519
rect 21925 3485 21959 3519
rect 21959 3485 21968 3519
rect 21916 3476 21968 3485
rect 9956 3408 10008 3460
rect 14832 3408 14884 3460
rect 16856 3408 16908 3460
rect 15200 3340 15252 3392
rect 16212 3340 16264 3392
rect 19708 3340 19760 3392
rect 20260 3383 20312 3392
rect 20260 3349 20269 3383
rect 20269 3349 20303 3383
rect 20303 3349 20312 3383
rect 20260 3340 20312 3349
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 22100 3340 22152 3392
rect 25596 3340 25648 3392
rect 26608 3340 26660 3392
rect 27436 3340 27488 3392
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 11436 3238 11488 3290
rect 11500 3238 11552 3290
rect 11564 3238 11616 3290
rect 11628 3238 11680 3290
rect 11692 3238 11744 3290
rect 19210 3238 19262 3290
rect 19274 3238 19326 3290
rect 19338 3238 19390 3290
rect 19402 3238 19454 3290
rect 19466 3238 19518 3290
rect 26984 3238 27036 3290
rect 27048 3238 27100 3290
rect 27112 3238 27164 3290
rect 27176 3238 27228 3290
rect 27240 3238 27292 3290
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 7564 3136 7616 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 9772 3136 9824 3188
rect 10876 3136 10928 3188
rect 11152 3136 11204 3188
rect 11428 3136 11480 3188
rect 9956 3068 10008 3120
rect 11888 3136 11940 3188
rect 9680 3000 9732 3052
rect 5632 2932 5684 2984
rect 7104 2975 7156 2984
rect 7104 2941 7138 2975
rect 7138 2941 7156 2975
rect 7104 2932 7156 2941
rect 9864 2932 9916 2984
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 11060 3000 11112 3052
rect 10048 2864 10100 2916
rect 10968 2932 11020 2984
rect 11796 2932 11848 2984
rect 14924 3136 14976 3188
rect 17776 3136 17828 3188
rect 16120 3068 16172 3120
rect 22100 3136 22152 3188
rect 22192 3136 22244 3188
rect 24860 3136 24912 3188
rect 25596 3111 25648 3120
rect 25596 3077 25605 3111
rect 25605 3077 25639 3111
rect 25639 3077 25648 3111
rect 25596 3068 25648 3077
rect 27160 3136 27212 3188
rect 21916 3043 21968 3052
rect 13176 2932 13228 2984
rect 13544 2932 13596 2984
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 12440 2864 12492 2916
rect 15016 2932 15068 2984
rect 16028 2975 16080 2984
rect 16028 2941 16037 2975
rect 16037 2941 16071 2975
rect 16071 2941 16080 2975
rect 16028 2932 16080 2941
rect 16396 2932 16448 2984
rect 21916 3009 21925 3043
rect 21925 3009 21959 3043
rect 21959 3009 21968 3043
rect 21916 3000 21968 3009
rect 22376 3000 22428 3052
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25044 3000 25096 3009
rect 27528 3068 27580 3120
rect 26516 3043 26568 3052
rect 26516 3009 26525 3043
rect 26525 3009 26559 3043
rect 26559 3009 26568 3043
rect 26516 3000 26568 3009
rect 27436 3000 27488 3052
rect 16764 2932 16816 2984
rect 17316 2975 17368 2984
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 11520 2796 11572 2848
rect 11980 2796 12032 2848
rect 13084 2796 13136 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 14096 2839 14148 2848
rect 14096 2805 14105 2839
rect 14105 2805 14139 2839
rect 14139 2805 14148 2839
rect 14096 2796 14148 2805
rect 15016 2796 15068 2848
rect 20260 2932 20312 2984
rect 20996 2975 21048 2984
rect 20996 2941 21005 2975
rect 21005 2941 21039 2975
rect 21039 2941 21048 2975
rect 20996 2932 21048 2941
rect 19616 2864 19668 2916
rect 16396 2839 16448 2848
rect 16396 2805 16405 2839
rect 16405 2805 16439 2839
rect 16439 2805 16448 2839
rect 16396 2796 16448 2805
rect 16948 2796 17000 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 22008 2975 22060 2984
rect 22008 2941 22042 2975
rect 22042 2941 22060 2975
rect 22008 2932 22060 2941
rect 23664 2932 23716 2984
rect 25228 2975 25280 2984
rect 25228 2941 25246 2975
rect 25246 2941 25280 2975
rect 25228 2932 25280 2941
rect 25320 2975 25372 2984
rect 25320 2941 25329 2975
rect 25329 2941 25363 2975
rect 25363 2941 25372 2975
rect 25320 2932 25372 2941
rect 26240 2975 26292 2984
rect 26240 2941 26249 2975
rect 26249 2941 26283 2975
rect 26283 2941 26292 2975
rect 26240 2932 26292 2941
rect 26700 2975 26752 2984
rect 26700 2941 26709 2975
rect 26709 2941 26743 2975
rect 26743 2941 26752 2975
rect 26700 2932 26752 2941
rect 26792 2975 26844 2984
rect 26792 2941 26801 2975
rect 26801 2941 26835 2975
rect 26835 2941 26844 2975
rect 26792 2932 26844 2941
rect 27068 2932 27120 2984
rect 27988 3000 28040 3052
rect 28816 2975 28868 2984
rect 28816 2941 28825 2975
rect 28825 2941 28859 2975
rect 28859 2941 28868 2975
rect 28816 2932 28868 2941
rect 29092 2932 29144 2984
rect 27344 2864 27396 2916
rect 27436 2864 27488 2916
rect 30932 2932 30984 2984
rect 21640 2796 21692 2848
rect 22192 2796 22244 2848
rect 23756 2796 23808 2848
rect 26700 2796 26752 2848
rect 26884 2839 26936 2848
rect 26884 2805 26893 2839
rect 26893 2805 26927 2839
rect 26927 2805 26936 2839
rect 26884 2796 26936 2805
rect 27068 2839 27120 2848
rect 27068 2805 27095 2839
rect 27095 2805 27120 2839
rect 27068 2796 27120 2805
rect 28816 2796 28868 2848
rect 29000 2796 29052 2848
rect 29092 2839 29144 2848
rect 29092 2805 29101 2839
rect 29101 2805 29135 2839
rect 29135 2805 29144 2839
rect 29092 2796 29144 2805
rect 29368 2839 29420 2848
rect 29368 2805 29377 2839
rect 29377 2805 29411 2839
rect 29411 2805 29420 2839
rect 29368 2796 29420 2805
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 12096 2694 12148 2746
rect 12160 2694 12212 2746
rect 12224 2694 12276 2746
rect 12288 2694 12340 2746
rect 12352 2694 12404 2746
rect 19870 2694 19922 2746
rect 19934 2694 19986 2746
rect 19998 2694 20050 2746
rect 20062 2694 20114 2746
rect 20126 2694 20178 2746
rect 27644 2694 27696 2746
rect 27708 2694 27760 2746
rect 27772 2694 27824 2746
rect 27836 2694 27888 2746
rect 27900 2694 27952 2746
rect 9496 2456 9548 2508
rect 11244 2592 11296 2644
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10232 2456 10284 2508
rect 10692 2524 10744 2576
rect 11152 2567 11204 2576
rect 11152 2533 11179 2567
rect 11179 2533 11204 2567
rect 11152 2524 11204 2533
rect 10876 2456 10928 2508
rect 10968 2456 11020 2508
rect 10416 2388 10468 2440
rect 10692 2320 10744 2372
rect 9312 2252 9364 2304
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10232 2252 10284 2304
rect 11612 2456 11664 2508
rect 12348 2456 12400 2508
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 16948 2592 17000 2644
rect 23664 2592 23716 2644
rect 27436 2592 27488 2644
rect 13084 2567 13136 2576
rect 13084 2533 13093 2567
rect 13093 2533 13127 2567
rect 13127 2533 13136 2567
rect 13084 2524 13136 2533
rect 14096 2524 14148 2576
rect 14832 2524 14884 2576
rect 17500 2524 17552 2576
rect 19800 2524 19852 2576
rect 11704 2388 11756 2440
rect 12072 2388 12124 2440
rect 14004 2456 14056 2508
rect 11888 2320 11940 2372
rect 11152 2295 11204 2304
rect 11152 2261 11161 2295
rect 11161 2261 11195 2295
rect 11195 2261 11204 2295
rect 11152 2252 11204 2261
rect 11612 2252 11664 2304
rect 15384 2456 15436 2508
rect 16028 2456 16080 2508
rect 16212 2499 16264 2508
rect 16212 2465 16221 2499
rect 16221 2465 16255 2499
rect 16255 2465 16264 2499
rect 16212 2456 16264 2465
rect 15936 2388 15988 2440
rect 18236 2499 18288 2508
rect 18236 2465 18245 2499
rect 18245 2465 18279 2499
rect 18279 2465 18288 2499
rect 18236 2456 18288 2465
rect 19708 2499 19760 2508
rect 19708 2465 19717 2499
rect 19717 2465 19751 2499
rect 19751 2465 19760 2499
rect 19708 2456 19760 2465
rect 19984 2499 20036 2508
rect 19984 2465 20018 2499
rect 20018 2465 20036 2499
rect 19984 2456 20036 2465
rect 20996 2456 21048 2508
rect 21640 2499 21692 2508
rect 21640 2465 21649 2499
rect 21649 2465 21683 2499
rect 21683 2465 21692 2499
rect 21640 2456 21692 2465
rect 24124 2524 24176 2576
rect 26516 2524 26568 2576
rect 26792 2524 26844 2576
rect 29092 2524 29144 2576
rect 22652 2456 22704 2508
rect 23756 2499 23808 2508
rect 23756 2465 23765 2499
rect 23765 2465 23799 2499
rect 23799 2465 23808 2499
rect 23756 2456 23808 2465
rect 23848 2456 23900 2508
rect 25228 2456 25280 2508
rect 25780 2456 25832 2508
rect 26240 2456 26292 2508
rect 27160 2499 27212 2508
rect 27160 2465 27169 2499
rect 27169 2465 27203 2499
rect 27203 2465 27212 2499
rect 27160 2456 27212 2465
rect 27344 2456 27396 2508
rect 29368 2456 29420 2508
rect 21456 2431 21508 2440
rect 21456 2397 21465 2431
rect 21465 2397 21499 2431
rect 21499 2397 21508 2431
rect 21456 2388 21508 2397
rect 15200 2320 15252 2372
rect 15752 2252 15804 2304
rect 22008 2388 22060 2440
rect 22284 2431 22336 2440
rect 22284 2397 22293 2431
rect 22293 2397 22327 2431
rect 22327 2397 22336 2431
rect 22284 2388 22336 2397
rect 22100 2320 22152 2372
rect 16580 2252 16632 2304
rect 16856 2252 16908 2304
rect 21272 2295 21324 2304
rect 21272 2261 21281 2295
rect 21281 2261 21315 2295
rect 21315 2261 21324 2295
rect 21272 2252 21324 2261
rect 21364 2252 21416 2304
rect 22376 2295 22428 2304
rect 22376 2261 22385 2295
rect 22385 2261 22419 2295
rect 22419 2261 22428 2295
rect 22376 2252 22428 2261
rect 25320 2320 25372 2372
rect 24400 2252 24452 2304
rect 25228 2295 25280 2304
rect 25228 2261 25237 2295
rect 25237 2261 25271 2295
rect 25271 2261 25280 2295
rect 25228 2252 25280 2261
rect 25504 2320 25556 2372
rect 27252 2320 27304 2372
rect 27528 2320 27580 2372
rect 25872 2252 25924 2304
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 11436 2150 11488 2202
rect 11500 2150 11552 2202
rect 11564 2150 11616 2202
rect 11628 2150 11680 2202
rect 11692 2150 11744 2202
rect 19210 2150 19262 2202
rect 19274 2150 19326 2202
rect 19338 2150 19390 2202
rect 19402 2150 19454 2202
rect 19466 2150 19518 2202
rect 26984 2150 27036 2202
rect 27048 2150 27100 2202
rect 27112 2150 27164 2202
rect 27176 2150 27228 2202
rect 27240 2150 27292 2202
rect 9772 2048 9824 2100
rect 11336 1980 11388 2032
rect 9496 1844 9548 1896
rect 11244 1887 11296 1896
rect 11244 1853 11253 1887
rect 11253 1853 11287 1887
rect 11287 1853 11296 1887
rect 11244 1844 11296 1853
rect 11428 1844 11480 1896
rect 11796 2091 11848 2100
rect 11796 2057 11805 2091
rect 11805 2057 11839 2091
rect 11839 2057 11848 2091
rect 11796 2048 11848 2057
rect 14924 2048 14976 2100
rect 15752 2091 15804 2100
rect 15752 2057 15761 2091
rect 15761 2057 15795 2091
rect 15795 2057 15804 2091
rect 15752 2048 15804 2057
rect 15936 2091 15988 2100
rect 15936 2057 15945 2091
rect 15945 2057 15979 2091
rect 15979 2057 15988 2091
rect 15936 2048 15988 2057
rect 16672 2048 16724 2100
rect 11612 2023 11664 2032
rect 11612 1989 11621 2023
rect 11621 1989 11655 2023
rect 11655 1989 11664 2023
rect 11612 1980 11664 1989
rect 15384 2023 15436 2032
rect 15384 1989 15393 2023
rect 15393 1989 15427 2023
rect 15427 1989 15436 2023
rect 15384 1980 15436 1989
rect 17040 2048 17092 2100
rect 19984 2091 20036 2100
rect 19984 2057 19993 2091
rect 19993 2057 20027 2091
rect 20027 2057 20036 2091
rect 19984 2048 20036 2057
rect 20260 2048 20312 2100
rect 11796 1912 11848 1964
rect 11980 1912 12032 1964
rect 11704 1844 11756 1896
rect 11612 1776 11664 1828
rect 10232 1708 10284 1760
rect 11796 1751 11848 1760
rect 11796 1717 11813 1751
rect 11813 1717 11848 1751
rect 11796 1708 11848 1717
rect 12072 1887 12124 1896
rect 12072 1853 12081 1887
rect 12081 1853 12115 1887
rect 12115 1853 12124 1887
rect 12072 1844 12124 1853
rect 12348 1912 12400 1964
rect 12992 1844 13044 1896
rect 13544 1955 13596 1964
rect 13544 1921 13553 1955
rect 13553 1921 13587 1955
rect 13587 1921 13596 1955
rect 13544 1912 13596 1921
rect 17500 1980 17552 2032
rect 19708 1980 19760 2032
rect 20812 2048 20864 2100
rect 22008 2048 22060 2100
rect 22284 2048 22336 2100
rect 18236 1912 18288 1964
rect 11980 1819 12032 1828
rect 11980 1785 11989 1819
rect 11989 1785 12023 1819
rect 12023 1785 12032 1819
rect 11980 1776 12032 1785
rect 12164 1776 12216 1828
rect 14832 1819 14884 1828
rect 14832 1785 14841 1819
rect 14841 1785 14875 1819
rect 14875 1785 14884 1819
rect 14832 1776 14884 1785
rect 15016 1819 15068 1828
rect 15016 1785 15041 1819
rect 15041 1785 15068 1819
rect 16028 1887 16080 1896
rect 16028 1853 16037 1887
rect 16037 1853 16071 1887
rect 16071 1853 16080 1887
rect 16028 1844 16080 1853
rect 16120 1844 16172 1896
rect 17776 1844 17828 1896
rect 19800 1912 19852 1964
rect 20628 1980 20680 2032
rect 21456 1980 21508 2032
rect 22652 2091 22704 2100
rect 22652 2057 22661 2091
rect 22661 2057 22695 2091
rect 22695 2057 22704 2091
rect 22652 2048 22704 2057
rect 24124 2048 24176 2100
rect 24400 2048 24452 2100
rect 25320 2048 25372 2100
rect 25872 2048 25924 2100
rect 26884 2048 26936 2100
rect 27344 2048 27396 2100
rect 23756 1980 23808 2032
rect 23848 2023 23900 2032
rect 23848 1989 23857 2023
rect 23857 1989 23891 2023
rect 23891 1989 23900 2023
rect 23848 1980 23900 1989
rect 23940 1980 23992 2032
rect 15016 1776 15068 1785
rect 16488 1776 16540 1828
rect 20996 1844 21048 1896
rect 22008 1889 22060 1896
rect 22008 1855 22017 1889
rect 22017 1855 22051 1889
rect 22051 1855 22060 1889
rect 22008 1844 22060 1855
rect 22192 1844 22244 1896
rect 21272 1776 21324 1828
rect 21456 1776 21508 1828
rect 21732 1819 21784 1828
rect 21732 1785 21741 1819
rect 21741 1785 21775 1819
rect 21775 1785 21784 1819
rect 21732 1776 21784 1785
rect 13084 1751 13136 1760
rect 13084 1717 13093 1751
rect 13093 1717 13127 1751
rect 13127 1717 13136 1751
rect 13084 1708 13136 1717
rect 13268 1751 13320 1760
rect 13268 1717 13277 1751
rect 13277 1717 13311 1751
rect 13311 1717 13320 1751
rect 13268 1708 13320 1717
rect 13820 1708 13872 1760
rect 17592 1751 17644 1760
rect 17592 1717 17601 1751
rect 17601 1717 17635 1751
rect 17635 1717 17644 1751
rect 17592 1708 17644 1717
rect 17776 1751 17828 1760
rect 17776 1717 17785 1751
rect 17785 1717 17819 1751
rect 17819 1717 17828 1751
rect 17776 1708 17828 1717
rect 18328 1751 18380 1760
rect 18328 1717 18337 1751
rect 18337 1717 18371 1751
rect 18371 1717 18380 1751
rect 18328 1708 18380 1717
rect 19432 1751 19484 1760
rect 19432 1717 19441 1751
rect 19441 1717 19475 1751
rect 19475 1717 19484 1751
rect 19432 1708 19484 1717
rect 23204 1887 23256 1896
rect 23204 1853 23213 1887
rect 23213 1853 23247 1887
rect 23247 1853 23256 1887
rect 23204 1844 23256 1853
rect 24400 1887 24452 1896
rect 24400 1853 24409 1887
rect 24409 1853 24443 1887
rect 24443 1853 24452 1887
rect 24400 1844 24452 1853
rect 25136 1887 25188 1896
rect 25136 1853 25145 1887
rect 25145 1853 25179 1887
rect 25179 1853 25188 1887
rect 25136 1844 25188 1853
rect 25228 1844 25280 1896
rect 23940 1776 23992 1828
rect 25596 1819 25648 1828
rect 25596 1785 25605 1819
rect 25605 1785 25639 1819
rect 25639 1785 25648 1819
rect 25596 1776 25648 1785
rect 25780 1887 25832 1896
rect 25780 1853 25789 1887
rect 25789 1853 25823 1887
rect 25823 1853 25832 1887
rect 25780 1844 25832 1853
rect 25872 1887 25924 1896
rect 25872 1853 25881 1887
rect 25881 1853 25915 1887
rect 25915 1853 25924 1887
rect 25872 1844 25924 1853
rect 26148 1980 26200 2032
rect 26516 1955 26568 1964
rect 26516 1921 26525 1955
rect 26525 1921 26559 1955
rect 26559 1921 26568 1955
rect 26516 1912 26568 1921
rect 27068 1844 27120 1896
rect 28448 1887 28500 1896
rect 28448 1853 28457 1887
rect 28457 1853 28491 1887
rect 28491 1853 28500 1887
rect 28448 1844 28500 1853
rect 27988 1776 28040 1828
rect 25412 1751 25464 1760
rect 25412 1717 25429 1751
rect 25429 1717 25464 1751
rect 25412 1708 25464 1717
rect 26148 1708 26200 1760
rect 26516 1751 26568 1760
rect 26516 1717 26525 1751
rect 26525 1717 26559 1751
rect 26559 1717 26568 1751
rect 26516 1708 26568 1717
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 12096 1606 12148 1658
rect 12160 1606 12212 1658
rect 12224 1606 12276 1658
rect 12288 1606 12340 1658
rect 12352 1606 12404 1658
rect 19870 1606 19922 1658
rect 19934 1606 19986 1658
rect 19998 1606 20050 1658
rect 20062 1606 20114 1658
rect 20126 1606 20178 1658
rect 27644 1606 27696 1658
rect 27708 1606 27760 1658
rect 27772 1606 27824 1658
rect 27836 1606 27888 1658
rect 27900 1606 27952 1658
rect 9956 1504 10008 1556
rect 11612 1504 11664 1556
rect 11980 1504 12032 1556
rect 16028 1504 16080 1556
rect 13084 1436 13136 1488
rect 14924 1436 14976 1488
rect 16764 1504 16816 1556
rect 19708 1504 19760 1556
rect 20996 1504 21048 1556
rect 21732 1504 21784 1556
rect 22192 1504 22244 1556
rect 23204 1504 23256 1556
rect 25136 1504 25188 1556
rect 25596 1504 25648 1556
rect 27068 1547 27120 1556
rect 27068 1513 27077 1547
rect 27077 1513 27111 1547
rect 27111 1513 27120 1547
rect 27068 1504 27120 1513
rect 28448 1504 28500 1556
rect 17592 1479 17644 1488
rect 17592 1445 17610 1479
rect 17610 1445 17644 1479
rect 17592 1436 17644 1445
rect 20260 1436 20312 1488
rect 22284 1436 22336 1488
rect 23756 1436 23808 1488
rect 26700 1436 26752 1488
rect 9312 1411 9364 1420
rect 9312 1377 9321 1411
rect 9321 1377 9355 1411
rect 9355 1377 9364 1411
rect 9312 1368 9364 1377
rect 9588 1411 9640 1420
rect 9588 1377 9622 1411
rect 9622 1377 9640 1411
rect 9588 1368 9640 1377
rect 11244 1368 11296 1420
rect 11888 1411 11940 1420
rect 11888 1377 11897 1411
rect 11897 1377 11931 1411
rect 11931 1377 11940 1411
rect 11888 1368 11940 1377
rect 13268 1368 13320 1420
rect 16488 1368 16540 1420
rect 19432 1368 19484 1420
rect 21364 1368 21416 1420
rect 21548 1411 21600 1420
rect 21548 1377 21582 1411
rect 21582 1377 21600 1411
rect 21548 1368 21600 1377
rect 23664 1368 23716 1420
rect 25412 1411 25464 1420
rect 25412 1377 25421 1411
rect 25421 1377 25455 1411
rect 25455 1377 25464 1411
rect 25412 1368 25464 1377
rect 26516 1368 26568 1420
rect 26884 1368 26936 1420
rect 27436 1411 27488 1420
rect 27436 1377 27445 1411
rect 27445 1377 27479 1411
rect 27479 1377 27488 1411
rect 27436 1368 27488 1377
rect 18328 1300 18380 1352
rect 26240 1300 26292 1352
rect 27988 1232 28040 1284
rect 11336 1164 11388 1216
rect 12992 1164 13044 1216
rect 25596 1207 25648 1216
rect 25596 1173 25605 1207
rect 25605 1173 25639 1207
rect 25639 1173 25648 1207
rect 25596 1164 25648 1173
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 11436 1062 11488 1114
rect 11500 1062 11552 1114
rect 11564 1062 11616 1114
rect 11628 1062 11680 1114
rect 11692 1062 11744 1114
rect 19210 1062 19262 1114
rect 19274 1062 19326 1114
rect 19338 1062 19390 1114
rect 19402 1062 19454 1114
rect 19466 1062 19518 1114
rect 26984 1062 27036 1114
rect 27048 1062 27100 1114
rect 27112 1062 27164 1114
rect 27176 1062 27228 1114
rect 27240 1062 27292 1114
rect 9588 960 9640 1012
rect 11336 1003 11388 1012
rect 11336 969 11345 1003
rect 11345 969 11379 1003
rect 11379 969 11388 1003
rect 11336 960 11388 969
rect 21548 960 21600 1012
rect 26240 960 26292 1012
rect 10232 935 10284 944
rect 10232 901 10241 935
rect 10241 901 10275 935
rect 10275 901 10284 935
rect 10232 892 10284 901
rect 9404 824 9456 876
rect 13820 824 13872 876
rect 9956 756 10008 808
rect 10692 799 10744 808
rect 10692 765 10701 799
rect 10701 765 10735 799
rect 10735 765 10744 799
rect 10692 756 10744 765
rect 11980 756 12032 808
rect 20812 799 20864 808
rect 20812 765 20821 799
rect 20821 765 20855 799
rect 20855 765 20864 799
rect 20812 756 20864 765
rect 22376 756 22428 808
rect 23664 756 23716 808
rect 25596 756 25648 808
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 12096 518 12148 570
rect 12160 518 12212 570
rect 12224 518 12276 570
rect 12288 518 12340 570
rect 12352 518 12404 570
rect 19870 518 19922 570
rect 19934 518 19986 570
rect 19998 518 20050 570
rect 20062 518 20114 570
rect 20126 518 20178 570
rect 27644 518 27696 570
rect 27708 518 27760 570
rect 27772 518 27824 570
rect 27836 518 27888 570
rect 27900 518 27952 570
<< metal2 >>
rect 11794 21992 11850 22001
rect 11794 21927 11850 21936
rect 12254 21992 12310 22001
rect 12254 21927 12310 21936
rect 23846 21992 23902 22001
rect 23846 21927 23902 21936
rect 24950 21992 25006 22001
rect 24950 21927 25006 21936
rect 25502 21992 25558 22001
rect 25502 21927 25558 21936
rect 26054 21992 26110 22001
rect 26054 21927 26110 21936
rect 27526 21992 27582 22001
rect 27526 21927 27582 21936
rect 28262 21992 28318 22001
rect 28262 21927 28318 21936
rect 8666 21856 8722 21865
rect 3662 21788 3970 21797
rect 8666 21791 8722 21800
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 6458 21720 6514 21729
rect 6458 21655 6460 21664
rect 6512 21655 6514 21664
rect 7286 21720 7342 21729
rect 7286 21655 7288 21664
rect 6460 21626 6512 21632
rect 7340 21655 7342 21664
rect 8390 21720 8446 21729
rect 8680 21690 8708 21791
rect 11436 21788 11744 21797
rect 11436 21786 11442 21788
rect 11498 21786 11522 21788
rect 11578 21786 11602 21788
rect 11658 21786 11682 21788
rect 11738 21786 11744 21788
rect 11498 21734 11500 21786
rect 11680 21734 11682 21786
rect 11436 21732 11442 21734
rect 11498 21732 11522 21734
rect 11578 21732 11602 21734
rect 11658 21732 11682 21734
rect 11738 21732 11744 21734
rect 9954 21720 10010 21729
rect 8390 21655 8392 21664
rect 7288 21626 7340 21632
rect 8444 21655 8446 21664
rect 8668 21684 8720 21690
rect 8392 21626 8444 21632
rect 9954 21655 9956 21664
rect 8668 21626 8720 21632
rect 10008 21655 10010 21664
rect 10322 21720 10378 21729
rect 11436 21723 11744 21732
rect 11808 21690 11836 21927
rect 12268 21690 12296 21927
rect 21638 21856 21694 21865
rect 19210 21788 19518 21797
rect 21638 21791 21694 21800
rect 19210 21786 19216 21788
rect 19272 21786 19296 21788
rect 19352 21786 19376 21788
rect 19432 21786 19456 21788
rect 19512 21786 19518 21788
rect 19272 21734 19274 21786
rect 19454 21734 19456 21786
rect 19210 21732 19216 21734
rect 19272 21732 19296 21734
rect 19352 21732 19376 21734
rect 19432 21732 19456 21734
rect 19512 21732 19518 21734
rect 12806 21720 12862 21729
rect 19210 21723 19518 21732
rect 10322 21655 10324 21664
rect 9956 21626 10008 21632
rect 10376 21655 10378 21664
rect 11796 21684 11848 21690
rect 10324 21626 10376 21632
rect 11796 21626 11848 21632
rect 12256 21684 12308 21690
rect 12806 21655 12808 21664
rect 12256 21626 12308 21632
rect 12860 21655 12862 21664
rect 12808 21626 12860 21632
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 4068 21616 4120 21622
rect 4068 21558 4120 21564
rect 11702 21584 11758 21593
rect 3344 21486 3372 21558
rect 3516 21548 3568 21554
rect 3516 21490 3568 21496
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 2412 21412 2464 21418
rect 2412 21354 2464 21360
rect 2424 21010 2452 21354
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2516 21010 2544 21286
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2504 21004 2556 21010
rect 2504 20946 2556 20952
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2240 20398 2268 20742
rect 2332 20602 2360 20946
rect 2700 20806 2728 21422
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 2792 20398 2820 21286
rect 3252 21146 3280 21422
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1964 19922 1992 20198
rect 1952 19916 2004 19922
rect 1952 19858 2004 19864
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 1860 18148 1912 18154
rect 1860 18090 1912 18096
rect 1308 18080 1360 18086
rect 1308 18022 1360 18028
rect 1320 17746 1348 18022
rect 1308 17740 1360 17746
rect 1308 17682 1360 17688
rect 1872 16726 1900 18090
rect 1860 16720 1912 16726
rect 1860 16662 1912 16668
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16114 1624 16594
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1596 14958 1624 16050
rect 1688 15570 1716 16390
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 1964 15065 1992 19246
rect 2148 18970 2176 19246
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2056 18154 2084 18702
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2148 18154 2176 18566
rect 2240 18222 2268 20334
rect 3252 20330 3280 21082
rect 3344 20398 3372 21422
rect 3424 21412 3476 21418
rect 3424 21354 3476 21360
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3240 20324 3292 20330
rect 3240 20266 3292 20272
rect 2412 19984 2464 19990
rect 2412 19926 2464 19932
rect 2424 19514 2452 19926
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 3252 19446 3280 20266
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3240 19440 3292 19446
rect 2976 19378 3188 19394
rect 3240 19382 3292 19388
rect 2976 19372 3200 19378
rect 2976 19366 3148 19372
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2424 18834 2452 19246
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2044 18148 2096 18154
rect 2044 18090 2096 18096
rect 2136 18148 2188 18154
rect 2136 18090 2188 18096
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 17338 2268 17682
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2424 16046 2452 16526
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 1950 15056 2006 15065
rect 1950 14991 2006 15000
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14482 1716 14758
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1964 14074 1992 14894
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2240 14550 2268 14758
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1872 11608 1900 12650
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12306 1992 12582
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 2056 11626 2084 12718
rect 2516 11694 2544 19246
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2608 19122 2636 19178
rect 2608 19094 2728 19122
rect 2700 18834 2728 19094
rect 2976 18902 3004 19366
rect 3148 19314 3200 19320
rect 3344 19310 3372 20198
rect 3436 19922 3464 21354
rect 3528 21078 3556 21490
rect 4080 21486 4108 21558
rect 8024 21548 8076 21554
rect 11702 21519 11758 21528
rect 16670 21584 16726 21593
rect 16670 21519 16726 21528
rect 19430 21584 19486 21593
rect 19430 21519 19486 21528
rect 8024 21490 8076 21496
rect 4068 21480 4120 21486
rect 3988 21440 4068 21468
rect 3988 21146 4016 21440
rect 4068 21422 4120 21428
rect 4252 21480 4304 21486
rect 4252 21422 4304 21428
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 3516 21072 3568 21078
rect 3516 21014 3568 21020
rect 4080 21010 4108 21286
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 4264 20602 4292 21422
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 6196 21078 6224 21286
rect 6274 21176 6330 21185
rect 6274 21111 6276 21120
rect 6328 21111 6330 21120
rect 6276 21082 6328 21088
rect 5356 21072 5408 21078
rect 5356 21014 5408 21020
rect 6184 21072 6236 21078
rect 6184 21014 6236 21020
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 4448 20466 4476 20946
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 4632 20398 4660 20946
rect 5092 20466 5212 20482
rect 5080 20460 5212 20466
rect 5132 20454 5212 20460
rect 5080 20402 5132 20408
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4620 20392 4672 20398
rect 4804 20392 4856 20398
rect 4672 20352 4752 20380
rect 4620 20334 4672 20340
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2688 18828 2740 18834
rect 2740 18788 2820 18816
rect 2688 18770 2740 18776
rect 2608 18426 2636 18770
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2700 17814 2728 18158
rect 2688 17808 2740 17814
rect 2688 17750 2740 17756
rect 2792 17134 2820 18788
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2884 17134 2912 18090
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2700 16182 2728 17070
rect 2688 16176 2740 16182
rect 2688 16118 2740 16124
rect 2792 15314 2820 17070
rect 2976 16590 3004 17274
rect 3068 17270 3096 19246
rect 3528 19174 3556 19858
rect 4080 19718 4108 20334
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 4724 19990 4752 20352
rect 4804 20334 4856 20340
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4816 19854 4844 20334
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4908 19786 4936 20198
rect 5000 20058 5028 20334
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 4080 19310 4108 19654
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 3148 17128 3200 17134
rect 3068 17088 3148 17116
rect 3068 16658 3096 17088
rect 3436 17105 3464 18770
rect 3620 18766 3648 19178
rect 3974 18864 4030 18873
rect 3974 18799 4030 18808
rect 3988 18766 4016 18799
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3528 17882 3556 18634
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3528 17746 3556 17818
rect 3804 17746 3832 18022
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3976 17536 4028 17542
rect 4080 17524 4108 19246
rect 4172 19174 4200 19654
rect 4908 19378 4936 19722
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4264 18873 4292 19314
rect 4712 19236 4764 19242
rect 4712 19178 4764 19184
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 4250 18864 4306 18873
rect 4250 18799 4306 18808
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 18086 4200 18702
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18154 4384 18566
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4264 17882 4292 18090
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4028 17496 4108 17524
rect 4160 17536 4212 17542
rect 3976 17478 4028 17484
rect 4160 17478 4212 17484
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 4172 17134 4200 17478
rect 4160 17128 4212 17134
rect 3148 17070 3200 17076
rect 3422 17096 3478 17105
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3332 17060 3384 17066
rect 4160 17070 4212 17076
rect 3422 17031 3478 17040
rect 3332 17002 3384 17008
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2976 16250 3004 16526
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2884 15586 2912 16118
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15706 3004 15846
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2884 15558 3004 15586
rect 2976 15434 3004 15558
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2872 15360 2924 15366
rect 2792 15308 2872 15314
rect 2792 15302 2924 15308
rect 3068 15314 3096 16594
rect 3160 15502 3188 16730
rect 3252 16658 3280 17002
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 2792 15286 2912 15302
rect 3068 15286 3188 15314
rect 2792 15042 2820 15286
rect 2608 15014 2820 15042
rect 2608 14958 2636 15014
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2792 13530 2820 14894
rect 3068 14074 3096 14894
rect 3160 14770 3188 15286
rect 3252 14958 3280 16594
rect 3344 16590 3372 17002
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3344 16182 3372 16526
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3344 16046 3372 16118
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3436 15434 3464 16934
rect 4264 16658 4292 17682
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4448 17202 4476 17614
rect 4724 17610 4752 19178
rect 5092 18970 5120 19178
rect 5184 18970 5212 20454
rect 5368 20058 5396 21014
rect 6472 21010 6500 21422
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 6840 21010 6868 21286
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 5460 20466 5488 20742
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5368 19922 5396 19994
rect 6012 19922 6040 20402
rect 6288 19922 6316 20742
rect 7024 20330 7052 21286
rect 8036 20398 8064 21490
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 8312 21146 8340 21422
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 8482 21176 8538 21185
rect 8300 21140 8352 21146
rect 8482 21111 8484 21120
rect 8300 21082 8352 21088
rect 8536 21111 8538 21120
rect 8484 21082 8536 21088
rect 8312 21010 8340 21082
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6012 19786 6040 19858
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6012 19334 6040 19722
rect 6288 19514 6316 19858
rect 6472 19514 6500 19858
rect 7024 19854 7052 20266
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5920 19306 6040 19334
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5184 18834 5212 18906
rect 5828 18902 5856 19246
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5184 17746 5212 18770
rect 5920 18426 5948 19306
rect 6368 19304 6420 19310
rect 6366 19272 6368 19281
rect 6460 19304 6512 19310
rect 6420 19272 6422 19281
rect 6184 19236 6236 19242
rect 6460 19246 6512 19252
rect 6366 19207 6422 19216
rect 6184 19178 6236 19184
rect 6196 18970 6224 19178
rect 6276 19168 6328 19174
rect 6472 19156 6500 19246
rect 6328 19128 6500 19156
rect 6276 19110 6328 19116
rect 6564 18970 6592 19722
rect 6920 19304 6972 19310
rect 6642 19272 6698 19281
rect 6920 19246 6972 19252
rect 6642 19207 6644 19216
rect 6696 19207 6698 19216
rect 6644 19178 6696 19184
rect 6184 18964 6236 18970
rect 6552 18964 6604 18970
rect 6236 18924 6316 18952
rect 6184 18906 6236 18912
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5816 17808 5868 17814
rect 5920 17796 5948 18362
rect 5868 17768 5948 17796
rect 5816 17750 5868 17756
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 4080 16250 4108 16526
rect 5828 16454 5856 17750
rect 6104 17746 6132 18838
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 3896 15706 3924 15846
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3988 15638 4016 15846
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3712 15473 3740 15506
rect 3698 15464 3754 15473
rect 3424 15428 3476 15434
rect 3698 15399 3754 15408
rect 3424 15370 3476 15376
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3436 14890 3464 15370
rect 3804 15366 3832 15506
rect 4080 15366 4108 15846
rect 4172 15638 4200 15914
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3160 14742 3280 14770
rect 3252 14346 3280 14742
rect 3436 14618 3464 14826
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3528 14482 3556 15302
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 4172 15026 4200 15574
rect 4264 15434 4292 15982
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4724 15706 4752 15914
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 5644 15570 5672 15982
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5540 15496 5592 15502
rect 5262 15464 5318 15473
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4804 15428 4856 15434
rect 5540 15438 5592 15444
rect 5262 15399 5318 15408
rect 4804 15370 4856 15376
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14482 3648 14758
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3160 13870 3188 14214
rect 3252 13938 3280 14282
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 3252 13462 3280 13670
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3528 13190 3556 14418
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 4172 13530 4200 14962
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 14482 4292 14758
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4724 13802 4752 15030
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 12434 2820 12718
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 2792 12406 2912 12434
rect 2792 12306 2820 12406
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 1952 11620 2004 11626
rect 1872 11580 1952 11608
rect 1952 11562 2004 11568
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2056 11218 2084 11562
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2056 10606 2084 11154
rect 2608 10810 2636 11154
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2792 10606 2820 11562
rect 2884 10674 2912 12406
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3436 11830 3464 12242
rect 3528 11898 3556 12650
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3790 11792 3846 11801
rect 3436 11694 3464 11766
rect 4080 11778 4108 12310
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4448 11801 4476 12242
rect 4816 12238 4844 15370
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4908 14521 4936 15098
rect 5000 14550 5028 15302
rect 4988 14544 5040 14550
rect 4894 14512 4950 14521
rect 4988 14486 5040 14492
rect 4894 14447 4950 14456
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4434 11792 4490 11801
rect 3988 11762 4200 11778
rect 4264 11762 4384 11778
rect 3790 11727 3846 11736
rect 3884 11756 3936 11762
rect 3804 11694 3832 11727
rect 3884 11698 3936 11704
rect 3988 11756 4212 11762
rect 3988 11750 4160 11756
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3528 11354 3556 11562
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3620 10996 3648 11562
rect 3896 11540 3924 11698
rect 3988 11694 4016 11750
rect 4160 11698 4212 11704
rect 4264 11756 4396 11762
rect 4264 11750 4344 11756
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 4080 11540 4108 11591
rect 3896 11512 4108 11540
rect 3528 10968 3648 10996
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 10130 1992 10406
rect 2056 10198 2084 10542
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9722 1624 9998
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9178 1716 9454
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1780 8974 1808 9862
rect 2056 9722 2084 10134
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2056 9110 2084 9658
rect 2884 9518 2912 10610
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2976 9722 3004 10066
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3068 9674 3096 10746
rect 3528 10198 3556 10968
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3240 9920 3292 9926
rect 3238 9888 3240 9897
rect 3292 9888 3294 9897
rect 3238 9823 3294 9832
rect 3238 9752 3294 9761
rect 3294 9710 3372 9738
rect 3238 9687 3294 9696
rect 3068 9646 3188 9674
rect 3160 9602 3188 9646
rect 3160 9574 3280 9602
rect 3252 9518 3280 9574
rect 2872 9512 2924 9518
rect 3240 9512 3292 9518
rect 2872 9454 2924 9460
rect 3146 9480 3202 9489
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 2332 8634 2360 9386
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2884 8430 2912 9454
rect 3240 9454 3292 9460
rect 3146 9415 3148 9424
rect 3200 9415 3202 9424
rect 3148 9386 3200 9392
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9178 3004 9318
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3068 8430 3096 9046
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 1400 8016 1452 8022
rect 1400 7958 1452 7964
rect 3054 7984 3110 7993
rect 1412 7342 1440 7958
rect 3054 7919 3110 7928
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 7342 1992 7686
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1216 7200 1268 7206
rect 1216 7142 1268 7148
rect 1228 6866 1256 7142
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1412 5778 1440 7278
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1964 6458 1992 6802
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2134 6352 2190 6361
rect 2332 6322 2360 7754
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7002 2820 7686
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6497 2544 6598
rect 2502 6488 2558 6497
rect 2502 6423 2558 6432
rect 2134 6287 2190 6296
rect 2320 6316 2372 6322
rect 2148 6254 2176 6287
rect 2320 6258 2372 6264
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2240 5778 2268 6054
rect 2332 5778 2360 6258
rect 2596 6248 2648 6254
rect 2594 6216 2596 6225
rect 2780 6248 2832 6254
rect 2648 6216 2650 6225
rect 2780 6190 2832 6196
rect 2594 6151 2650 6160
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2700 5930 2728 6122
rect 2792 6118 2820 6190
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2700 5902 2820 5930
rect 2884 5914 2912 6802
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 1412 5166 1440 5714
rect 2792 5642 2820 5902
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2976 5778 3004 6598
rect 3068 6322 3096 7919
rect 3160 7206 3188 9386
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9042 3280 9318
rect 3344 9110 3372 9710
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7546 3280 7822
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3344 7274 3372 8910
rect 3436 8498 3464 9998
rect 3712 9926 3740 10066
rect 3804 10033 3832 10066
rect 4080 10033 4108 11512
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3790 10024 3846 10033
rect 3790 9959 3792 9968
rect 3844 9959 3846 9968
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 3792 9930 3844 9936
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3528 9654 3556 9862
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 3746 9716 3798 9722
rect 3712 9664 3746 9674
rect 3712 9658 3798 9664
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4066 9688 4122 9697
rect 3516 9648 3568 9654
rect 3712 9646 3786 9658
rect 3516 9590 3568 9596
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3516 9444 3568 9450
rect 3620 9432 3648 9551
rect 3712 9518 3740 9646
rect 3700 9512 3752 9518
rect 3988 9489 4016 9658
rect 4066 9623 4122 9632
rect 3700 9454 3752 9460
rect 3974 9480 4030 9489
rect 3568 9404 3648 9432
rect 3516 9386 3568 9392
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3424 7336 3476 7342
rect 3528 7324 3556 8978
rect 3620 8974 3648 9404
rect 3712 9081 3740 9454
rect 3974 9415 4030 9424
rect 3988 9110 4016 9415
rect 3976 9104 4028 9110
rect 3698 9072 3754 9081
rect 3976 9046 4028 9052
rect 3698 9007 3700 9016
rect 3752 9007 3754 9016
rect 3700 8978 3752 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 3476 7296 3556 7324
rect 3884 7336 3936 7342
rect 3882 7304 3884 7313
rect 3936 7304 3938 7313
rect 3424 7278 3476 7284
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 6390 3188 7142
rect 3344 6934 3372 7210
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3148 6384 3200 6390
rect 3240 6384 3292 6390
rect 3148 6326 3200 6332
rect 3238 6352 3240 6361
rect 3292 6352 3294 6361
rect 3056 6316 3108 6322
rect 3238 6287 3294 6296
rect 3056 6258 3108 6264
rect 3344 6186 3372 6870
rect 3436 6866 3464 7278
rect 3882 7239 3938 7248
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6254 3464 6802
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3514 6488 3570 6497
rect 3662 6491 3970 6500
rect 3514 6423 3570 6432
rect 3528 6254 3556 6423
rect 4080 6254 4108 9623
rect 4172 9042 4200 10474
rect 4264 10130 4292 11750
rect 4434 11727 4490 11736
rect 4344 11698 4396 11704
rect 4448 11694 4476 11727
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 4816 10538 4844 12174
rect 4908 11762 4936 14447
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9518 4384 9998
rect 4448 9722 4476 10134
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4264 8838 4292 9386
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4724 8922 4752 10134
rect 4908 9722 4936 11494
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4908 9110 4936 9522
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4632 8906 4752 8922
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4620 8900 4752 8906
rect 4672 8894 4752 8900
rect 4620 8842 4672 8848
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 8634 4752 8774
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4264 7886 4292 8366
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4434 7440 4490 7449
rect 4724 7410 4752 8570
rect 5000 8362 5028 8910
rect 4988 8356 5040 8362
rect 4988 8298 5040 8304
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7954 4936 8230
rect 5000 8022 5028 8298
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4434 7375 4490 7384
rect 4712 7404 4764 7410
rect 4448 7342 4476 7375
rect 4712 7346 4764 7352
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4160 7200 4212 7206
rect 4448 7188 4476 7278
rect 4160 7142 4212 7148
rect 4264 7160 4476 7188
rect 4172 7002 4200 7142
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 3424 6248 3476 6254
rect 3422 6216 3424 6225
rect 3516 6248 3568 6254
rect 3476 6216 3478 6225
rect 3332 6180 3384 6186
rect 3516 6190 3568 6196
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4172 6186 4200 6938
rect 3422 6151 3478 6160
rect 4160 6180 4212 6186
rect 3332 6122 3384 6128
rect 4160 6122 4212 6128
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1688 4690 1716 5510
rect 1964 5166 1992 5510
rect 2792 5370 2820 5578
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 3160 4690 3188 5510
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 2516 4282 2544 4626
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 3344 4078 3372 4694
rect 3436 4690 3464 4966
rect 3528 4826 3556 4966
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3620 4570 3648 5238
rect 3528 4542 3648 4570
rect 3528 4078 3556 4542
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 4080 4282 4108 5306
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3332 4072 3384 4078
rect 3252 4020 3332 4026
rect 3252 4014 3384 4020
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3252 3998 3372 4014
rect 3252 3602 3280 3998
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3738 3372 3878
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3528 3602 3556 4014
rect 3804 3738 3832 4014
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3988 3738 4016 3946
rect 4080 3738 4108 4218
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4172 3670 4200 5714
rect 4264 5098 4292 7160
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4264 4554 4292 5034
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 4908 4758 4936 7890
rect 5092 6866 5120 12854
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5184 11354 5212 12378
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5276 11257 5304 15399
rect 5552 15162 5580 15438
rect 5644 15162 5672 15506
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5552 14618 5580 14962
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5552 12850 5580 14010
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5736 12646 5764 13262
rect 5920 12850 5948 14486
rect 6012 14482 6040 15438
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6012 14074 6040 14418
rect 6104 14414 6132 17478
rect 6196 16794 6224 18770
rect 6288 18222 6316 18924
rect 6552 18906 6604 18912
rect 6932 18834 6960 19246
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6932 18358 6960 18770
rect 7116 18630 7144 19994
rect 7196 19984 7248 19990
rect 7196 19926 7248 19932
rect 7208 19854 7236 19926
rect 8036 19922 8064 20334
rect 8220 19990 8248 20878
rect 8312 20398 8340 20946
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8404 20058 8432 20946
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8574 20632 8630 20641
rect 8574 20567 8576 20576
rect 8628 20567 8630 20576
rect 8576 20538 8628 20544
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7208 18970 7236 19790
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6656 17746 6684 18090
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6656 17338 6684 17682
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6840 17270 6868 17682
rect 6932 17678 6960 18294
rect 7668 18222 7696 19858
rect 8220 19310 8248 19926
rect 8496 19922 8524 20198
rect 8680 19990 8708 20742
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8956 20058 8984 20334
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 9784 19718 9812 21354
rect 9876 21146 9904 21422
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9784 19514 9812 19654
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 17746 7328 18022
rect 7392 17814 7420 18090
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7576 17746 7604 18022
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6932 17338 6960 17614
rect 7760 17338 7788 18158
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 7852 17066 7880 17818
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 7392 16726 7420 17002
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 16794 7696 16934
rect 7852 16810 7880 17002
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7760 16782 7880 16810
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6196 14890 6224 16594
rect 7760 16522 7788 16782
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7760 16182 7788 16458
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 7748 16176 7800 16182
rect 7748 16118 7800 16124
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 15706 6960 15914
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6748 15026 6776 15302
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6932 14890 6960 15642
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6104 13818 6132 14350
rect 6196 13870 6224 14826
rect 7024 14822 7052 16118
rect 7760 16046 7788 16118
rect 7852 16046 7880 16594
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15638 7236 15846
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7576 15366 7604 15914
rect 7852 15706 7880 15982
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7944 15366 7972 17070
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8036 16046 8064 16526
rect 8128 16250 8156 18770
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18222 8248 18566
rect 9416 18222 9444 18702
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9508 17882 9536 18090
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8220 16658 8248 17070
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8404 16590 8432 17478
rect 8680 17338 8708 17478
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 9402 17096 9458 17105
rect 8588 16794 8616 17070
rect 9402 17031 9458 17040
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7378 15056 7434 15065
rect 7378 14991 7434 15000
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 14618 7144 14758
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7208 14414 7236 14894
rect 7392 14822 7420 14991
rect 7380 14816 7432 14822
rect 7300 14776 7380 14804
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6012 13790 6132 13818
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6012 13274 6040 13790
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 13394 6132 13670
rect 6656 13462 6684 14214
rect 6932 13462 6960 14350
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13530 7236 14214
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6012 13246 6132 13274
rect 6104 12850 6132 13246
rect 7116 13190 7144 13330
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 7116 12714 7144 13126
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12442 6960 12582
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6932 12306 6960 12378
rect 7116 12306 7144 12650
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5262 11248 5318 11257
rect 5262 11183 5318 11192
rect 5356 11212 5408 11218
rect 5276 11150 5304 11183
rect 5356 11154 5408 11160
rect 5264 11144 5316 11150
rect 5184 11104 5264 11132
rect 5184 10810 5212 11104
rect 5264 11086 5316 11092
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5276 10606 5304 10950
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5368 10198 5396 11154
rect 5552 10606 5580 11630
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5736 11218 5764 11562
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11218 5856 11494
rect 5920 11342 6224 11370
rect 5920 11286 5948 11342
rect 6196 11286 6224 11342
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10470 5580 10542
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5552 9654 5580 10406
rect 5736 9926 5764 11154
rect 6104 10810 6132 11222
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6288 10538 6316 11698
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6460 10532 6512 10538
rect 6460 10474 6512 10480
rect 5920 10266 5948 10474
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 6288 10062 6316 10474
rect 6472 10198 6500 10474
rect 6460 10192 6512 10198
rect 6564 10169 6592 11290
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6460 10134 6512 10140
rect 6550 10160 6606 10169
rect 6748 10130 6776 10746
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6550 10095 6552 10104
rect 6604 10095 6606 10104
rect 6736 10124 6788 10130
rect 6552 10066 6604 10072
rect 6736 10066 6788 10072
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6840 9926 6868 10134
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5184 8430 5212 9590
rect 7024 9586 7052 12106
rect 7012 9580 7064 9586
rect 6840 9540 7012 9568
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 5184 7954 5212 8366
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 6104 7342 6132 7958
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6196 7410 6224 7890
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6092 6656 6144 6662
rect 6090 6624 6092 6633
rect 6144 6624 6146 6633
rect 6090 6559 6146 6568
rect 6104 6322 6132 6559
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6196 5642 6224 6734
rect 6288 6730 6316 8366
rect 6380 7886 6408 9318
rect 6840 9178 6868 9540
rect 7012 9522 7064 9528
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7024 9178 7052 9386
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6840 8430 6868 9114
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6932 8090 6960 8434
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6380 6866 6408 7822
rect 6564 7478 6592 7890
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 6748 7410 6776 7958
rect 6840 7562 6868 8026
rect 7024 7954 7052 8026
rect 7012 7948 7064 7954
rect 7116 7936 7144 12106
rect 7208 11694 7236 13466
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7208 10266 7236 10678
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7300 10130 7328 14776
rect 7380 14758 7432 14764
rect 7576 14618 7604 15302
rect 7840 14952 7892 14958
rect 8220 14940 8248 16458
rect 8496 16182 8524 16594
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8496 15570 8524 16118
rect 9048 15978 9076 16594
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 9048 15502 9076 15914
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9048 15026 9076 15438
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8300 14952 8352 14958
rect 8220 14912 8300 14940
rect 7840 14894 7892 14900
rect 8300 14894 8352 14900
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13870 7512 14214
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 13326 7512 13670
rect 7852 13394 7880 14894
rect 9048 14550 9076 14962
rect 9036 14544 9088 14550
rect 9036 14486 9088 14492
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7944 13734 7972 14350
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 9416 13394 9444 17031
rect 9508 16658 9536 17614
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9508 16250 9536 16594
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9508 16017 9536 16050
rect 9600 16046 9628 17070
rect 9692 16182 9720 17478
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9784 16250 9812 16390
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9588 16040 9640 16046
rect 9494 16008 9550 16017
rect 9588 15982 9640 15988
rect 9494 15943 9550 15952
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9600 15162 9628 15574
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9496 14952 9548 14958
rect 9692 14940 9720 15370
rect 9876 15026 9904 16934
rect 9968 16726 9996 21286
rect 10152 20398 10180 21286
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10244 20058 10272 20946
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10336 20602 10364 20878
rect 10520 20777 10548 21422
rect 11348 20942 11376 21422
rect 11716 21078 11744 21519
rect 16684 21486 16712 21519
rect 19444 21486 19472 21519
rect 21652 21486 21680 21791
rect 23860 21486 23888 21927
rect 24398 21856 24454 21865
rect 24398 21791 24454 21800
rect 24412 21486 24440 21791
rect 24964 21486 24992 21927
rect 25516 21486 25544 21927
rect 26068 21486 26096 21927
rect 26514 21856 26570 21865
rect 26514 21791 26570 21800
rect 26528 21554 26556 21791
rect 26984 21788 27292 21797
rect 26984 21786 26990 21788
rect 27046 21786 27070 21788
rect 27126 21786 27150 21788
rect 27206 21786 27230 21788
rect 27286 21786 27292 21788
rect 27046 21734 27048 21786
rect 27228 21734 27230 21786
rect 26984 21732 26990 21734
rect 27046 21732 27070 21734
rect 27126 21732 27150 21734
rect 27206 21732 27230 21734
rect 27286 21732 27292 21734
rect 26984 21723 27292 21732
rect 27540 21690 27568 21927
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 26884 21616 26936 21622
rect 26884 21558 26936 21564
rect 26516 21548 26568 21554
rect 26516 21490 26568 21496
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 18604 21480 18656 21486
rect 19432 21480 19484 21486
rect 18604 21422 18656 21428
rect 19246 21448 19302 21457
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12096 21244 12404 21253
rect 12096 21242 12102 21244
rect 12158 21242 12182 21244
rect 12238 21242 12262 21244
rect 12318 21242 12342 21244
rect 12398 21242 12404 21244
rect 12158 21190 12160 21242
rect 12340 21190 12342 21242
rect 12096 21188 12102 21190
rect 12158 21188 12182 21190
rect 12238 21188 12262 21190
rect 12318 21188 12342 21190
rect 12398 21188 12404 21190
rect 12096 21179 12404 21188
rect 11704 21072 11756 21078
rect 11704 21014 11756 21020
rect 12820 21010 12848 21286
rect 13740 21010 13768 21422
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 13818 21176 13874 21185
rect 13818 21111 13820 21120
rect 13872 21111 13874 21120
rect 13820 21082 13872 21088
rect 15474 21040 15530 21049
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12808 21004 12860 21010
rect 13728 21004 13780 21010
rect 12808 20946 12860 20952
rect 13648 20964 13728 20992
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 10506 20768 10562 20777
rect 10506 20703 10562 20712
rect 11436 20700 11744 20709
rect 11436 20698 11442 20700
rect 11498 20698 11522 20700
rect 11578 20698 11602 20700
rect 11658 20698 11682 20700
rect 11738 20698 11744 20700
rect 11498 20646 11500 20698
rect 11680 20646 11682 20698
rect 11436 20644 11442 20646
rect 11498 20644 11522 20646
rect 11578 20644 11602 20646
rect 11658 20644 11682 20646
rect 11738 20644 11744 20646
rect 11436 20635 11744 20644
rect 12084 20602 12112 20946
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12912 20641 12940 20810
rect 12898 20632 12954 20641
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 12072 20596 12124 20602
rect 12898 20567 12954 20576
rect 12072 20538 12124 20544
rect 13648 20398 13676 20964
rect 13728 20946 13780 20952
rect 15292 21004 15344 21010
rect 15474 20975 15476 20984
rect 15292 20946 15344 20952
rect 15528 20975 15530 20984
rect 15476 20946 15528 20952
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13740 20466 13768 20742
rect 13832 20641 13860 20810
rect 13818 20632 13874 20641
rect 13818 20567 13874 20576
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 20058 11100 20266
rect 12096 20156 12404 20165
rect 12096 20154 12102 20156
rect 12158 20154 12182 20156
rect 12238 20154 12262 20156
rect 12318 20154 12342 20156
rect 12398 20154 12404 20156
rect 12158 20102 12160 20154
rect 12340 20102 12342 20154
rect 12096 20100 12102 20102
rect 12158 20100 12182 20102
rect 12238 20100 12262 20102
rect 12318 20100 12342 20102
rect 12398 20100 12404 20102
rect 12096 20091 12404 20100
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11072 19310 11100 19858
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10048 18216 10100 18222
rect 10046 18184 10048 18193
rect 10100 18184 10102 18193
rect 10046 18119 10102 18128
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 16726 10088 18022
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10152 17785 10180 17818
rect 10138 17776 10194 17785
rect 10138 17711 10194 17720
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9968 16454 9996 16662
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 10060 16250 10088 16526
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9548 14912 9720 14940
rect 9496 14894 9548 14900
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13462 9628 14282
rect 9968 14278 9996 15506
rect 10152 15434 10180 17274
rect 10244 15570 10272 19246
rect 11072 18834 11100 19246
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10980 18426 11008 18702
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10520 18329 10548 18362
rect 10506 18320 10562 18329
rect 10506 18255 10562 18264
rect 10520 18222 10548 18255
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10704 17882 10732 18158
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10428 17134 10456 17478
rect 10520 17338 10548 17682
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10704 17134 10732 17818
rect 10888 17814 10916 18090
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10980 17270 11008 18362
rect 11164 17762 11192 19722
rect 11256 18970 11284 19790
rect 11436 19612 11744 19621
rect 11436 19610 11442 19612
rect 11498 19610 11522 19612
rect 11578 19610 11602 19612
rect 11658 19610 11682 19612
rect 11738 19610 11744 19612
rect 11498 19558 11500 19610
rect 11680 19558 11682 19610
rect 11436 19556 11442 19558
rect 11498 19556 11522 19558
rect 11578 19556 11602 19558
rect 11658 19556 11682 19558
rect 11738 19556 11744 19558
rect 11436 19547 11744 19556
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11440 18902 11468 19110
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11072 17734 11284 17762
rect 11348 17746 11376 18634
rect 11436 18524 11744 18533
rect 11436 18522 11442 18524
rect 11498 18522 11522 18524
rect 11578 18522 11602 18524
rect 11658 18522 11682 18524
rect 11738 18522 11744 18524
rect 11498 18470 11500 18522
rect 11680 18470 11682 18522
rect 11436 18468 11442 18470
rect 11498 18468 11522 18470
rect 11578 18468 11602 18470
rect 11658 18468 11682 18470
rect 11738 18468 11744 18470
rect 11436 18459 11744 18468
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11624 17882 11652 18090
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11072 17678 11100 17734
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10336 16046 10364 16594
rect 10428 16250 10456 17070
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15638 10364 15982
rect 10520 15978 10548 16458
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10508 15972 10560 15978
rect 10508 15914 10560 15920
rect 10324 15632 10376 15638
rect 10324 15574 10376 15580
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10230 15464 10286 15473
rect 10140 15428 10192 15434
rect 10230 15399 10232 15408
rect 10140 15370 10192 15376
rect 10284 15399 10286 15408
rect 10232 15370 10284 15376
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 7484 12782 7512 13262
rect 8220 12782 8248 13262
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12782 9076 13126
rect 9416 12918 9444 13330
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 7484 12306 7512 12718
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7392 11762 7420 12106
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7668 11694 7696 12582
rect 7760 12442 7788 12718
rect 9600 12442 9628 13398
rect 9968 13394 9996 14214
rect 10060 13802 10088 15030
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10244 14906 10272 15370
rect 10336 15162 10364 15574
rect 10612 15570 10640 16186
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10152 14550 10180 14894
rect 10244 14878 10364 14906
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10336 13394 10364 14878
rect 10428 14618 10456 15098
rect 10520 14890 10548 15370
rect 10612 15042 10640 15506
rect 10704 15434 10732 16594
rect 11072 16590 11100 17070
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16176 11020 16182
rect 11164 16164 11192 17546
rect 11020 16136 11192 16164
rect 10968 16118 11020 16124
rect 10784 16040 10836 16046
rect 10782 16008 10784 16017
rect 11152 16040 11204 16046
rect 10836 16008 10838 16017
rect 10782 15943 10838 15952
rect 10888 16000 11152 16028
rect 10796 15570 10824 15943
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10612 15026 10732 15042
rect 10612 15020 10744 15026
rect 10612 15014 10692 15020
rect 10692 14962 10744 14968
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10612 14618 10640 14894
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10704 14550 10732 14962
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 10508 14476 10560 14482
rect 10796 14464 10824 15506
rect 10888 14958 10916 16000
rect 11256 16028 11284 17734
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11348 17338 11376 17682
rect 11808 17649 11836 18770
rect 11900 18737 11928 19926
rect 12096 19068 12404 19077
rect 12096 19066 12102 19068
rect 12158 19066 12182 19068
rect 12238 19066 12262 19068
rect 12318 19066 12342 19068
rect 12398 19066 12404 19068
rect 12158 19014 12160 19066
rect 12340 19014 12342 19066
rect 12096 19012 12102 19014
rect 12158 19012 12182 19014
rect 12238 19012 12262 19014
rect 12318 19012 12342 19014
rect 12398 19012 12404 19014
rect 12096 19003 12404 19012
rect 11886 18728 11942 18737
rect 11886 18663 11942 18672
rect 12636 18222 12664 20334
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13372 19922 13400 20198
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13832 18970 13860 20334
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 19310 14596 19790
rect 14752 19310 14780 19994
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14844 18834 14872 19246
rect 15212 18902 15240 20198
rect 15304 19990 15332 20946
rect 15488 20058 15516 20946
rect 15580 20466 15608 21286
rect 15764 21010 15792 21286
rect 16592 21010 16620 21422
rect 16684 21146 16712 21422
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 15752 21004 15804 21010
rect 15752 20946 15804 20952
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15488 19718 15516 19858
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15304 19310 15332 19654
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 15304 18834 15332 19246
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 12096 17980 12404 17989
rect 12096 17978 12102 17980
rect 12158 17978 12182 17980
rect 12238 17978 12262 17980
rect 12318 17978 12342 17980
rect 12398 17978 12404 17980
rect 12158 17926 12160 17978
rect 12340 17926 12342 17978
rect 12096 17924 12102 17926
rect 12158 17924 12182 17926
rect 12238 17924 12262 17926
rect 12318 17924 12342 17926
rect 12398 17924 12404 17926
rect 12096 17915 12404 17924
rect 13266 17912 13322 17921
rect 13266 17847 13268 17856
rect 13320 17847 13322 17856
rect 13268 17818 13320 17824
rect 13648 17814 13676 18158
rect 14200 17882 14228 18158
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 13636 17808 13688 17814
rect 11978 17776 12034 17785
rect 13636 17750 13688 17756
rect 13818 17776 13874 17785
rect 11978 17711 12034 17720
rect 11992 17678 12020 17711
rect 11888 17672 11940 17678
rect 11794 17640 11850 17649
rect 11888 17614 11940 17620
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 11794 17575 11850 17584
rect 11436 17436 11744 17445
rect 11436 17434 11442 17436
rect 11498 17434 11522 17436
rect 11578 17434 11602 17436
rect 11658 17434 11682 17436
rect 11738 17434 11744 17436
rect 11498 17382 11500 17434
rect 11680 17382 11682 17434
rect 11436 17380 11442 17382
rect 11498 17380 11522 17382
rect 11578 17380 11602 17382
rect 11658 17380 11682 17382
rect 11738 17380 11744 17382
rect 11436 17371 11744 17380
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11900 17218 11928 17614
rect 11992 17338 12020 17614
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11808 17202 11928 17218
rect 11796 17196 11928 17202
rect 11848 17190 11928 17196
rect 11796 17138 11848 17144
rect 11436 16348 11744 16357
rect 11436 16346 11442 16348
rect 11498 16346 11522 16348
rect 11578 16346 11602 16348
rect 11658 16346 11682 16348
rect 11738 16346 11744 16348
rect 11498 16294 11500 16346
rect 11680 16294 11682 16346
rect 11436 16292 11442 16294
rect 11498 16292 11522 16294
rect 11578 16292 11602 16294
rect 11658 16292 11682 16294
rect 11738 16292 11744 16294
rect 11436 16283 11744 16292
rect 11204 16000 11284 16028
rect 11152 15982 11204 15988
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 10980 15502 11008 15846
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 14958 11008 15438
rect 11072 15366 11100 15846
rect 11532 15570 11560 15846
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10888 14770 10916 14894
rect 10888 14742 11008 14770
rect 10876 14476 10928 14482
rect 10560 14436 10640 14464
rect 10796 14436 10876 14464
rect 10508 14418 10560 14424
rect 10612 14074 10640 14436
rect 10876 14418 10928 14424
rect 10980 14362 11008 14742
rect 11164 14414 11192 15302
rect 11436 15260 11744 15269
rect 11436 15258 11442 15260
rect 11498 15258 11522 15260
rect 11578 15258 11602 15260
rect 11658 15258 11682 15260
rect 11738 15258 11744 15260
rect 11498 15206 11500 15258
rect 11680 15206 11682 15258
rect 11436 15204 11442 15206
rect 11498 15204 11522 15206
rect 11578 15204 11602 15206
rect 11658 15204 11682 15206
rect 11738 15204 11744 15206
rect 11436 15195 11744 15204
rect 11242 14920 11298 14929
rect 11242 14855 11298 14864
rect 11256 14822 11284 14855
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 10796 14334 11008 14362
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9968 13274 9996 13330
rect 9784 12782 9812 13262
rect 9968 13246 10272 13274
rect 10244 13190 10272 13246
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 7760 11898 7788 12378
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8668 12300 8720 12306
rect 8720 12260 8984 12288
rect 8668 12242 8720 12248
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 8024 11688 8076 11694
rect 8128 11665 8156 12174
rect 8024 11630 8076 11636
rect 8114 11656 8170 11665
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7300 9674 7328 10066
rect 7208 8090 7236 9658
rect 7300 9646 7420 9674
rect 7286 9072 7342 9081
rect 7286 9007 7288 9016
rect 7340 9007 7342 9016
rect 7288 8978 7340 8984
rect 7300 8566 7328 8978
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7392 7993 7420 9646
rect 7484 8498 7512 11630
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11354 7604 11494
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7576 9110 7604 11290
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7668 8430 7696 11222
rect 8036 10606 8064 11630
rect 8114 11591 8170 11600
rect 8404 11558 8432 12242
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11694 8524 12038
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8300 11212 8352 11218
rect 8404 11200 8432 11494
rect 8588 11354 8616 12242
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8576 11212 8628 11218
rect 8404 11172 8576 11200
rect 8300 11154 8352 11160
rect 8576 11154 8628 11160
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 10198 7788 10406
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 8312 9722 8340 11154
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10130 8432 10950
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8496 9926 8524 11018
rect 8588 10169 8616 11154
rect 8680 10198 8708 11154
rect 8772 10810 8800 11154
rect 8956 11014 8984 12260
rect 9048 11626 9076 12378
rect 10152 12306 10180 13126
rect 10244 12306 10272 13126
rect 10428 12986 10456 13330
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10600 12912 10652 12918
rect 10598 12880 10600 12889
rect 10652 12880 10654 12889
rect 10598 12815 10654 12824
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 9508 12102 9536 12242
rect 10336 12102 10364 12242
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 9048 11082 9076 11562
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11218 9352 11494
rect 9312 11212 9364 11218
rect 9364 11172 9444 11200
rect 9312 11154 9364 11160
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8668 10192 8720 10198
rect 8574 10160 8630 10169
rect 8668 10134 8720 10140
rect 8574 10095 8630 10104
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 9042 7788 9522
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8404 9382 8432 9454
rect 8496 9450 8524 9862
rect 8588 9586 8616 10095
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 7852 9178 7880 9318
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 8106 7696 8366
rect 7576 8078 7696 8106
rect 7378 7984 7434 7993
rect 7196 7948 7248 7954
rect 7116 7908 7196 7936
rect 7012 7890 7064 7896
rect 7378 7919 7434 7928
rect 7196 7890 7248 7896
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6840 7534 6960 7562
rect 6932 7478 6960 7534
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6564 6866 6592 7278
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6274 6488 6330 6497
rect 6274 6423 6330 6432
rect 6288 6390 6316 6423
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6380 6254 6408 6802
rect 6472 6254 6500 6802
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6564 6118 6592 6802
rect 6656 6236 6684 7210
rect 6748 6934 6776 7346
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6932 6497 6960 7278
rect 7024 6866 7052 7686
rect 7208 7274 7236 7890
rect 7576 7750 7604 8078
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7668 7546 7696 7890
rect 7760 7546 7788 7890
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7208 6798 7236 7210
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6918 6488 6974 6497
rect 6918 6423 6974 6432
rect 6736 6248 6788 6254
rect 6656 6208 6736 6236
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 5092 4690 5120 4966
rect 5184 4826 5212 5306
rect 6196 5166 6224 5578
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6656 4826 6684 6208
rect 6736 6190 6788 6196
rect 6826 6216 6882 6225
rect 6826 6151 6828 6160
rect 6880 6151 6882 6160
rect 6828 6122 6880 6128
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4632 3602 4660 3674
rect 4724 3602 4752 4218
rect 5092 3602 5120 4626
rect 5184 4282 5212 4762
rect 6932 4758 6960 6423
rect 7392 5234 7420 6870
rect 7576 6798 7604 7346
rect 7852 7002 7880 7890
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 8220 6866 8248 7686
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7484 6633 7512 6666
rect 7470 6624 7526 6633
rect 7470 6559 7526 6568
rect 7484 6254 7512 6559
rect 7576 6390 7604 6734
rect 8036 6458 8064 6802
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 8312 6322 8340 7822
rect 8404 7313 8432 9318
rect 8680 8906 8708 10134
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 9518 8800 9862
rect 8864 9654 8892 10678
rect 8956 10674 8984 10950
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8772 8430 8800 9454
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8576 8288 8628 8294
rect 8864 8276 8892 9590
rect 8956 9450 8984 10610
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 10266 9352 10542
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9324 9518 9352 10202
rect 9416 9518 9444 11172
rect 9508 10606 9536 12038
rect 10046 11928 10102 11937
rect 10046 11863 10048 11872
rect 10100 11863 10102 11872
rect 10048 11834 10100 11840
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9968 11286 9996 11630
rect 10060 11286 10088 11834
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 8576 8230 8628 8236
rect 8772 8248 8892 8276
rect 8496 7750 8524 8230
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8588 7342 8616 8230
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8576 7336 8628 7342
rect 8390 7304 8446 7313
rect 8576 7278 8628 7284
rect 8390 7239 8446 7248
rect 8576 6928 8628 6934
rect 8680 6916 8708 7822
rect 8772 7698 8800 8248
rect 9140 7954 9168 9454
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 8634 9352 8978
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8864 7818 8892 7890
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9324 7698 9352 7754
rect 8772 7670 8892 7698
rect 8628 6888 8708 6916
rect 8576 6870 8628 6876
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6390 8432 6598
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8312 5370 8340 5782
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8404 5370 8432 5714
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8496 5302 8524 5714
rect 8588 5642 8616 6870
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8680 6322 8708 6598
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8864 5234 8892 7670
rect 8956 7670 9352 7698
rect 8956 7546 8984 7670
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6798 9076 7278
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 6866 9352 7142
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 6186 9168 6598
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8956 5914 8984 6122
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9416 5846 9444 9454
rect 9508 8022 9536 10542
rect 9692 9654 9720 10542
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10130 9812 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9876 9058 9904 11154
rect 10336 11082 10364 11562
rect 10612 11218 10640 12038
rect 10796 11694 10824 14334
rect 11256 14074 11284 14418
rect 11624 14346 11652 14418
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 11436 14172 11744 14181
rect 11436 14170 11442 14172
rect 11498 14170 11522 14172
rect 11578 14170 11602 14172
rect 11658 14170 11682 14172
rect 11738 14170 11744 14172
rect 11498 14118 11500 14170
rect 11680 14118 11682 14170
rect 11436 14116 11442 14118
rect 11498 14116 11522 14118
rect 11578 14116 11602 14118
rect 11658 14116 11682 14118
rect 11738 14116 11744 14118
rect 11436 14107 11744 14116
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11808 13734 11836 17138
rect 12544 17134 12572 17478
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12636 17134 12664 17274
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12624 17128 12676 17134
rect 12676 17088 12756 17116
rect 12624 17070 12676 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12096 16892 12404 16901
rect 12096 16890 12102 16892
rect 12158 16890 12182 16892
rect 12238 16890 12262 16892
rect 12318 16890 12342 16892
rect 12398 16890 12404 16892
rect 12158 16838 12160 16890
rect 12340 16838 12342 16890
rect 12096 16836 12102 16838
rect 12158 16836 12182 16838
rect 12238 16836 12262 16838
rect 12318 16836 12342 16838
rect 12398 16836 12404 16838
rect 12096 16827 12404 16836
rect 12544 16046 12572 16934
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11992 15366 12020 15914
rect 12096 15804 12404 15813
rect 12096 15802 12102 15804
rect 12158 15802 12182 15804
rect 12238 15802 12262 15804
rect 12318 15802 12342 15804
rect 12398 15802 12404 15804
rect 12158 15750 12160 15802
rect 12340 15750 12342 15802
rect 12096 15748 12102 15750
rect 12158 15748 12182 15750
rect 12238 15748 12262 15750
rect 12318 15748 12342 15750
rect 12398 15748 12404 15750
rect 12096 15739 12404 15748
rect 12636 15434 12664 15982
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 12622 14920 12678 14929
rect 12622 14855 12678 14864
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14550 11928 14758
rect 12096 14716 12404 14725
rect 12096 14714 12102 14716
rect 12158 14714 12182 14716
rect 12238 14714 12262 14716
rect 12318 14714 12342 14716
rect 12398 14714 12404 14716
rect 12158 14662 12160 14714
rect 12340 14662 12342 14714
rect 12096 14660 12102 14662
rect 12158 14660 12182 14662
rect 12238 14660 12262 14662
rect 12318 14660 12342 14662
rect 12398 14660 12404 14662
rect 12096 14651 12404 14660
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11992 14006 12020 14486
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11900 13326 11928 13806
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10130 10088 10406
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9692 9042 9904 9058
rect 10060 9042 10088 9318
rect 9680 9036 9904 9042
rect 9732 9030 9904 9036
rect 9680 8978 9732 8984
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8634 9812 8774
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 6322 9536 7754
rect 9600 6866 9628 8298
rect 9876 8090 9904 9030
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 8430 9996 8910
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7002 9720 7890
rect 9784 7410 9812 8026
rect 10152 7993 10180 9658
rect 10244 9518 10272 10542
rect 10428 10470 10456 10950
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10612 8838 10640 11154
rect 10980 10198 11008 12582
rect 11072 12442 11100 12650
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11164 12306 11192 13126
rect 11256 12306 11284 13262
rect 11436 13084 11744 13093
rect 11436 13082 11442 13084
rect 11498 13082 11522 13084
rect 11578 13082 11602 13084
rect 11658 13082 11682 13084
rect 11738 13082 11744 13084
rect 11498 13030 11500 13082
rect 11680 13030 11682 13082
rect 11436 13028 11442 13030
rect 11498 13028 11522 13030
rect 11578 13028 11602 13030
rect 11658 13028 11682 13030
rect 11738 13028 11744 13030
rect 11436 13019 11744 13028
rect 11900 12782 11928 13262
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11532 12306 11560 12718
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10796 9518 10824 9862
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 11072 9178 11100 11222
rect 11256 10130 11284 12106
rect 11436 11996 11744 12005
rect 11436 11994 11442 11996
rect 11498 11994 11522 11996
rect 11578 11994 11602 11996
rect 11658 11994 11682 11996
rect 11738 11994 11744 11996
rect 11498 11942 11500 11994
rect 11680 11942 11682 11994
rect 11436 11940 11442 11942
rect 11498 11940 11522 11942
rect 11578 11940 11602 11942
rect 11658 11940 11682 11942
rect 11738 11940 11744 11942
rect 11436 11931 11744 11940
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11164 8974 11192 10066
rect 11256 9722 11284 10066
rect 11348 10062 11376 10950
rect 11436 10908 11744 10917
rect 11436 10906 11442 10908
rect 11498 10906 11522 10908
rect 11578 10906 11602 10908
rect 11658 10906 11682 10908
rect 11738 10906 11744 10908
rect 11498 10854 11500 10906
rect 11680 10854 11682 10906
rect 11436 10852 11442 10854
rect 11498 10852 11522 10854
rect 11578 10852 11602 10854
rect 11658 10852 11682 10854
rect 11738 10852 11744 10854
rect 11436 10843 11744 10852
rect 11808 10606 11836 11630
rect 11900 11082 11928 12174
rect 11992 11665 12020 13942
rect 12636 13870 12664 14855
rect 12728 14618 12756 17088
rect 12820 16454 12848 17614
rect 13648 17202 13676 17750
rect 13818 17711 13820 17720
rect 13872 17711 13874 17720
rect 13820 17682 13872 17688
rect 14844 17678 14872 18770
rect 15304 18714 15332 18770
rect 15304 18686 15424 18714
rect 15396 18630 15424 18686
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 14922 18456 14978 18465
rect 14922 18391 14978 18400
rect 15290 18456 15346 18465
rect 15290 18391 15292 18400
rect 14936 17746 14964 18391
rect 15344 18391 15346 18400
rect 15292 18362 15344 18368
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15212 17746 15240 18090
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15304 17270 15332 18022
rect 15396 17746 15424 18566
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13004 16658 13032 16934
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12728 13802 12756 14214
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12096 13628 12404 13637
rect 12096 13626 12102 13628
rect 12158 13626 12182 13628
rect 12238 13626 12262 13628
rect 12318 13626 12342 13628
rect 12398 13626 12404 13628
rect 12158 13574 12160 13626
rect 12340 13574 12342 13626
rect 12096 13572 12102 13574
rect 12158 13572 12182 13574
rect 12238 13572 12262 13574
rect 12318 13572 12342 13574
rect 12398 13572 12404 13574
rect 12096 13563 12404 13572
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12096 12540 12404 12549
rect 12096 12538 12102 12540
rect 12158 12538 12182 12540
rect 12238 12538 12262 12540
rect 12318 12538 12342 12540
rect 12398 12538 12404 12540
rect 12158 12486 12160 12538
rect 12340 12486 12342 12538
rect 12096 12484 12102 12486
rect 12158 12484 12182 12486
rect 12238 12484 12262 12486
rect 12318 12484 12342 12486
rect 12398 12484 12404 12486
rect 12096 12475 12404 12484
rect 12452 12306 12480 12582
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12452 11898 12480 12106
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 11978 11656 12034 11665
rect 11978 11591 12034 11600
rect 12096 11452 12404 11461
rect 12096 11450 12102 11452
rect 12158 11450 12182 11452
rect 12238 11450 12262 11452
rect 12318 11450 12342 11452
rect 12398 11450 12404 11452
rect 12158 11398 12160 11450
rect 12340 11398 12342 11450
rect 12096 11396 12102 11398
rect 12158 11396 12182 11398
rect 12238 11396 12262 11398
rect 12318 11396 12342 11398
rect 12398 11396 12404 11398
rect 12096 11387 12404 11396
rect 12728 11150 12756 13738
rect 12820 13190 12848 14418
rect 12912 13870 12940 16458
rect 13188 16046 13216 17138
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15120 16726 15148 17070
rect 15212 16794 15240 17070
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 15108 16720 15160 16726
rect 15108 16662 15160 16668
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13648 14958 13676 15642
rect 14004 15428 14056 15434
rect 14004 15370 14056 15376
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12912 13530 12940 13806
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 13004 12714 13032 13194
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 13188 12434 13216 14894
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13266 14648 13322 14657
rect 13266 14583 13268 14592
rect 13320 14583 13322 14592
rect 13268 14554 13320 14560
rect 13280 13530 13308 14554
rect 13556 14550 13584 14826
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13740 14482 13768 15098
rect 14016 15026 14044 15370
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14108 14822 14136 15982
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14200 15609 14228 15642
rect 14186 15600 14242 15609
rect 14660 15570 14688 16662
rect 15304 16182 15332 17206
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15396 16028 15424 17682
rect 15488 17626 15516 19654
rect 15580 19446 15608 19926
rect 15672 19514 15700 20334
rect 15764 20074 15792 20742
rect 15856 20466 15884 20742
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 15764 20046 15884 20074
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15856 19310 15884 20046
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15764 19174 15792 19246
rect 15752 19168 15804 19174
rect 15658 19136 15714 19145
rect 15752 19110 15804 19116
rect 15658 19071 15714 19080
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15580 17785 15608 18770
rect 15566 17776 15622 17785
rect 15672 17762 15700 19071
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15764 17882 15792 18770
rect 15844 18692 15896 18698
rect 15844 18634 15896 18640
rect 15856 18222 15884 18634
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15948 18086 15976 19926
rect 16040 19922 16068 20198
rect 16592 20058 16620 20946
rect 16776 20913 16804 21286
rect 17500 20936 17552 20942
rect 16762 20904 16818 20913
rect 16684 20862 16762 20890
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16302 19952 16358 19961
rect 16028 19916 16080 19922
rect 16684 19922 16712 20862
rect 17500 20878 17552 20884
rect 16762 20839 16818 20848
rect 16946 20768 17002 20777
rect 16946 20703 17002 20712
rect 16960 20602 16988 20703
rect 17512 20602 17540 20878
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16080 19896 16302 19904
rect 16080 19876 16304 19896
rect 16028 19858 16080 19864
rect 16356 19887 16358 19896
rect 16396 19916 16448 19922
rect 16304 19858 16356 19864
rect 16396 19858 16448 19864
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16408 19718 16436 19858
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16396 19712 16448 19718
rect 16316 19660 16396 19666
rect 16316 19654 16448 19660
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16316 19638 16436 19654
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18630 16068 19246
rect 16132 18834 16160 19314
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16224 18222 16252 18702
rect 16316 18601 16344 19638
rect 16500 19530 16528 19654
rect 16408 19502 16528 19530
rect 16408 19242 16436 19502
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16500 18970 16528 19382
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16488 18624 16540 18630
rect 16302 18592 16358 18601
rect 16488 18566 16540 18572
rect 16302 18527 16358 18536
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 15936 18080 15988 18086
rect 16316 18057 16344 18090
rect 15936 18022 15988 18028
rect 16302 18048 16358 18057
rect 16302 17983 16358 17992
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 15672 17734 15884 17762
rect 15566 17711 15622 17720
rect 15488 17610 15608 17626
rect 15488 17604 15620 17610
rect 15488 17598 15568 17604
rect 15568 17546 15620 17552
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17202 15700 17478
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15476 16992 15528 16998
rect 15764 16980 15792 17070
rect 15528 16952 15792 16980
rect 15476 16934 15528 16940
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15580 16046 15608 16186
rect 15304 16000 15424 16028
rect 15568 16040 15620 16046
rect 14186 15535 14242 15544
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14482 14136 14758
rect 14384 14618 14412 14826
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 13740 13870 13768 14418
rect 13820 14408 13872 14414
rect 14016 14362 14044 14418
rect 13872 14356 14044 14362
rect 13820 14350 14044 14356
rect 13832 14334 14044 14350
rect 14016 14006 14044 14334
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 13394 13308 13466
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13464 12646 13492 13806
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13556 12850 13584 13126
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13096 12406 13216 12434
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 10130 11744 10406
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11716 10010 11744 10066
rect 11716 9982 11836 10010
rect 11436 9820 11744 9829
rect 11436 9818 11442 9820
rect 11498 9818 11522 9820
rect 11578 9818 11602 9820
rect 11658 9818 11682 9820
rect 11738 9818 11744 9820
rect 11498 9766 11500 9818
rect 11680 9766 11682 9818
rect 11436 9764 11442 9766
rect 11498 9764 11522 9766
rect 11578 9764 11602 9766
rect 11658 9764 11682 9766
rect 11738 9764 11744 9766
rect 11436 9755 11744 9764
rect 11244 9716 11296 9722
rect 11808 9704 11836 9982
rect 11244 9658 11296 9664
rect 11716 9676 11836 9704
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 9110 11652 9318
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11716 9042 11744 9676
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10612 8362 10640 8774
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 9862 7984 9918 7993
rect 9862 7919 9864 7928
rect 9916 7919 9918 7928
rect 10138 7984 10194 7993
rect 10138 7919 10194 7928
rect 10598 7984 10654 7993
rect 10980 7954 11008 8230
rect 10598 7919 10654 7928
rect 10968 7948 11020 7954
rect 9864 7890 9916 7896
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10322 7848 10378 7857
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9784 6322 9812 7142
rect 9864 6452 9916 6458
rect 9968 6440 9996 7822
rect 10322 7783 10378 7792
rect 10336 7478 10364 7783
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10336 7342 10364 7414
rect 10612 7342 10640 7919
rect 10968 7890 11020 7896
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9916 6412 9996 6440
rect 9864 6394 9916 6400
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9588 5772 9640 5778
rect 9640 5732 9720 5760
rect 9588 5714 9640 5720
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 7392 4826 7420 5170
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5368 3738 5396 4014
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5828 3738 5856 3946
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 6182 3632 6238 3641
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5632 3596 5684 3602
rect 6288 3602 6316 4422
rect 6828 4276 6880 4282
rect 6932 4264 6960 4694
rect 6880 4236 6960 4264
rect 6828 4218 6880 4224
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6182 3567 6184 3576
rect 5632 3538 5684 3544
rect 6236 3567 6238 3576
rect 6276 3596 6328 3602
rect 6184 3538 6236 3544
rect 6276 3538 6328 3544
rect 4724 3398 4752 3538
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 5644 2990 5672 3538
rect 6656 3194 6684 4014
rect 6932 3602 6960 4236
rect 7392 3738 7420 4762
rect 7852 4690 7880 5034
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7668 3602 7696 4558
rect 7852 4282 7880 4626
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 8220 3602 8248 4694
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3738 8616 3878
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8680 3670 8708 4014
rect 8668 3664 8720 3670
rect 8666 3632 8668 3641
rect 8720 3632 8722 3641
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8484 3596 8536 3602
rect 8666 3567 8722 3576
rect 8484 3538 8536 3544
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 7116 2990 7144 3334
rect 7576 3194 7604 3538
rect 7668 3398 7696 3538
rect 8220 3466 8248 3538
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7656 3392 7708 3398
rect 8312 3346 8340 3538
rect 8496 3398 8524 3538
rect 8668 3528 8720 3534
rect 8772 3516 8800 4218
rect 8944 3528 8996 3534
rect 8720 3488 8944 3516
rect 8668 3470 8720 3476
rect 8944 3470 8996 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 7656 3334 7708 3340
rect 8220 3318 8340 3346
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8220 3194 8248 3318
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 9324 1426 9352 2246
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 9416 882 9444 3470
rect 9692 3058 9720 5732
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 3194 9812 3538
rect 9876 3482 9904 5034
rect 9968 4434 9996 5578
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4554 10088 5102
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9968 4406 10088 4434
rect 10060 4010 10088 4406
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9876 3466 9996 3482
rect 9876 3460 10008 3466
rect 9876 3454 9956 3460
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9876 2990 9904 3454
rect 9956 3402 10008 3408
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9508 1902 9536 2450
rect 9968 2446 9996 3062
rect 10060 2922 10088 3946
rect 10244 3534 10272 6938
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6662 10364 6734
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6458 10364 6598
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10428 6186 10456 7142
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10428 4826 10456 5102
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 2990 10272 3470
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 2106 9812 2246
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 9496 1896 9548 1902
rect 9496 1838 9548 1844
rect 9968 1562 9996 2382
rect 10244 2310 10272 2450
rect 10428 2446 10456 3538
rect 10704 2825 10732 7414
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10796 7002 10824 7278
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 11072 6866 11100 7210
rect 11164 7188 11192 8774
rect 11256 7886 11284 8978
rect 11716 8838 11744 8978
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11436 8732 11744 8741
rect 11436 8730 11442 8732
rect 11498 8730 11522 8732
rect 11578 8730 11602 8732
rect 11658 8730 11682 8732
rect 11738 8730 11744 8732
rect 11498 8678 11500 8730
rect 11680 8678 11682 8730
rect 11436 8676 11442 8678
rect 11498 8676 11522 8678
rect 11578 8676 11602 8678
rect 11658 8676 11682 8678
rect 11738 8676 11744 8678
rect 11436 8667 11744 8676
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11624 8022 11652 8570
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11348 7342 11376 7958
rect 11436 7644 11744 7653
rect 11436 7642 11442 7644
rect 11498 7642 11522 7644
rect 11578 7642 11602 7644
rect 11658 7642 11682 7644
rect 11738 7642 11744 7644
rect 11498 7590 11500 7642
rect 11680 7590 11682 7642
rect 11436 7588 11442 7590
rect 11498 7588 11522 7590
rect 11578 7588 11602 7590
rect 11658 7588 11682 7590
rect 11738 7588 11744 7590
rect 11436 7579 11744 7588
rect 11808 7426 11836 9386
rect 11900 9110 11928 11018
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11992 9602 12020 10474
rect 12176 10470 12204 10542
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12096 10364 12404 10373
rect 12096 10362 12102 10364
rect 12158 10362 12182 10364
rect 12238 10362 12262 10364
rect 12318 10362 12342 10364
rect 12398 10362 12404 10364
rect 12158 10310 12160 10362
rect 12340 10310 12342 10362
rect 12096 10308 12102 10310
rect 12158 10308 12182 10310
rect 12238 10308 12262 10310
rect 12318 10308 12342 10310
rect 12398 10308 12404 10310
rect 12096 10299 12404 10308
rect 12452 10198 12480 10474
rect 12072 10192 12124 10198
rect 12070 10160 12072 10169
rect 12440 10192 12492 10198
rect 12124 10160 12126 10169
rect 12440 10134 12492 10140
rect 12070 10095 12126 10104
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12360 10033 12388 10066
rect 12346 10024 12402 10033
rect 12346 9959 12402 9968
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9738 12480 9862
rect 12360 9722 12480 9738
rect 12348 9716 12480 9722
rect 12400 9710 12480 9716
rect 12348 9658 12400 9664
rect 11992 9574 12112 9602
rect 12084 9518 12112 9574
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11992 9178 12020 9454
rect 12096 9276 12404 9285
rect 12096 9274 12102 9276
rect 12158 9274 12182 9276
rect 12238 9274 12262 9276
rect 12318 9274 12342 9276
rect 12398 9274 12404 9276
rect 12158 9222 12160 9274
rect 12340 9222 12342 9274
rect 12096 9220 12102 9222
rect 12158 9220 12182 9222
rect 12238 9220 12262 9222
rect 12318 9220 12342 9222
rect 12398 9220 12404 9222
rect 12096 9211 12404 9220
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11888 9104 11940 9110
rect 11886 9072 11888 9081
rect 11940 9072 11942 9081
rect 11886 9007 11942 9016
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12084 8922 12112 8978
rect 12544 8974 12572 10542
rect 12636 10130 12664 10746
rect 12820 10606 12848 11018
rect 13004 11014 13032 11630
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13004 10606 13032 10950
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12728 9722 12756 10474
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 13096 9178 13124 12406
rect 13464 12238 13492 12582
rect 13740 12442 13768 13806
rect 14016 13530 14044 13806
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13924 13410 13952 13466
rect 13924 13382 14044 13410
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13832 11898 13860 12650
rect 13924 12102 13952 13262
rect 14016 12186 14044 13382
rect 14108 12782 14136 14418
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 13870 14228 14214
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14200 12374 14228 13806
rect 14568 12986 14596 14418
rect 14660 13394 14688 15506
rect 15304 15162 15332 16000
rect 15568 15982 15620 15988
rect 15672 15910 15700 16526
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15396 15162 15424 15438
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15212 13802 15240 14486
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15212 13462 15240 13738
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14016 12158 14228 12186
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13556 11082 13584 11630
rect 13648 11354 13676 11766
rect 14016 11558 14044 12038
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14108 11393 14136 11630
rect 14094 11384 14150 11393
rect 13636 11348 13688 11354
rect 14094 11319 14150 11328
rect 13636 11290 13688 11296
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13188 9674 13216 11018
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10266 13584 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13188 9646 13400 9674
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12806 9072 12862 9081
rect 12806 9007 12862 9016
rect 11992 8894 12112 8922
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12716 8900 12768 8906
rect 11992 8430 12020 8894
rect 12716 8842 12768 8848
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11992 7954 12020 8366
rect 12096 8188 12404 8197
rect 12096 8186 12102 8188
rect 12158 8186 12182 8188
rect 12238 8186 12262 8188
rect 12318 8186 12342 8188
rect 12398 8186 12404 8188
rect 12158 8134 12160 8186
rect 12340 8134 12342 8186
rect 12096 8132 12102 8134
rect 12158 8132 12182 8134
rect 12238 8132 12262 8134
rect 12318 8132 12342 8134
rect 12398 8132 12404 8134
rect 12096 8123 12404 8132
rect 12728 7954 12756 8842
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 11716 7398 11836 7426
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11164 7160 11376 7188
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10980 5817 11008 6802
rect 10966 5808 11022 5817
rect 10888 5766 10966 5794
rect 10888 3194 10916 5766
rect 10966 5743 11022 5752
rect 11072 4690 11100 6802
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11256 6322 11284 6666
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 5370 11192 5510
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11256 4826 11284 6258
rect 11348 5760 11376 7160
rect 11624 6934 11652 7210
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11716 6746 11744 7398
rect 11796 7336 11848 7342
rect 11794 7304 11796 7313
rect 11888 7336 11940 7342
rect 11848 7304 11850 7313
rect 11888 7278 11940 7284
rect 11794 7239 11850 7248
rect 11900 7002 11928 7278
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11992 6866 12020 7890
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12096 7100 12404 7109
rect 12096 7098 12102 7100
rect 12158 7098 12182 7100
rect 12238 7098 12262 7100
rect 12318 7098 12342 7100
rect 12398 7098 12404 7100
rect 12158 7046 12160 7098
rect 12340 7046 12342 7098
rect 12096 7044 12102 7046
rect 12158 7044 12182 7046
rect 12238 7044 12262 7046
rect 12318 7044 12342 7046
rect 12398 7044 12404 7046
rect 12096 7035 12404 7044
rect 12544 6866 12572 7686
rect 12728 6866 12756 7890
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 11716 6718 11836 6746
rect 11436 6556 11744 6565
rect 11436 6554 11442 6556
rect 11498 6554 11522 6556
rect 11578 6554 11602 6556
rect 11658 6554 11682 6556
rect 11738 6554 11744 6556
rect 11498 6502 11500 6554
rect 11680 6502 11682 6554
rect 11436 6500 11442 6502
rect 11498 6500 11522 6502
rect 11578 6500 11602 6502
rect 11658 6500 11682 6502
rect 11738 6500 11744 6502
rect 11436 6491 11744 6500
rect 11808 6338 11836 6718
rect 11624 6310 11836 6338
rect 11520 5772 11572 5778
rect 11348 5732 11520 5760
rect 11520 5714 11572 5720
rect 11624 5642 11652 6310
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11716 5914 11744 6190
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11436 5468 11744 5477
rect 11436 5466 11442 5468
rect 11498 5466 11522 5468
rect 11578 5466 11602 5468
rect 11658 5466 11682 5468
rect 11738 5466 11744 5468
rect 11498 5414 11500 5466
rect 11680 5414 11682 5466
rect 11436 5412 11442 5414
rect 11498 5412 11522 5414
rect 11578 5412 11602 5414
rect 11658 5412 11682 5414
rect 11738 5412 11744 5414
rect 11436 5403 11744 5412
rect 11808 5370 11836 5782
rect 11900 5778 11928 6054
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11072 4078 11100 4626
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3602 11008 3878
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11072 3482 11100 3674
rect 11164 3482 11192 4626
rect 11436 4380 11744 4389
rect 11436 4378 11442 4380
rect 11498 4378 11522 4380
rect 11578 4378 11602 4380
rect 11658 4378 11682 4380
rect 11738 4378 11744 4380
rect 11498 4326 11500 4378
rect 11680 4326 11682 4378
rect 11436 4324 11442 4326
rect 11498 4324 11522 4326
rect 11578 4324 11602 4326
rect 11658 4324 11682 4326
rect 11738 4324 11744 4326
rect 11436 4315 11744 4324
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11072 3454 11192 3482
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11072 3058 11100 3454
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2984 11020 2990
rect 11164 2938 11192 3130
rect 11020 2932 11192 2938
rect 10968 2926 11192 2932
rect 10980 2910 11192 2926
rect 10876 2848 10928 2854
rect 10690 2816 10746 2825
rect 10876 2790 10928 2796
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10690 2751 10746 2760
rect 10704 2582 10732 2751
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10888 2514 10916 2790
rect 10980 2514 11008 2790
rect 11164 2582 11192 2910
rect 11256 2650 11284 4014
rect 11436 3292 11744 3301
rect 11436 3290 11442 3292
rect 11498 3290 11522 3292
rect 11578 3290 11602 3292
rect 11658 3290 11682 3292
rect 11738 3290 11744 3292
rect 11498 3238 11500 3290
rect 11680 3238 11682 3290
rect 11436 3236 11442 3238
rect 11498 3236 11522 3238
rect 11578 3236 11602 3238
rect 11658 3236 11682 3238
rect 11738 3236 11744 3238
rect 11436 3227 11744 3236
rect 11900 3194 11928 5578
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11440 2774 11468 3130
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11520 2848 11572 2854
rect 11348 2746 11468 2774
rect 11518 2816 11520 2825
rect 11572 2816 11574 2825
rect 11518 2751 11574 2760
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 1766 10272 2246
rect 10232 1760 10284 1766
rect 10232 1702 10284 1708
rect 9956 1556 10008 1562
rect 9956 1498 10008 1504
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9600 1018 9628 1362
rect 9588 1012 9640 1018
rect 9588 954 9640 960
rect 9404 876 9456 882
rect 9404 818 9456 824
rect 9968 814 9996 1498
rect 10244 950 10272 1702
rect 10232 944 10284 950
rect 10232 886 10284 892
rect 10704 814 10732 2314
rect 10888 2292 10916 2450
rect 11152 2304 11204 2310
rect 10888 2264 11152 2292
rect 11152 2246 11204 2252
rect 11348 2038 11376 2746
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11624 2310 11652 2450
rect 11704 2440 11756 2446
rect 11702 2408 11704 2417
rect 11756 2408 11758 2417
rect 11702 2343 11758 2352
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11436 2204 11744 2213
rect 11436 2202 11442 2204
rect 11498 2202 11522 2204
rect 11578 2202 11602 2204
rect 11658 2202 11682 2204
rect 11738 2202 11744 2204
rect 11498 2150 11500 2202
rect 11680 2150 11682 2202
rect 11436 2148 11442 2150
rect 11498 2148 11522 2150
rect 11578 2148 11602 2150
rect 11658 2148 11682 2150
rect 11738 2148 11744 2150
rect 11436 2139 11744 2148
rect 11808 2106 11836 2926
rect 11992 2854 12020 6190
rect 12820 6118 12848 9007
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 12900 7948 12952 7954
rect 13176 7948 13228 7954
rect 12900 7890 12952 7896
rect 13096 7908 13176 7936
rect 12912 6866 12940 7890
rect 13096 7177 13124 7908
rect 13176 7890 13228 7896
rect 13280 7818 13308 7958
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13280 7478 13308 7754
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13082 7168 13138 7177
rect 13082 7103 13138 7112
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 6390 12940 6802
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 13096 6225 13124 7103
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13082 6216 13138 6225
rect 13082 6151 13138 6160
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12096 6012 12404 6021
rect 12096 6010 12102 6012
rect 12158 6010 12182 6012
rect 12238 6010 12262 6012
rect 12318 6010 12342 6012
rect 12398 6010 12404 6012
rect 12158 5958 12160 6010
rect 12340 5958 12342 6010
rect 12096 5956 12102 5958
rect 12158 5956 12182 5958
rect 12238 5956 12262 5958
rect 12318 5956 12342 5958
rect 12398 5956 12404 5958
rect 12096 5947 12404 5956
rect 12162 5808 12218 5817
rect 12162 5743 12164 5752
rect 12216 5743 12218 5752
rect 12164 5714 12216 5720
rect 12820 5642 12848 6054
rect 12898 5672 12954 5681
rect 12808 5636 12860 5642
rect 12898 5607 12954 5616
rect 12808 5578 12860 5584
rect 12820 5098 12848 5578
rect 12912 5574 12940 5607
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12912 5166 12940 5510
rect 13096 5166 13124 6054
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12096 4924 12404 4933
rect 12096 4922 12102 4924
rect 12158 4922 12182 4924
rect 12238 4922 12262 4924
rect 12318 4922 12342 4924
rect 12398 4922 12404 4924
rect 12158 4870 12160 4922
rect 12340 4870 12342 4922
rect 12096 4868 12102 4870
rect 12158 4868 12182 4870
rect 12238 4868 12262 4870
rect 12318 4868 12342 4870
rect 12398 4868 12404 4870
rect 12096 4859 12404 4868
rect 13096 4282 13124 5102
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12096 3836 12404 3845
rect 12096 3834 12102 3836
rect 12158 3834 12182 3836
rect 12238 3834 12262 3836
rect 12318 3834 12342 3836
rect 12398 3834 12404 3836
rect 12158 3782 12160 3834
rect 12340 3782 12342 3834
rect 12096 3780 12102 3782
rect 12158 3780 12182 3782
rect 12238 3780 12262 3782
rect 12318 3780 12342 3782
rect 12398 3780 12404 3782
rect 12096 3771 12404 3780
rect 13188 2990 13216 6598
rect 13280 5914 13308 6802
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13372 5658 13400 9646
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 7954 13584 9318
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13464 7274 13492 7890
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13464 6746 13492 7210
rect 13556 6934 13584 7890
rect 13648 7342 13676 10202
rect 13740 9042 13768 10474
rect 14016 10266 14044 10542
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13740 7546 13768 7686
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13648 6866 13676 7278
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13740 7002 13768 7210
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13832 6866 13860 7142
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13544 6792 13596 6798
rect 13464 6740 13544 6746
rect 13464 6734 13596 6740
rect 13464 6718 13584 6734
rect 13924 6730 13952 7686
rect 14016 7546 14044 7822
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5778 13768 6054
rect 14200 5817 14228 12158
rect 14292 11898 14320 12242
rect 14660 12238 14688 12582
rect 14752 12442 14780 13126
rect 14936 12986 14964 13330
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14292 9586 14320 11834
rect 15212 11762 15240 13398
rect 15396 12850 15424 14962
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 12986 15516 13670
rect 15580 13530 15608 15302
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15396 12646 15424 12786
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15488 12306 15516 12922
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 14568 10130 14596 10406
rect 15028 10198 15056 10406
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 15212 9722 15240 10542
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 14384 9110 14412 9386
rect 14476 9178 14504 9454
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14844 9110 14872 9318
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 15200 9036 15252 9042
rect 15304 9024 15332 12242
rect 15488 11762 15516 12242
rect 15672 12186 15700 15846
rect 15856 15094 15884 17734
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16224 16658 16252 17614
rect 16316 16794 16344 17818
rect 16408 17746 16436 18226
rect 16500 18086 16528 18566
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16500 17610 16528 18022
rect 16592 17746 16620 19722
rect 16684 19145 16712 19858
rect 16776 19514 16804 20334
rect 16960 19922 16988 20538
rect 17604 20398 17632 21354
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 17684 21072 17736 21078
rect 17684 21014 17736 21020
rect 17696 20777 17724 21014
rect 17788 21010 17816 21286
rect 18524 21010 18552 21286
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 17868 20800 17920 20806
rect 17682 20768 17738 20777
rect 17868 20742 17920 20748
rect 17682 20703 17738 20712
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 17052 19802 17080 20198
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17132 19984 17184 19990
rect 17592 19984 17644 19990
rect 17132 19926 17184 19932
rect 17590 19952 17592 19961
rect 17644 19952 17646 19961
rect 16960 19774 17080 19802
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16776 19310 16804 19450
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16856 19304 16908 19310
rect 16960 19281 16988 19774
rect 17144 19310 17172 19926
rect 17590 19887 17646 19896
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17604 19514 17632 19722
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17236 19310 17264 19450
rect 17132 19304 17184 19310
rect 16856 19246 16908 19252
rect 16946 19272 17002 19281
rect 16670 19136 16726 19145
rect 16670 19071 16726 19080
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 17814 16712 18566
rect 16776 18034 16804 19246
rect 16868 18358 16896 19246
rect 17130 19272 17132 19281
rect 17224 19304 17276 19310
rect 17184 19272 17186 19281
rect 16946 19207 16948 19216
rect 17000 19207 17002 19216
rect 17040 19236 17092 19242
rect 16948 19178 17000 19184
rect 17224 19246 17276 19252
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17130 19207 17186 19216
rect 17040 19178 17092 19184
rect 17052 19145 17080 19178
rect 17038 19136 17094 19145
rect 17038 19071 17094 19080
rect 17038 19000 17094 19009
rect 17236 18952 17264 19246
rect 17604 18970 17632 19246
rect 17038 18935 17094 18944
rect 16946 18864 17002 18873
rect 17052 18834 17080 18935
rect 17144 18924 17264 18952
rect 17316 18964 17368 18970
rect 16946 18799 16948 18808
rect 17000 18799 17002 18808
rect 17040 18828 17092 18834
rect 16948 18770 17000 18776
rect 17040 18770 17092 18776
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16776 18006 16896 18034
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16776 17610 16804 17682
rect 16868 17678 16896 18006
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16670 17368 16726 17377
rect 16670 17303 16672 17312
rect 16724 17303 16726 17312
rect 16672 17274 16724 17280
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16224 16250 16252 16594
rect 16316 16454 16344 16730
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15706 16160 16050
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15764 14346 15792 14894
rect 15752 14340 15804 14346
rect 15804 14300 15884 14328
rect 15752 14282 15804 14288
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15764 13530 15792 13806
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15856 12782 15884 14300
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 13462 15976 13670
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 16040 13258 16068 15506
rect 16316 15042 16344 16390
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16408 15162 16436 15982
rect 16592 15162 16620 16934
rect 16776 16590 16804 17546
rect 16960 17338 16988 18770
rect 17052 17921 17080 18770
rect 17144 18306 17172 18924
rect 17316 18906 17368 18912
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17236 18465 17264 18770
rect 17328 18698 17356 18906
rect 17696 18834 17724 19994
rect 17788 18970 17816 20198
rect 17880 19310 17908 20742
rect 17972 20058 18000 20946
rect 18248 20913 18276 20946
rect 18234 20904 18290 20913
rect 18234 20839 18290 20848
rect 18616 20618 18644 21422
rect 19432 21422 19484 21428
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 21548 21480 21600 21486
rect 21548 21422 21600 21428
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 19246 21383 19248 21392
rect 19300 21383 19302 21392
rect 19248 21354 19300 21360
rect 19260 21146 19288 21354
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18524 20590 18644 20618
rect 18052 20528 18104 20534
rect 18050 20496 18052 20505
rect 18104 20496 18106 20505
rect 18050 20431 18106 20440
rect 18236 20392 18288 20398
rect 18328 20392 18380 20398
rect 18236 20334 18288 20340
rect 18326 20360 18328 20369
rect 18420 20392 18472 20398
rect 18380 20360 18382 20369
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 18064 18834 18092 19450
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17408 18624 17460 18630
rect 17512 18601 17540 18702
rect 17696 18698 17724 18770
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17408 18566 17460 18572
rect 17498 18592 17554 18601
rect 17222 18456 17278 18465
rect 17420 18426 17448 18566
rect 17498 18527 17554 18536
rect 17498 18456 17554 18465
rect 17222 18391 17278 18400
rect 17408 18420 17460 18426
rect 17498 18391 17554 18400
rect 17408 18362 17460 18368
rect 17144 18290 17448 18306
rect 17512 18290 17540 18391
rect 17144 18284 17460 18290
rect 17144 18278 17408 18284
rect 17408 18226 17460 18232
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17038 17912 17094 17921
rect 17038 17847 17094 17856
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16960 17134 16988 17274
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16960 16726 16988 17070
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 17052 16590 17080 17847
rect 17144 17785 17172 18158
rect 17130 17776 17186 17785
rect 17130 17711 17186 17720
rect 17316 17740 17368 17746
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17144 16454 17172 17711
rect 17316 17682 17368 17688
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17236 16794 17264 16934
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 15366 16712 16050
rect 16868 15570 16896 16390
rect 17144 15910 17172 16390
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16316 15014 16436 15042
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 16132 13802 16160 14826
rect 16210 14512 16266 14521
rect 16210 14447 16212 14456
rect 16264 14447 16266 14456
rect 16304 14476 16356 14482
rect 16212 14418 16264 14424
rect 16304 14418 16356 14424
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 13870 16252 14214
rect 16316 14074 16344 14418
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16408 13954 16436 15014
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16316 13926 16436 13954
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 15934 12880 15990 12889
rect 15934 12815 15990 12824
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15764 12186 15792 12242
rect 15672 12158 15792 12186
rect 15672 11898 15700 12158
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15764 11694 15792 12038
rect 15948 11694 15976 12815
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 11218 15424 11494
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15396 10674 15424 11154
rect 15856 10810 15884 11154
rect 16040 11082 16068 13194
rect 16316 12889 16344 13926
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16408 13394 16436 13670
rect 16500 13394 16528 14962
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16500 12986 16528 13330
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16302 12880 16358 12889
rect 16302 12815 16358 12824
rect 16486 12880 16542 12889
rect 16486 12815 16542 12824
rect 16500 12782 16528 12815
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16408 12434 16436 12718
rect 16408 12406 16528 12434
rect 16500 12170 16528 12406
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16132 11218 16160 12038
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16408 10674 16436 12038
rect 16500 10674 16528 12106
rect 16592 11694 16620 15098
rect 16960 15094 16988 15506
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16948 14952 17000 14958
rect 17144 14940 17172 15846
rect 17000 14912 17172 14940
rect 17224 14952 17276 14958
rect 16948 14894 17000 14900
rect 17224 14894 17276 14900
rect 16868 14414 16896 14894
rect 16960 14822 16988 14894
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16776 13394 16804 14350
rect 16960 14346 16988 14758
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16868 13530 16896 13738
rect 17052 13530 17080 13806
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17236 13462 17264 14894
rect 17328 14618 17356 17682
rect 17420 17320 17448 18226
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17420 17292 17540 17320
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17420 16794 17448 17138
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17512 16658 17540 17292
rect 17604 16998 17632 17614
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17604 16794 17632 16934
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16684 12782 16712 13126
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16684 12306 16712 12582
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 15252 8996 15332 9024
rect 15396 9908 15424 10610
rect 15476 9920 15528 9926
rect 15396 9880 15476 9908
rect 15200 8978 15252 8984
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14568 8090 14596 8570
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14476 7546 14504 7822
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14568 7342 14596 8026
rect 14660 7426 14688 8978
rect 15396 8906 15424 9880
rect 15476 9862 15528 9868
rect 15948 9450 15976 10610
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16040 10130 16068 10542
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16316 10169 16344 10474
rect 16302 10160 16358 10169
rect 16028 10124 16080 10130
rect 16302 10095 16358 10104
rect 16028 10066 16080 10072
rect 16040 10033 16068 10066
rect 16026 10024 16082 10033
rect 16026 9959 16082 9968
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16224 9518 16252 9862
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15566 9072 15622 9081
rect 15476 9036 15528 9042
rect 15566 9007 15568 9016
rect 15476 8978 15528 8984
rect 15620 9007 15622 9016
rect 15568 8978 15620 8984
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15488 8838 15516 8978
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 8566 15516 8774
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7546 14780 7686
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14660 7398 14780 7426
rect 14844 7410 14872 8230
rect 15304 7954 15332 8230
rect 15856 8022 15884 9318
rect 15948 8974 15976 9386
rect 16132 9178 16160 9454
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8566 15976 8910
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15108 7948 15160 7954
rect 15028 7908 15108 7936
rect 14922 7576 14978 7585
rect 14922 7511 14978 7520
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14002 5808 14058 5817
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13728 5772 13780 5778
rect 14186 5808 14242 5817
rect 14002 5743 14004 5752
rect 13728 5714 13780 5720
rect 14056 5743 14058 5752
rect 14096 5772 14148 5778
rect 14004 5714 14056 5720
rect 14186 5743 14242 5752
rect 14096 5714 14148 5720
rect 13556 5681 13584 5714
rect 13542 5672 13598 5681
rect 13280 5630 13492 5658
rect 13280 5234 13308 5630
rect 13464 5574 13492 5630
rect 13542 5607 13598 5616
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13648 5522 13676 5714
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13372 4690 13400 5510
rect 13648 5494 13768 5522
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13648 5234 13676 5306
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13740 5148 13768 5494
rect 13832 5273 13860 5646
rect 14108 5642 14136 5714
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 13818 5264 13874 5273
rect 13818 5199 13874 5208
rect 13820 5160 13872 5166
rect 13740 5120 13820 5148
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13556 4486 13584 5102
rect 13740 4826 13768 5120
rect 13820 5102 13872 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13832 4078 13860 4966
rect 14292 4570 14320 6802
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14384 5302 14412 5714
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14476 5166 14504 5714
rect 14568 5234 14596 5714
rect 14648 5704 14700 5710
rect 14752 5681 14780 7398
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14936 7342 14964 7511
rect 15028 7449 15056 7908
rect 15292 7948 15344 7954
rect 15108 7890 15160 7896
rect 15212 7908 15292 7936
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15120 7478 15148 7686
rect 15108 7472 15160 7478
rect 15014 7440 15070 7449
rect 15108 7414 15160 7420
rect 15014 7375 15070 7384
rect 15028 7342 15056 7375
rect 15212 7342 15240 7908
rect 15292 7890 15344 7896
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15384 7880 15436 7886
rect 15580 7857 15608 7890
rect 15384 7822 15436 7828
rect 15566 7848 15622 7857
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15396 7002 15424 7822
rect 15566 7783 15622 7792
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15488 7002 15516 7686
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15580 7342 15608 7414
rect 15672 7342 15700 7686
rect 15856 7342 15884 7958
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15568 7200 15620 7206
rect 15660 7200 15712 7206
rect 15568 7142 15620 7148
rect 15658 7168 15660 7177
rect 15752 7200 15804 7206
rect 15712 7168 15714 7177
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15580 6934 15608 7142
rect 15948 7188 15976 8502
rect 15752 7142 15804 7148
rect 15856 7160 15976 7188
rect 15658 7103 15714 7112
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 5778 14872 6190
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14648 5646 14700 5652
rect 14738 5672 14794 5681
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14660 5166 14688 5646
rect 14738 5607 14794 5616
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14936 5166 14964 5510
rect 15028 5370 15056 6802
rect 15488 6458 15516 6802
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15672 5914 15700 6802
rect 15764 6798 15792 7142
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15764 5817 15792 5850
rect 15750 5808 15806 5817
rect 15750 5743 15806 5752
rect 15198 5672 15254 5681
rect 15198 5607 15254 5616
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15212 5166 15240 5607
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 14660 4826 14688 5102
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14016 4542 14320 4570
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 14016 4010 14044 4542
rect 14752 4282 14780 5102
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 4690 14964 4966
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14004 4004 14056 4010
rect 14004 3946 14056 3952
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 11980 2848 12032 2854
rect 11886 2816 11942 2825
rect 11980 2790 12032 2796
rect 11886 2751 11942 2760
rect 11900 2496 11928 2751
rect 11992 2632 12020 2790
rect 12096 2748 12404 2757
rect 12096 2746 12102 2748
rect 12158 2746 12182 2748
rect 12238 2746 12262 2748
rect 12318 2746 12342 2748
rect 12398 2746 12404 2748
rect 12158 2694 12160 2746
rect 12340 2694 12342 2746
rect 12096 2692 12102 2694
rect 12158 2692 12182 2694
rect 12238 2692 12262 2694
rect 12318 2692 12342 2694
rect 12398 2692 12404 2694
rect 12096 2683 12404 2692
rect 12452 2632 12480 2858
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 11992 2604 12204 2632
rect 11900 2468 12020 2496
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 11428 1896 11480 1902
rect 11428 1838 11480 1844
rect 11256 1426 11284 1838
rect 11440 1578 11468 1838
rect 11624 1834 11652 1974
rect 11796 1964 11848 1970
rect 11796 1906 11848 1912
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 11716 1578 11744 1838
rect 11808 1766 11836 1906
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11440 1556 11744 1578
rect 11440 1550 11612 1556
rect 11664 1550 11744 1556
rect 11612 1498 11664 1504
rect 11900 1426 11928 2314
rect 11992 1970 12020 2468
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 11980 1964 12032 1970
rect 11980 1906 12032 1912
rect 12084 1902 12112 2382
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 12176 1834 12204 2604
rect 12360 2604 12480 2632
rect 12360 2514 12388 2604
rect 13096 2582 13124 2790
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12360 1970 12388 2450
rect 13556 1970 13584 2926
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 11980 1828 12032 1834
rect 11980 1770 12032 1776
rect 12164 1828 12216 1834
rect 12164 1770 12216 1776
rect 11992 1562 12020 1770
rect 12096 1660 12404 1669
rect 12096 1658 12102 1660
rect 12158 1658 12182 1660
rect 12238 1658 12262 1660
rect 12318 1658 12342 1660
rect 12398 1658 12404 1660
rect 12158 1606 12160 1658
rect 12340 1606 12342 1658
rect 12096 1604 12102 1606
rect 12158 1604 12182 1606
rect 12238 1604 12262 1606
rect 12318 1604 12342 1606
rect 12398 1604 12404 1606
rect 12096 1595 12404 1604
rect 11980 1556 12032 1562
rect 11980 1498 12032 1504
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11888 1420 11940 1426
rect 11888 1362 11940 1368
rect 11336 1216 11388 1222
rect 11336 1158 11388 1164
rect 11348 1018 11376 1158
rect 11436 1116 11744 1125
rect 11436 1114 11442 1116
rect 11498 1114 11522 1116
rect 11578 1114 11602 1116
rect 11658 1114 11682 1116
rect 11738 1114 11744 1116
rect 11498 1062 11500 1114
rect 11680 1062 11682 1114
rect 11436 1060 11442 1062
rect 11498 1060 11522 1062
rect 11578 1060 11602 1062
rect 11658 1060 11682 1062
rect 11738 1060 11744 1062
rect 11436 1051 11744 1060
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 11992 814 12020 1498
rect 13004 1222 13032 1838
rect 13832 1766 13860 2790
rect 14016 2514 14044 3946
rect 14384 3738 14412 4014
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 14108 2582 14136 2790
rect 14844 2582 14872 3402
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14844 1834 14872 2518
rect 14936 2106 14964 3130
rect 15028 2990 15056 5102
rect 15856 5030 15884 7160
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15764 4690 15792 4966
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15856 4214 15884 4966
rect 15948 4486 15976 5034
rect 16040 4758 16068 8842
rect 16224 8430 16252 9454
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16408 9110 16436 9386
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16396 8016 16448 8022
rect 16396 7958 16448 7964
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7585 16344 7686
rect 16302 7576 16358 7585
rect 16302 7511 16358 7520
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16132 6934 16160 7278
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16408 6866 16436 7958
rect 16592 7313 16620 11630
rect 16776 11098 16804 13330
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 12782 17080 13262
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16868 11898 16896 12242
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16684 11070 16804 11098
rect 16684 9654 16712 11070
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 10606 16804 10950
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16684 7886 16712 8298
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16578 7304 16634 7313
rect 16578 7239 16634 7248
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 6322 16344 6734
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16408 5778 16436 6802
rect 16500 6662 16528 7142
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16118 5264 16174 5273
rect 16118 5199 16174 5208
rect 16132 5166 16160 5199
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16500 4758 16528 4966
rect 16684 4758 16712 7346
rect 16776 7342 16804 10406
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 9518 16896 9862
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17144 9178 17172 9454
rect 17420 9432 17448 14282
rect 17512 14278 17540 15574
rect 17590 15056 17646 15065
rect 17590 14991 17646 15000
rect 17604 14958 17632 14991
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17512 13938 17540 14214
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17696 13190 17724 18634
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17880 18426 17908 18566
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 17882 17908 18090
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17880 16697 17908 17818
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17866 16688 17922 16697
rect 17866 16623 17922 16632
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17972 15570 18000 15642
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17788 14006 17816 14826
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 14482 17908 14758
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17972 14006 18000 15506
rect 18064 14657 18092 17206
rect 18156 16726 18184 19858
rect 18248 19514 18276 20334
rect 18420 20334 18472 20340
rect 18326 20295 18382 20304
rect 18432 20058 18460 20334
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18524 19922 18552 20590
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18512 19916 18564 19922
rect 18616 19904 18644 20470
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18892 20369 18920 20402
rect 18878 20360 18934 20369
rect 18878 20295 18934 20304
rect 18984 20058 19012 20878
rect 19210 20700 19518 20709
rect 19210 20698 19216 20700
rect 19272 20698 19296 20700
rect 19352 20698 19376 20700
rect 19432 20698 19456 20700
rect 19512 20698 19518 20700
rect 19272 20646 19274 20698
rect 19454 20646 19456 20698
rect 19210 20644 19216 20646
rect 19272 20644 19296 20646
rect 19352 20644 19376 20646
rect 19432 20644 19456 20646
rect 19512 20644 19518 20646
rect 19210 20635 19518 20644
rect 19062 20496 19118 20505
rect 19062 20431 19118 20440
rect 19076 20398 19104 20431
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19628 20346 19656 21286
rect 19720 21010 19748 21286
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19812 20398 19840 21422
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 19870 21244 20178 21253
rect 19870 21242 19876 21244
rect 19932 21242 19956 21244
rect 20012 21242 20036 21244
rect 20092 21242 20116 21244
rect 20172 21242 20178 21244
rect 19932 21190 19934 21242
rect 20114 21190 20116 21242
rect 19870 21188 19876 21190
rect 19932 21188 19956 21190
rect 20012 21188 20036 21190
rect 20092 21188 20116 21190
rect 20172 21188 20178 21190
rect 19870 21179 20178 21188
rect 19892 21140 19944 21146
rect 19892 21082 19944 21088
rect 19800 20392 19852 20398
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 19352 19922 19380 20198
rect 19444 20058 19472 20334
rect 19628 20330 19748 20346
rect 19800 20334 19852 20340
rect 19628 20324 19760 20330
rect 19628 20318 19708 20324
rect 19708 20266 19760 20272
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19628 19922 19656 20198
rect 18696 19916 18748 19922
rect 18616 19876 18696 19904
rect 18512 19858 18564 19864
rect 18696 19858 18748 19864
rect 19340 19916 19392 19922
rect 19616 19916 19668 19922
rect 19392 19876 19564 19904
rect 19340 19858 19392 19864
rect 18524 19825 18552 19858
rect 18510 19816 18566 19825
rect 18510 19751 18566 19760
rect 19062 19816 19118 19825
rect 19536 19802 19564 19876
rect 19616 19858 19668 19864
rect 19536 19774 19656 19802
rect 19062 19751 19064 19760
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18524 19009 18552 19751
rect 19116 19751 19118 19760
rect 19064 19722 19116 19728
rect 19210 19612 19518 19621
rect 19210 19610 19216 19612
rect 19272 19610 19296 19612
rect 19352 19610 19376 19612
rect 19432 19610 19456 19612
rect 19512 19610 19518 19612
rect 19272 19558 19274 19610
rect 19454 19558 19456 19610
rect 19210 19556 19216 19558
rect 19272 19556 19296 19558
rect 19352 19556 19376 19558
rect 19432 19556 19456 19558
rect 19512 19556 19518 19558
rect 19210 19547 19518 19556
rect 19628 19310 19656 19774
rect 19720 19378 19748 20266
rect 19904 20262 19932 21082
rect 20272 20602 20300 21354
rect 21560 21078 21588 21422
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20272 20398 20300 20538
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 19870 20156 20178 20165
rect 19870 20154 19876 20156
rect 19932 20154 19956 20156
rect 20012 20154 20036 20156
rect 20092 20154 20116 20156
rect 20172 20154 20178 20156
rect 19932 20102 19934 20154
rect 20114 20102 20116 20154
rect 19870 20100 19876 20102
rect 19932 20100 19956 20102
rect 20012 20100 20036 20102
rect 20092 20100 20116 20102
rect 20172 20100 20178 20102
rect 19870 20091 20178 20100
rect 20272 19446 20300 20198
rect 20350 20088 20406 20097
rect 20350 20023 20352 20032
rect 20404 20023 20406 20032
rect 20352 19994 20404 20000
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 18972 19304 19024 19310
rect 19156 19304 19208 19310
rect 18972 19246 19024 19252
rect 19154 19272 19156 19281
rect 19616 19304 19668 19310
rect 19208 19272 19210 19281
rect 18510 19000 18566 19009
rect 18510 18935 18566 18944
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 18057 18276 18226
rect 18234 18048 18290 18057
rect 18234 17983 18290 17992
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18708 16046 18736 16662
rect 18800 16658 18828 18770
rect 18984 18766 19012 19246
rect 19616 19246 19668 19252
rect 19154 19207 19210 19216
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19708 18896 19760 18902
rect 19708 18838 19760 18844
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19210 18524 19518 18533
rect 19210 18522 19216 18524
rect 19272 18522 19296 18524
rect 19352 18522 19376 18524
rect 19432 18522 19456 18524
rect 19512 18522 19518 18524
rect 19272 18470 19274 18522
rect 19454 18470 19456 18522
rect 19210 18468 19216 18470
rect 19272 18468 19296 18470
rect 19352 18468 19376 18470
rect 19432 18468 19456 18470
rect 19512 18468 19518 18470
rect 19210 18459 19518 18468
rect 18880 18148 18932 18154
rect 18880 18090 18932 18096
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18236 15972 18288 15978
rect 18236 15914 18288 15920
rect 18248 15706 18276 15914
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18050 14648 18106 14657
rect 18050 14583 18106 14592
rect 18432 14550 18460 15438
rect 18892 14890 18920 18090
rect 19628 18086 19656 18702
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19210 17436 19518 17445
rect 19210 17434 19216 17436
rect 19272 17434 19296 17436
rect 19352 17434 19376 17436
rect 19432 17434 19456 17436
rect 19512 17434 19518 17436
rect 19272 17382 19274 17434
rect 19454 17382 19456 17434
rect 19210 17380 19216 17382
rect 19272 17380 19296 17382
rect 19352 17380 19376 17382
rect 19432 17380 19456 17382
rect 19512 17380 19518 17382
rect 19210 17371 19518 17380
rect 19248 17264 19300 17270
rect 19628 17218 19656 18022
rect 19248 17206 19300 17212
rect 19064 16720 19116 16726
rect 19064 16662 19116 16668
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 18984 15638 19012 16526
rect 19076 15706 19104 16662
rect 19260 16658 19288 17206
rect 19536 17190 19656 17218
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19536 16590 19564 17190
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19210 16348 19518 16357
rect 19210 16346 19216 16348
rect 19272 16346 19296 16348
rect 19352 16346 19376 16348
rect 19432 16346 19456 16348
rect 19512 16346 19518 16348
rect 19272 16294 19274 16346
rect 19454 16294 19456 16346
rect 19210 16292 19216 16294
rect 19272 16292 19296 16294
rect 19352 16292 19376 16294
rect 19432 16292 19456 16294
rect 19512 16292 19518 16294
rect 19210 16283 19518 16292
rect 19628 16046 19656 16934
rect 19720 16250 19748 18838
rect 19812 18222 19840 19178
rect 20258 19136 20314 19145
rect 19870 19068 20178 19077
rect 20258 19071 20314 19080
rect 19870 19066 19876 19068
rect 19932 19066 19956 19068
rect 20012 19066 20036 19068
rect 20092 19066 20116 19068
rect 20172 19066 20178 19068
rect 19932 19014 19934 19066
rect 20114 19014 20116 19066
rect 19870 19012 19876 19014
rect 19932 19012 19956 19014
rect 20012 19012 20036 19014
rect 20092 19012 20116 19014
rect 20172 19012 20178 19014
rect 19870 19003 20178 19012
rect 20272 18834 20300 19071
rect 20548 18834 20576 19382
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20272 18601 20300 18770
rect 20258 18592 20314 18601
rect 20258 18527 20314 18536
rect 20074 18456 20130 18465
rect 20272 18426 20300 18527
rect 20074 18391 20130 18400
rect 20260 18420 20312 18426
rect 20088 18222 20116 18391
rect 20260 18362 20312 18368
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20444 18216 20496 18222
rect 20548 18204 20576 18770
rect 20640 18442 20668 18770
rect 20732 18601 20760 18770
rect 20718 18592 20774 18601
rect 20718 18527 20774 18536
rect 20640 18426 20760 18442
rect 20640 18420 20772 18426
rect 20640 18414 20720 18420
rect 20720 18362 20772 18368
rect 20548 18176 20760 18204
rect 20444 18158 20496 18164
rect 20088 18068 20116 18158
rect 19812 18040 20116 18068
rect 20456 18057 20484 18158
rect 20442 18048 20498 18057
rect 19812 17270 19840 18040
rect 19870 17980 20178 17989
rect 20442 17983 20498 17992
rect 19870 17978 19876 17980
rect 19932 17978 19956 17980
rect 20012 17978 20036 17980
rect 20092 17978 20116 17980
rect 20172 17978 20178 17980
rect 19932 17926 19934 17978
rect 20114 17926 20116 17978
rect 19870 17924 19876 17926
rect 19932 17924 19956 17926
rect 20012 17924 20036 17926
rect 20092 17924 20116 17926
rect 20172 17924 20178 17926
rect 19870 17915 20178 17924
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20456 17270 20484 17478
rect 20548 17270 20576 17682
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 19812 16776 19840 17070
rect 19870 16892 20178 16901
rect 19870 16890 19876 16892
rect 19932 16890 19956 16892
rect 20012 16890 20036 16892
rect 20092 16890 20116 16892
rect 20172 16890 20178 16892
rect 19932 16838 19934 16890
rect 20114 16838 20116 16890
rect 19870 16836 19876 16838
rect 19932 16836 19956 16838
rect 20012 16836 20036 16838
rect 20092 16836 20116 16838
rect 20172 16836 20178 16838
rect 19870 16827 20178 16836
rect 20456 16833 20484 17070
rect 20442 16824 20498 16833
rect 19812 16748 19932 16776
rect 20442 16759 20498 16768
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19812 16130 19840 16526
rect 19904 16522 19932 16748
rect 20166 16688 20222 16697
rect 20166 16623 20222 16632
rect 20442 16688 20498 16697
rect 20442 16623 20498 16632
rect 20180 16572 20208 16623
rect 20352 16584 20404 16590
rect 20180 16544 20352 16572
rect 20352 16526 20404 16532
rect 19892 16516 19944 16522
rect 19892 16458 19944 16464
rect 19720 16102 19840 16130
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18984 14634 19012 15574
rect 19536 15570 19564 15846
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18892 14606 19012 14634
rect 19076 14618 19104 15370
rect 19210 15260 19518 15269
rect 19210 15258 19216 15260
rect 19272 15258 19296 15260
rect 19352 15258 19376 15260
rect 19432 15258 19456 15260
rect 19512 15258 19518 15260
rect 19272 15206 19274 15258
rect 19454 15206 19456 15258
rect 19210 15204 19216 15206
rect 19272 15204 19296 15206
rect 19352 15204 19376 15206
rect 19432 15204 19456 15206
rect 19512 15204 19518 15206
rect 19210 15195 19518 15204
rect 19628 15094 19656 15438
rect 19616 15088 19668 15094
rect 19616 15030 19668 15036
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19064 14612 19116 14618
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18340 14278 18368 14418
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17696 11393 17724 11562
rect 17682 11384 17738 11393
rect 17682 11319 17738 11328
rect 17696 11150 17724 11319
rect 17788 11257 17816 13942
rect 17972 13870 18000 13942
rect 18432 13938 18460 14486
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18892 13530 18920 14606
rect 19064 14554 19116 14560
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18984 14074 19012 14418
rect 19352 14414 19380 14962
rect 19628 14958 19656 15030
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19628 14482 19656 14894
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 12374 17908 13330
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18156 12442 18184 12650
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17972 11830 18000 12174
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18064 11694 18092 11834
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17774 11248 17830 11257
rect 17774 11183 17830 11192
rect 17684 11144 17736 11150
rect 18156 11132 18184 12378
rect 18892 12306 18920 13126
rect 19076 12986 19104 14214
rect 19210 14172 19518 14181
rect 19210 14170 19216 14172
rect 19272 14170 19296 14172
rect 19352 14170 19376 14172
rect 19432 14170 19456 14172
rect 19512 14170 19518 14172
rect 19272 14118 19274 14170
rect 19454 14118 19456 14170
rect 19210 14116 19216 14118
rect 19272 14116 19296 14118
rect 19352 14116 19376 14118
rect 19432 14116 19456 14118
rect 19512 14116 19518 14118
rect 19210 14107 19518 14116
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19260 13938 19288 14010
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19720 13394 19748 16102
rect 19904 15910 19932 16458
rect 20260 15972 20312 15978
rect 20260 15914 20312 15920
rect 19892 15904 19944 15910
rect 20272 15881 20300 15914
rect 19892 15846 19944 15852
rect 20258 15872 20314 15881
rect 19870 15804 20178 15813
rect 20258 15807 20314 15816
rect 19870 15802 19876 15804
rect 19932 15802 19956 15804
rect 20012 15802 20036 15804
rect 20092 15802 20116 15804
rect 20172 15802 20178 15804
rect 19932 15750 19934 15802
rect 20114 15750 20116 15802
rect 19870 15748 19876 15750
rect 19932 15748 19956 15750
rect 20012 15748 20036 15750
rect 20092 15748 20116 15750
rect 20172 15748 20178 15750
rect 19870 15739 20178 15748
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19812 13870 19840 15506
rect 19870 14716 20178 14725
rect 19870 14714 19876 14716
rect 19932 14714 19956 14716
rect 20012 14714 20036 14716
rect 20092 14714 20116 14716
rect 20172 14714 20178 14716
rect 19932 14662 19934 14714
rect 20114 14662 20116 14714
rect 19870 14660 19876 14662
rect 19932 14660 19956 14662
rect 20012 14660 20036 14662
rect 20092 14660 20116 14662
rect 20172 14660 20178 14662
rect 19870 14651 20178 14660
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 14249 19932 14350
rect 19890 14240 19946 14249
rect 19890 14175 19946 14184
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19870 13628 20178 13637
rect 19870 13626 19876 13628
rect 19932 13626 19956 13628
rect 20012 13626 20036 13628
rect 20092 13626 20116 13628
rect 20172 13626 20178 13628
rect 19932 13574 19934 13626
rect 20114 13574 20116 13626
rect 19870 13572 19876 13574
rect 19932 13572 19956 13574
rect 20012 13572 20036 13574
rect 20092 13572 20116 13574
rect 20172 13572 20178 13574
rect 19870 13563 20178 13572
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 19982 13424 20038 13433
rect 19708 13388 19760 13394
rect 20088 13394 20116 13466
rect 19982 13359 20038 13368
rect 20076 13388 20128 13394
rect 19708 13330 19760 13336
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19210 13084 19518 13093
rect 19210 13082 19216 13084
rect 19272 13082 19296 13084
rect 19352 13082 19376 13084
rect 19432 13082 19456 13084
rect 19512 13082 19518 13084
rect 19272 13030 19274 13082
rect 19454 13030 19456 13082
rect 19210 13028 19216 13030
rect 19272 13028 19296 13030
rect 19352 13028 19376 13030
rect 19432 13028 19456 13030
rect 19512 13028 19518 13030
rect 19210 13019 19518 13028
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19076 12442 19104 12582
rect 19064 12436 19116 12442
rect 19628 12434 19656 12922
rect 19720 12782 19748 13126
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19812 12714 19840 13126
rect 19996 12782 20024 13359
rect 20076 13330 20128 13336
rect 20088 12918 20116 13330
rect 20456 13326 20484 16623
rect 20548 16572 20576 17206
rect 20640 16697 20668 17682
rect 20732 17134 20760 18176
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20718 16824 20774 16833
rect 20718 16759 20774 16768
rect 20626 16688 20682 16697
rect 20626 16623 20682 16632
rect 20628 16584 20680 16590
rect 20548 16544 20628 16572
rect 20628 16526 20680 16532
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20548 13530 20576 15506
rect 20640 15434 20668 15982
rect 20732 15706 20760 16759
rect 20824 16674 20852 20742
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20916 19922 20944 20334
rect 21560 19922 21588 21014
rect 21836 21010 21864 21286
rect 24044 21078 24072 21286
rect 24032 21072 24084 21078
rect 24032 21014 24084 21020
rect 24596 21010 24624 21286
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 22926 20904 22982 20913
rect 22926 20839 22982 20848
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 22112 19825 22140 20266
rect 22204 20058 22232 20266
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22098 19816 22154 19825
rect 22098 19751 22154 19760
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20916 18698 20944 18906
rect 21008 18834 21036 19110
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 21008 18290 21036 18566
rect 21100 18290 21128 19314
rect 21192 18290 21220 19450
rect 21284 18834 21312 19654
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21376 18714 21404 19110
rect 21836 18902 21864 19246
rect 21548 18896 21600 18902
rect 21454 18864 21510 18873
rect 21548 18838 21600 18844
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21454 18799 21510 18808
rect 21284 18686 21404 18714
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21284 18170 21312 18686
rect 21192 18142 21312 18170
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20916 17746 20944 18022
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20824 16646 20944 16674
rect 20812 16040 20864 16046
rect 20810 16008 20812 16017
rect 20864 16008 20866 16017
rect 20810 15943 20866 15952
rect 20810 15736 20866 15745
rect 20720 15700 20772 15706
rect 20810 15671 20866 15680
rect 20720 15642 20772 15648
rect 20824 15638 20852 15671
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20628 15428 20680 15434
rect 20628 15370 20680 15376
rect 20732 15094 20760 15506
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19870 12540 20178 12549
rect 19870 12538 19876 12540
rect 19932 12538 19956 12540
rect 20012 12538 20036 12540
rect 20092 12538 20116 12540
rect 20172 12538 20178 12540
rect 19932 12486 19934 12538
rect 20114 12486 20116 12538
rect 19870 12484 19876 12486
rect 19932 12484 19956 12486
rect 20012 12484 20036 12486
rect 20092 12484 20116 12486
rect 20172 12484 20178 12486
rect 19870 12475 20178 12484
rect 20548 12434 20576 12718
rect 20640 12714 20668 14826
rect 20824 14482 20852 15302
rect 20916 15065 20944 16646
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 15570 21036 16390
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21100 15706 21128 15914
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21086 15464 21142 15473
rect 21086 15399 21142 15408
rect 20902 15056 20958 15065
rect 20902 14991 20958 15000
rect 20996 14816 21048 14822
rect 21100 14804 21128 15399
rect 21192 14929 21220 18142
rect 21270 17640 21326 17649
rect 21270 17575 21272 17584
rect 21324 17575 21326 17584
rect 21272 17546 21324 17552
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21284 15638 21312 16594
rect 21376 16114 21404 18158
rect 21468 17610 21496 18799
rect 21560 18630 21588 18838
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 22204 18426 22232 19858
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22296 19689 22324 19722
rect 22282 19680 22338 19689
rect 22282 19615 22338 19624
rect 22388 19394 22416 20334
rect 22480 20262 22508 20402
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22296 19378 22416 19394
rect 22296 19372 22428 19378
rect 22296 19366 22376 19372
rect 22296 18970 22324 19366
rect 22376 19314 22428 19320
rect 22664 19310 22692 20742
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22756 20074 22784 20402
rect 22940 20398 22968 20839
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 22756 20046 22876 20074
rect 22848 19990 22876 20046
rect 22836 19984 22888 19990
rect 22836 19926 22888 19932
rect 22744 19848 22796 19854
rect 22742 19816 22744 19825
rect 22836 19848 22888 19854
rect 22796 19816 22798 19825
rect 22836 19790 22888 19796
rect 22742 19751 22798 19760
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 22756 19310 22784 19654
rect 22848 19514 22876 19790
rect 22940 19689 22968 20198
rect 23110 20088 23166 20097
rect 23110 20023 23166 20032
rect 23124 19922 23152 20023
rect 23492 19922 23520 20198
rect 23768 19922 23796 20334
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24136 19922 24164 20198
rect 24228 19990 24256 20742
rect 25148 20398 25176 21286
rect 26252 21078 26280 21286
rect 26240 21072 26292 21078
rect 26240 21014 26292 21020
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25792 20398 25820 20878
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 24216 19984 24268 19990
rect 24216 19926 24268 19932
rect 25792 19922 25820 20334
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 23020 19712 23072 19718
rect 22926 19680 22982 19689
rect 23020 19654 23072 19660
rect 22926 19615 22982 19624
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 22388 18970 22416 19178
rect 22940 19156 22968 19615
rect 23032 19310 23060 19654
rect 23216 19514 23244 19858
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 23020 19168 23072 19174
rect 22940 19136 23020 19156
rect 24584 19168 24636 19174
rect 23072 19136 23074 19145
rect 22940 19128 23018 19136
rect 24584 19110 24636 19116
rect 24676 19168 24728 19174
rect 25044 19168 25096 19174
rect 24676 19110 24728 19116
rect 24964 19116 25044 19122
rect 24964 19110 25096 19116
rect 23018 19071 23074 19080
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 24596 18834 24624 19110
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 24584 18828 24636 18834
rect 24584 18770 24636 18776
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 22848 18426 22876 18566
rect 22940 18465 22968 18770
rect 22926 18456 22982 18465
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22836 18420 22888 18426
rect 24044 18426 24072 18770
rect 22926 18391 22982 18400
rect 24032 18420 24084 18426
rect 22836 18362 22888 18368
rect 24032 18362 24084 18368
rect 23296 18352 23348 18358
rect 22466 18320 22522 18329
rect 23296 18294 23348 18300
rect 22466 18255 22522 18264
rect 21914 18184 21970 18193
rect 21914 18119 21970 18128
rect 21928 17746 21956 18119
rect 22480 18057 22508 18255
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 22466 18048 22522 18057
rect 22466 17983 22522 17992
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21560 17270 21588 17614
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21272 15632 21324 15638
rect 21272 15574 21324 15580
rect 21284 15162 21312 15574
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21178 14920 21234 14929
rect 21178 14855 21234 14864
rect 21100 14776 21220 14804
rect 20996 14758 21048 14764
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 14362 20852 14418
rect 20824 14334 20944 14362
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13258 20760 13874
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20916 12850 20944 14334
rect 21008 14074 21036 14758
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21008 13326 21036 13806
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 19628 12406 19932 12434
rect 19064 12378 19116 12384
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18708 12102 18736 12242
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18524 11694 18552 12038
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18236 11144 18288 11150
rect 18156 11104 18236 11132
rect 17684 11086 17736 11092
rect 18236 11086 18288 11092
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18248 10606 18276 10746
rect 18236 10600 18288 10606
rect 18156 10560 18236 10588
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 10130 18000 10406
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17500 9444 17552 9450
rect 17420 9404 17500 9432
rect 17500 9386 17552 9392
rect 17960 9376 18012 9382
rect 18064 9364 18092 10066
rect 18012 9336 18092 9364
rect 17960 9318 18012 9324
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17052 7410 17080 7822
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17040 7404 17092 7410
rect 16868 7364 17040 7392
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 6798 16804 7142
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15948 4146 15976 4422
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 16580 4072 16632 4078
rect 16500 4032 16580 4060
rect 16500 3602 16528 4032
rect 16580 4014 16632 4020
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15028 2417 15056 2790
rect 15212 2650 15240 3334
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15014 2408 15070 2417
rect 15212 2378 15240 2586
rect 16040 2514 16068 2926
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15014 2343 15070 2352
rect 15200 2372 15252 2378
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 14832 1828 14884 1834
rect 14832 1770 14884 1776
rect 13084 1760 13136 1766
rect 13084 1702 13136 1708
rect 13268 1760 13320 1766
rect 13268 1702 13320 1708
rect 13820 1760 13872 1766
rect 13820 1702 13872 1708
rect 13096 1494 13124 1702
rect 13084 1488 13136 1494
rect 13084 1430 13136 1436
rect 13280 1426 13308 1702
rect 13268 1420 13320 1426
rect 13268 1362 13320 1368
rect 12992 1216 13044 1222
rect 12992 1158 13044 1164
rect 13832 882 13860 1702
rect 14936 1494 14964 2042
rect 15028 1834 15056 2343
rect 15200 2314 15252 2320
rect 15396 2038 15424 2450
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 2106 15792 2246
rect 15948 2106 15976 2382
rect 15752 2100 15804 2106
rect 15752 2042 15804 2048
rect 15936 2100 15988 2106
rect 15936 2042 15988 2048
rect 15384 2032 15436 2038
rect 15384 1974 15436 1980
rect 16132 1902 16160 3062
rect 16224 2514 16252 3334
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16408 2854 16436 2926
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16028 1896 16080 1902
rect 16028 1838 16080 1844
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 15016 1828 15068 1834
rect 15016 1770 15068 1776
rect 16040 1562 16068 1838
rect 16500 1834 16528 3538
rect 16776 2990 16804 6734
rect 16868 3466 16896 7364
rect 17040 7346 17092 7352
rect 17420 7342 17448 7754
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17144 5370 17172 6394
rect 17972 5846 18000 9318
rect 18156 8838 18184 10560
rect 18236 10542 18288 10548
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18340 10198 18368 10474
rect 18432 10266 18460 11494
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 18432 9738 18460 10202
rect 18432 9710 18552 9738
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18248 8634 18276 8978
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18432 8430 18460 9522
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18524 7886 18552 9710
rect 18616 9500 18644 11698
rect 18708 10742 18736 12038
rect 19210 11996 19518 12005
rect 19210 11994 19216 11996
rect 19272 11994 19296 11996
rect 19352 11994 19376 11996
rect 19432 11994 19456 11996
rect 19512 11994 19518 11996
rect 19272 11942 19274 11994
rect 19454 11942 19456 11994
rect 19210 11940 19216 11942
rect 19272 11940 19296 11942
rect 19352 11940 19376 11942
rect 19432 11940 19456 11942
rect 19512 11940 19518 11942
rect 19210 11931 19518 11940
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11558 19288 11698
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19628 11354 19656 12310
rect 19800 11688 19852 11694
rect 19720 11636 19800 11642
rect 19720 11630 19852 11636
rect 19720 11614 19840 11630
rect 19720 11558 19748 11614
rect 19904 11558 19932 12406
rect 20456 12406 20576 12434
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 19996 11694 20024 12310
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20180 11694 20208 12242
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19812 11354 19840 11494
rect 19870 11452 20178 11461
rect 19870 11450 19876 11452
rect 19932 11450 19956 11452
rect 20012 11450 20036 11452
rect 20092 11450 20116 11452
rect 20172 11450 20178 11452
rect 19932 11398 19934 11450
rect 20114 11398 20116 11450
rect 19870 11396 19876 11398
rect 19932 11396 19956 11398
rect 20012 11396 20036 11398
rect 20092 11396 20116 11398
rect 20172 11396 20178 11398
rect 19870 11387 20178 11396
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 20364 11286 20392 12038
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18800 10606 18828 11018
rect 19210 10908 19518 10917
rect 19210 10906 19216 10908
rect 19272 10906 19296 10908
rect 19352 10906 19376 10908
rect 19432 10906 19456 10908
rect 19512 10906 19518 10908
rect 19272 10854 19274 10906
rect 19454 10854 19456 10906
rect 19210 10852 19216 10854
rect 19272 10852 19296 10854
rect 19352 10852 19376 10854
rect 19432 10852 19456 10854
rect 19512 10852 19518 10854
rect 19210 10843 19518 10852
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18708 10266 18736 10542
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 9518 18920 10066
rect 18696 9512 18748 9518
rect 18616 9472 18696 9500
rect 18696 9454 18748 9460
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18708 8276 18736 9454
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18800 9110 18828 9318
rect 18892 9178 18920 9454
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18984 8922 19012 10406
rect 18892 8894 19012 8922
rect 18892 8430 18920 8894
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18788 8288 18840 8294
rect 18708 8248 18788 8276
rect 18788 8230 18840 8236
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18248 6458 18276 6802
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18340 5778 18368 6190
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17144 4282 17172 5102
rect 17604 4622 17632 5102
rect 18064 4622 18092 5306
rect 18340 5166 18368 5510
rect 18432 5234 18460 6258
rect 18524 6186 18552 7822
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18524 5370 18552 5510
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18524 4826 18552 5034
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18616 4758 18644 8026
rect 18708 6254 18736 8026
rect 18800 7342 18828 8230
rect 18892 8090 18920 8366
rect 18984 8362 19012 8774
rect 19076 8412 19104 10474
rect 19210 9820 19518 9829
rect 19210 9818 19216 9820
rect 19272 9818 19296 9820
rect 19352 9818 19376 9820
rect 19432 9818 19456 9820
rect 19512 9818 19518 9820
rect 19272 9766 19274 9818
rect 19454 9766 19456 9818
rect 19210 9764 19216 9766
rect 19272 9764 19296 9766
rect 19352 9764 19376 9766
rect 19432 9764 19456 9766
rect 19512 9764 19518 9766
rect 19210 9755 19518 9764
rect 19210 8732 19518 8741
rect 19210 8730 19216 8732
rect 19272 8730 19296 8732
rect 19352 8730 19376 8732
rect 19432 8730 19456 8732
rect 19512 8730 19518 8732
rect 19272 8678 19274 8730
rect 19454 8678 19456 8730
rect 19210 8676 19216 8678
rect 19272 8676 19296 8678
rect 19352 8676 19376 8678
rect 19432 8676 19456 8678
rect 19512 8676 19518 8678
rect 19210 8667 19518 8676
rect 19156 8424 19208 8430
rect 19076 8384 19156 8412
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 19076 7970 19104 8384
rect 19156 8366 19208 8372
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19628 8090 19656 8366
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 18892 7954 19104 7970
rect 18880 7948 19104 7954
rect 18932 7942 19104 7948
rect 18880 7890 18932 7896
rect 18892 7698 18920 7890
rect 18892 7670 19012 7698
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18892 7342 18920 7482
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18800 6798 18828 7278
rect 18984 7002 19012 7670
rect 19210 7644 19518 7653
rect 19210 7642 19216 7644
rect 19272 7642 19296 7644
rect 19352 7642 19376 7644
rect 19432 7642 19456 7644
rect 19512 7642 19518 7644
rect 19272 7590 19274 7642
rect 19454 7590 19456 7642
rect 19210 7588 19216 7590
rect 19272 7588 19296 7590
rect 19352 7588 19376 7590
rect 19432 7588 19456 7590
rect 19512 7588 19518 7590
rect 19210 7579 19518 7588
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 18788 6792 18840 6798
rect 18984 6746 19012 6938
rect 18788 6734 18840 6740
rect 18800 6458 18828 6734
rect 18892 6718 19012 6746
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18708 5574 18736 5782
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18696 5296 18748 5302
rect 18800 5284 18828 6394
rect 18892 6118 18920 6718
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 6254 19012 6598
rect 19210 6556 19518 6565
rect 19210 6554 19216 6556
rect 19272 6554 19296 6556
rect 19352 6554 19376 6556
rect 19432 6554 19456 6556
rect 19512 6554 19518 6556
rect 19272 6502 19274 6554
rect 19454 6502 19456 6554
rect 19210 6500 19216 6502
rect 19272 6500 19296 6502
rect 19352 6500 19376 6502
rect 19432 6500 19456 6502
rect 19512 6500 19518 6502
rect 19210 6491 19518 6500
rect 19720 6322 19748 11018
rect 20272 10470 20300 11086
rect 20456 10810 20484 12406
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20640 11762 20668 12242
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20732 11626 20760 12582
rect 21008 12442 21036 13126
rect 21100 12782 21128 13738
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21192 12628 21220 14776
rect 21284 14550 21312 15098
rect 21376 14618 21404 16050
rect 21456 15904 21508 15910
rect 21652 15881 21680 17138
rect 21824 17128 21876 17134
rect 21744 17088 21824 17116
rect 21744 16998 21772 17088
rect 21824 17070 21876 17076
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21456 15846 21508 15852
rect 21638 15872 21694 15881
rect 21468 15570 21496 15846
rect 21638 15807 21694 15816
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21652 15434 21680 15807
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21468 14890 21496 15302
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21468 13190 21496 14826
rect 21560 14414 21588 14894
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 13326 21588 14350
rect 21652 14074 21680 14418
rect 21744 14249 21772 16934
rect 22098 16144 22154 16153
rect 22098 16079 22154 16088
rect 22112 16046 22140 16079
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21928 15722 21956 15914
rect 22100 15904 22152 15910
rect 22204 15892 22232 17682
rect 22480 17610 22508 17983
rect 23032 17678 23060 18158
rect 23308 18154 23336 18294
rect 23296 18148 23348 18154
rect 23296 18090 23348 18096
rect 23308 17746 23336 18090
rect 23296 17740 23348 17746
rect 23296 17682 23348 17688
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 22376 17536 22428 17542
rect 22376 17478 22428 17484
rect 22388 16046 22416 17478
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22664 16998 22692 17138
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22466 16824 22522 16833
rect 22466 16759 22522 16768
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22152 15864 22232 15892
rect 22100 15846 22152 15852
rect 22296 15722 22324 15982
rect 21928 15694 22324 15722
rect 21822 15600 21878 15609
rect 21822 15535 21824 15544
rect 21876 15535 21878 15544
rect 22100 15564 22152 15570
rect 21824 15506 21876 15512
rect 22100 15506 22152 15512
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 21928 14482 21956 15030
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 22020 14414 22048 14894
rect 22008 14408 22060 14414
rect 21928 14356 22008 14362
rect 21928 14350 22060 14356
rect 21928 14334 22048 14350
rect 22112 14346 22140 15506
rect 22388 14618 22416 15982
rect 22480 15706 22508 16759
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22572 15094 22600 16934
rect 22940 16250 22968 17070
rect 23032 16794 23060 17614
rect 23124 17270 23152 17614
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22742 16144 22798 16153
rect 22742 16079 22798 16088
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22560 15088 22612 15094
rect 22560 15030 22612 15036
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22100 14340 22152 14346
rect 21730 14240 21786 14249
rect 21730 14175 21786 14184
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 21652 13394 21680 14010
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21744 13530 21772 13738
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21928 13394 21956 14334
rect 22100 14282 22152 14288
rect 22468 14272 22520 14278
rect 22098 14240 22154 14249
rect 22468 14214 22520 14220
rect 22098 14175 22154 14184
rect 22112 13462 22140 14175
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22204 13530 22232 13738
rect 22296 13530 22324 13806
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21100 12600 21220 12628
rect 21364 12640 21416 12646
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 19870 10364 20178 10373
rect 19870 10362 19876 10364
rect 19932 10362 19956 10364
rect 20012 10362 20036 10364
rect 20092 10362 20116 10364
rect 20172 10362 20178 10364
rect 19932 10310 19934 10362
rect 20114 10310 20116 10362
rect 19870 10308 19876 10310
rect 19932 10308 19956 10310
rect 20012 10308 20036 10310
rect 20092 10308 20116 10310
rect 20172 10308 20178 10310
rect 19870 10299 20178 10308
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20088 9382 20116 9454
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19870 9276 20178 9285
rect 19870 9274 19876 9276
rect 19932 9274 19956 9276
rect 20012 9274 20036 9276
rect 20092 9274 20116 9276
rect 20172 9274 20178 9276
rect 19932 9222 19934 9274
rect 20114 9222 20116 9274
rect 19870 9220 19876 9222
rect 19932 9220 19956 9222
rect 20012 9220 20036 9222
rect 20092 9220 20116 9222
rect 20172 9220 20178 9222
rect 19870 9211 20178 9220
rect 20272 8838 20300 10406
rect 20456 10198 20484 10542
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20364 9110 20392 9454
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20456 9042 20484 10134
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20456 8430 20484 8978
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19812 8022 19840 8230
rect 19870 8188 20178 8197
rect 19870 8186 19876 8188
rect 19932 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20178 8188
rect 19932 8134 19934 8186
rect 20114 8134 20116 8186
rect 19870 8132 19876 8134
rect 19932 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20178 8134
rect 19870 8123 20178 8132
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 20456 7410 20484 8366
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 19870 7100 20178 7109
rect 19870 7098 19876 7100
rect 19932 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20178 7100
rect 19932 7046 19934 7098
rect 20114 7046 20116 7098
rect 19870 7044 19876 7046
rect 19932 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20178 7046
rect 19870 7035 20178 7044
rect 20456 6866 20484 7346
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20548 6746 20576 11290
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20640 9178 20668 9454
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20732 8106 20760 10746
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20732 8078 20852 8106
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20732 7342 20760 7890
rect 20628 7336 20680 7342
rect 20626 7304 20628 7313
rect 20720 7336 20772 7342
rect 20680 7304 20682 7313
rect 20720 7278 20772 7284
rect 20626 7239 20682 7248
rect 20456 6730 20576 6746
rect 20444 6724 20576 6730
rect 20496 6718 20576 6724
rect 20444 6666 20496 6672
rect 20456 6390 20484 6666
rect 20444 6384 20496 6390
rect 20444 6326 20496 6332
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19616 6180 19668 6186
rect 19616 6122 19668 6128
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5778 18920 6054
rect 19076 5846 19104 6122
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19628 5778 19656 6122
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 19210 5468 19518 5477
rect 19210 5466 19216 5468
rect 19272 5466 19296 5468
rect 19352 5466 19376 5468
rect 19432 5466 19456 5468
rect 19512 5466 19518 5468
rect 19272 5414 19274 5466
rect 19454 5414 19456 5466
rect 19210 5412 19216 5414
rect 19272 5412 19296 5414
rect 19352 5412 19376 5414
rect 19432 5412 19456 5414
rect 19512 5412 19518 5414
rect 19210 5403 19518 5412
rect 18748 5256 18828 5284
rect 18696 5238 18748 5244
rect 19628 5030 19656 5714
rect 19720 5642 19748 6258
rect 20640 6254 20668 7239
rect 20824 6882 20852 8078
rect 20916 7954 20944 8230
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 21008 7750 21036 12378
rect 21100 9450 21128 12600
rect 21364 12582 21416 12588
rect 21376 12374 21404 12582
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21468 11762 21496 12106
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21192 11286 21220 11630
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21284 11218 21312 11494
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21284 10266 21312 10474
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21376 10062 21404 11630
rect 21468 10538 21496 11698
rect 21560 11694 21588 13262
rect 21652 12986 21680 13330
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21732 13252 21784 13258
rect 21732 13194 21784 13200
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21744 12782 21772 13194
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 22020 12646 22048 13262
rect 22480 13190 22508 14214
rect 22572 13977 22600 15030
rect 22664 14822 22692 15982
rect 22756 15706 22784 16079
rect 22926 16008 22982 16017
rect 23032 15994 23060 16526
rect 23124 16182 23152 17206
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23216 16998 23244 17138
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23216 16658 23244 16730
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23112 16176 23164 16182
rect 23112 16118 23164 16124
rect 23216 16046 23244 16390
rect 22982 15966 23060 15994
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 22926 15943 22982 15952
rect 22940 15910 22968 15943
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 14521 22692 14758
rect 22650 14512 22706 14521
rect 22650 14447 22706 14456
rect 22558 13968 22614 13977
rect 22558 13903 22614 13912
rect 22756 13870 22784 15370
rect 22940 15094 22968 15846
rect 23124 15706 23152 15846
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23308 15502 23336 17682
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23400 16658 23428 17478
rect 23492 17134 23520 17682
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23492 16046 23520 16934
rect 23584 16658 23612 17478
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23676 16522 23704 17478
rect 24136 17338 24164 18770
rect 24688 18737 24716 19110
rect 24964 19094 25084 19110
rect 24674 18728 24730 18737
rect 24674 18663 24730 18672
rect 24492 18216 24544 18222
rect 24544 18164 24716 18170
rect 24492 18158 24716 18164
rect 24504 18142 24716 18158
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24596 17746 24624 18022
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23952 16794 23980 16934
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23664 16516 23716 16522
rect 23664 16458 23716 16464
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23676 15706 23704 16050
rect 24136 16046 24164 17274
rect 24228 16658 24256 17682
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24412 17202 24440 17274
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24412 16697 24440 17138
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 24398 16688 24454 16697
rect 24216 16652 24268 16658
rect 24398 16623 24454 16632
rect 24492 16652 24544 16658
rect 24216 16594 24268 16600
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 23664 15700 23716 15706
rect 23664 15642 23716 15648
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22848 14074 22876 14418
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22848 13870 22876 14010
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22940 13734 22968 14894
rect 23400 14822 23428 15506
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23216 13938 23244 14350
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 13938 23336 14214
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23400 13734 23428 14758
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23584 13870 23612 14554
rect 23676 14482 23704 15030
rect 23860 14482 23888 15982
rect 24136 15094 24164 15982
rect 24412 15502 24440 16623
rect 24492 16594 24544 16600
rect 24504 16250 24532 16594
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24596 15910 24624 17002
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24596 15745 24624 15846
rect 24582 15736 24638 15745
rect 24688 15706 24716 18142
rect 24964 18086 24992 19094
rect 25148 18970 25176 19654
rect 25608 19310 25636 19790
rect 25792 19378 25820 19858
rect 25884 19786 25912 20198
rect 26436 20058 26464 20742
rect 26528 20330 26556 21286
rect 26896 20330 26924 21558
rect 28276 21486 28304 21927
rect 28998 21856 29054 21865
rect 28998 21791 29054 21800
rect 29012 21554 29040 21791
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 29184 21480 29236 21486
rect 29184 21422 29236 21428
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 27644 21244 27952 21253
rect 27644 21242 27650 21244
rect 27706 21242 27730 21244
rect 27786 21242 27810 21244
rect 27866 21242 27890 21244
rect 27946 21242 27952 21244
rect 27706 21190 27708 21242
rect 27888 21190 27890 21242
rect 27644 21188 27650 21190
rect 27706 21188 27730 21190
rect 27786 21188 27810 21190
rect 27866 21188 27890 21190
rect 27946 21188 27952 21190
rect 27644 21179 27952 21188
rect 28000 21026 28028 21286
rect 28184 21078 28212 21286
rect 27816 20998 28028 21026
rect 28172 21072 28224 21078
rect 28172 21014 28224 21020
rect 27816 20942 27844 20998
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 26984 20700 27292 20709
rect 26984 20698 26990 20700
rect 27046 20698 27070 20700
rect 27126 20698 27150 20700
rect 27206 20698 27230 20700
rect 27286 20698 27292 20700
rect 27046 20646 27048 20698
rect 27228 20646 27230 20698
rect 26984 20644 26990 20646
rect 27046 20644 27070 20646
rect 27126 20644 27150 20646
rect 27206 20644 27230 20646
rect 27286 20644 27292 20646
rect 26984 20635 27292 20644
rect 27816 20398 27844 20878
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 26516 20324 26568 20330
rect 26516 20266 26568 20272
rect 26884 20324 26936 20330
rect 26884 20266 26936 20272
rect 27644 20156 27952 20165
rect 27644 20154 27650 20156
rect 27706 20154 27730 20156
rect 27786 20154 27810 20156
rect 27866 20154 27890 20156
rect 27946 20154 27952 20156
rect 27706 20102 27708 20154
rect 27888 20102 27890 20154
rect 27644 20100 27650 20102
rect 27706 20100 27730 20102
rect 27786 20100 27810 20102
rect 27866 20100 27890 20102
rect 27946 20100 27952 20102
rect 27644 20091 27952 20100
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 27528 19984 27580 19990
rect 26514 19952 26570 19961
rect 26514 19887 26570 19896
rect 27526 19952 27528 19961
rect 27580 19952 27582 19961
rect 27526 19887 27582 19896
rect 27988 19916 28040 19922
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24964 17746 24992 18022
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24780 17542 24808 17682
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24872 17134 24900 17546
rect 25056 17490 25084 18158
rect 24964 17462 25084 17490
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24872 16726 24900 17070
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24780 15706 24808 15982
rect 24582 15671 24638 15680
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24688 15586 24716 15642
rect 24492 15564 24544 15570
rect 24688 15558 24808 15586
rect 24872 15570 24900 16662
rect 24964 16454 24992 17462
rect 25148 17338 25176 18158
rect 25240 17882 25268 18226
rect 25332 18193 25360 19246
rect 25516 19174 25544 19246
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 25608 18970 25636 19246
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25504 18624 25556 18630
rect 25424 18572 25504 18578
rect 25424 18566 25556 18572
rect 25424 18550 25544 18566
rect 25318 18184 25374 18193
rect 25318 18119 25374 18128
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25228 16992 25280 16998
rect 25332 16980 25360 18022
rect 25424 17202 25452 18550
rect 25608 17202 25636 18906
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25280 16952 25360 16980
rect 25228 16934 25280 16940
rect 25044 16720 25096 16726
rect 25044 16662 25096 16668
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24964 15978 24992 16390
rect 25056 16046 25084 16662
rect 25240 16590 25268 16934
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25044 16040 25096 16046
rect 25044 15982 25096 15988
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24492 15506 24544 15512
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24124 15088 24176 15094
rect 24124 15030 24176 15036
rect 24504 15026 24532 15506
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23768 13530 23796 14418
rect 24136 14414 24164 14894
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23952 13394 23980 14214
rect 24228 13394 24256 14758
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24320 14278 24348 14418
rect 24412 14385 24440 14894
rect 24504 14618 24532 14962
rect 24596 14958 24624 15302
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24398 14376 24454 14385
rect 24398 14311 24454 14320
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24412 13530 24440 14311
rect 24596 14074 24624 14418
rect 24688 14414 24716 15438
rect 24780 14482 24808 15558
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24964 14958 24992 15914
rect 25424 15366 25452 17138
rect 25608 17066 25636 17138
rect 25504 17060 25556 17066
rect 25504 17002 25556 17008
rect 25596 17060 25648 17066
rect 25596 17002 25648 17008
rect 25516 16794 25544 17002
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25700 16454 25728 16594
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25792 15570 25820 19314
rect 25884 18057 25912 19314
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 26068 18222 26096 18906
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 26148 18148 26200 18154
rect 26148 18090 26200 18096
rect 25870 18048 25926 18057
rect 25870 17983 25926 17992
rect 25872 17060 25924 17066
rect 25872 17002 25924 17008
rect 25884 16658 25912 17002
rect 26056 16992 26108 16998
rect 26056 16934 26108 16940
rect 26068 16658 26096 16934
rect 26160 16833 26188 18090
rect 26332 17808 26384 17814
rect 26332 17750 26384 17756
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 26252 17134 26280 17478
rect 26344 17134 26372 17750
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26146 16824 26202 16833
rect 26146 16759 26202 16768
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 25976 16538 26004 16594
rect 25884 16510 26004 16538
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25884 15450 25912 16510
rect 26160 16250 26188 16594
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 25608 15422 25912 15450
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 25228 14952 25280 14958
rect 25608 14906 25636 15422
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25280 14900 25636 14906
rect 25228 14894 25636 14900
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24596 13462 24624 14010
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24872 13530 24900 13806
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24584 13456 24636 13462
rect 24584 13398 24636 13404
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 24412 12850 24440 13262
rect 24964 13258 24992 14894
rect 25056 14618 25084 14894
rect 25240 14890 25636 14894
rect 25136 14884 25188 14890
rect 25136 14826 25188 14832
rect 25240 14884 25648 14890
rect 25240 14878 25596 14884
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 25148 13530 25176 14826
rect 25240 14482 25268 14878
rect 25596 14826 25648 14832
rect 25504 14816 25556 14822
rect 25504 14758 25556 14764
rect 25516 14550 25544 14758
rect 25504 14544 25556 14550
rect 25504 14486 25556 14492
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25240 14074 25268 14282
rect 25700 14278 25728 15302
rect 25964 15156 26016 15162
rect 25964 15098 26016 15104
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25884 14482 25912 14758
rect 25976 14482 26004 15098
rect 25872 14476 25924 14482
rect 25872 14418 25924 14424
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25240 13462 25268 14010
rect 25608 13870 25636 14214
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25332 13530 25360 13806
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25228 13456 25280 13462
rect 25228 13398 25280 13404
rect 25700 13326 25728 14214
rect 26068 13394 26096 16050
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26160 14346 26188 14418
rect 26252 14385 26280 17070
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26238 14376 26294 14385
rect 26148 14340 26200 14346
rect 26344 14346 26372 14554
rect 26238 14311 26294 14320
rect 26332 14340 26384 14346
rect 26148 14282 26200 14288
rect 26332 14282 26384 14288
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26344 13394 26372 13806
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21652 10282 21680 12582
rect 21824 12368 21876 12374
rect 21824 12310 21876 12316
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21744 11830 21772 12038
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 21744 11354 21772 11630
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21560 10254 21680 10282
rect 21560 10130 21588 10254
rect 21744 10130 21772 10950
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21284 9178 21312 9318
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 20824 6866 21036 6882
rect 20720 6860 20772 6866
rect 20824 6860 21048 6866
rect 20824 6854 20996 6860
rect 20720 6802 20772 6808
rect 20996 6802 21048 6808
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 19870 6012 20178 6021
rect 19870 6010 19876 6012
rect 19932 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20178 6012
rect 19932 5958 19934 6010
rect 20114 5958 20116 6010
rect 19870 5956 19876 5958
rect 19932 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20178 5958
rect 19870 5947 20178 5956
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 19628 4690 19656 4966
rect 19870 4924 20178 4933
rect 19870 4922 19876 4924
rect 19932 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20178 4924
rect 19932 4870 19934 4922
rect 20114 4870 20116 4922
rect 19870 4868 19876 4870
rect 19932 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20178 4870
rect 19870 4859 20178 4868
rect 20732 4842 20760 6802
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21008 6390 21036 6598
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 20640 4814 20760 4842
rect 20640 4758 20668 4814
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16580 2304 16632 2310
rect 16632 2252 16712 2258
rect 16580 2246 16712 2252
rect 16592 2230 16712 2246
rect 16684 2106 16712 2230
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 16488 1828 16540 1834
rect 16488 1770 16540 1776
rect 16028 1556 16080 1562
rect 16028 1498 16080 1504
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 16500 1426 16528 1770
rect 16776 1562 16804 2926
rect 16868 2310 16896 3402
rect 17328 2990 17356 4082
rect 17788 3194 17816 4218
rect 17868 3936 17920 3942
rect 17972 3890 18000 4422
rect 17920 3884 18000 3890
rect 17868 3878 18000 3884
rect 17880 3862 18000 3878
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 16960 2650 16988 2790
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 17052 2106 17080 2790
rect 17512 2582 17540 2790
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 17512 2038 17540 2518
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17788 1902 17816 3130
rect 18248 2514 18276 4626
rect 19210 4380 19518 4389
rect 19210 4378 19216 4380
rect 19272 4378 19296 4380
rect 19352 4378 19376 4380
rect 19432 4378 19456 4380
rect 19512 4378 19518 4380
rect 19272 4326 19274 4378
rect 19454 4326 19456 4378
rect 19210 4324 19216 4326
rect 19272 4324 19296 4326
rect 19352 4324 19376 4326
rect 19432 4324 19456 4326
rect 19512 4324 19518 4326
rect 19210 4315 19518 4324
rect 19628 4282 19656 4626
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20088 4282 20116 4558
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 18340 4078 18368 4218
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 19210 3292 19518 3301
rect 19210 3290 19216 3292
rect 19272 3290 19296 3292
rect 19352 3290 19376 3292
rect 19432 3290 19456 3292
rect 19512 3290 19518 3292
rect 19272 3238 19274 3290
rect 19454 3238 19456 3290
rect 19210 3236 19216 3238
rect 19272 3236 19296 3238
rect 19352 3236 19376 3238
rect 19432 3236 19456 3238
rect 19512 3236 19518 3238
rect 19210 3227 19518 3236
rect 19628 2922 19656 4218
rect 20088 4078 20116 4218
rect 20732 4214 20760 4626
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19870 3836 20178 3845
rect 19870 3834 19876 3836
rect 19932 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20178 3836
rect 19932 3782 19934 3834
rect 20114 3782 20116 3834
rect 19870 3780 19876 3782
rect 19932 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20178 3782
rect 19870 3771 20178 3780
rect 21008 3670 21036 6326
rect 21100 6254 21128 9046
rect 21560 8498 21588 10066
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 21468 6186 21496 7346
rect 21836 6866 21864 12310
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 10130 21956 12038
rect 22020 11218 22048 12582
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22112 10810 22140 11086
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22848 10606 22876 12242
rect 23032 11830 23060 12242
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 23124 10606 23152 12718
rect 23768 12646 23796 12786
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23768 12306 23796 12582
rect 23756 12300 23808 12306
rect 23756 12242 23808 12248
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23492 11830 23520 12038
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23308 11218 23336 11494
rect 23492 11354 23520 11562
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23584 11218 23612 12038
rect 23860 11762 23888 12038
rect 26436 11830 26464 12106
rect 26424 11824 26476 11830
rect 26424 11766 26476 11772
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25596 11688 25648 11694
rect 25596 11630 25648 11636
rect 25780 11688 25832 11694
rect 25780 11630 25832 11636
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 24216 11620 24268 11626
rect 24216 11562 24268 11568
rect 24228 11286 24256 11562
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25240 11354 25268 11494
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23768 10810 23796 11154
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 22836 10600 22888 10606
rect 23112 10600 23164 10606
rect 22888 10548 23060 10554
rect 22836 10542 23060 10548
rect 23112 10542 23164 10548
rect 22008 10532 22060 10538
rect 22848 10526 23060 10542
rect 24228 10538 24256 11222
rect 25332 11082 25360 11630
rect 25608 11286 25636 11630
rect 25792 11354 25820 11630
rect 25780 11348 25832 11354
rect 25780 11290 25832 11296
rect 25596 11280 25648 11286
rect 25596 11222 25648 11228
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24872 10606 24900 10950
rect 25884 10810 25912 11630
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 22008 10474 22060 10480
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21928 9722 21956 10066
rect 22020 10062 22048 10474
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21928 9110 21956 9658
rect 22020 9518 22048 9998
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9586 22140 9862
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 22020 8906 22048 9454
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 22112 8378 22140 8978
rect 22296 8974 22324 9318
rect 22388 9178 22416 10134
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22468 9444 22520 9450
rect 22468 9386 22520 9392
rect 22480 9178 22508 9386
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22940 9042 22968 9862
rect 23032 9674 23060 10526
rect 24216 10532 24268 10538
rect 24216 10474 24268 10480
rect 24228 10198 24256 10474
rect 24872 10198 24900 10542
rect 25884 10266 25912 10610
rect 26160 10606 26188 10950
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 26344 10266 26372 10542
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 23032 9646 23152 9674
rect 23492 9654 23520 10066
rect 23124 9586 23152 9646
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22848 8906 22876 8978
rect 22836 8900 22888 8906
rect 22836 8842 22888 8848
rect 22848 8498 22876 8842
rect 23124 8634 23152 9522
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 23124 8430 23152 8570
rect 23216 8430 23244 8570
rect 22020 8350 22140 8378
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 21824 6860 21876 6866
rect 21744 6820 21824 6848
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21456 6180 21508 6186
rect 21456 6122 21508 6128
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21192 4758 21220 4966
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21284 4690 21312 5510
rect 21468 5370 21496 6122
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21468 5114 21496 5306
rect 21560 5234 21588 6598
rect 21744 6254 21772 6820
rect 21824 6802 21876 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21836 6458 21864 6666
rect 21928 6458 21956 6802
rect 22020 6746 22048 8350
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 22112 7954 22140 8230
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22664 7562 22692 8366
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22204 7534 22692 7562
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22112 7002 22140 7210
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22020 6718 22140 6746
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21640 5160 21692 5166
rect 21468 5108 21640 5114
rect 21468 5102 21692 5108
rect 21468 5086 21680 5102
rect 21744 5098 21772 6190
rect 21836 5710 21864 6394
rect 22020 6254 22048 6598
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22112 6100 22140 6718
rect 21928 6072 22140 6100
rect 21928 5778 21956 6072
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21836 5302 21864 5646
rect 21824 5296 21876 5302
rect 21824 5238 21876 5244
rect 21928 5234 21956 5714
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22020 5302 22048 5510
rect 22008 5296 22060 5302
rect 22008 5238 22060 5244
rect 22100 5296 22152 5302
rect 22204 5284 22232 7534
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22296 6866 22324 7142
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22284 6180 22336 6186
rect 22284 6122 22336 6128
rect 22152 5256 22232 5284
rect 22100 5238 22152 5244
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 22020 5166 22048 5238
rect 22008 5160 22060 5166
rect 22296 5148 22324 6122
rect 22388 5914 22416 7346
rect 22756 7342 22784 8298
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 7954 23060 8230
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23400 7410 23428 8366
rect 24044 8362 24072 8774
rect 24228 8362 24256 10134
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 25872 10124 25924 10130
rect 25872 10066 25924 10072
rect 25056 9518 25084 10066
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 9722 25176 9862
rect 25792 9722 25820 10066
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 24492 9444 24544 9450
rect 24492 9386 24544 9392
rect 24504 9330 24532 9386
rect 24504 9302 24624 9330
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24504 8634 24532 8978
rect 24596 8974 24624 9302
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24596 8566 24624 8910
rect 24584 8560 24636 8566
rect 24584 8502 24636 8508
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24320 7954 24348 8434
rect 24596 8090 24624 8502
rect 24872 8362 24900 9454
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 9110 24992 9318
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 25240 8906 25268 9454
rect 25424 9042 25452 9454
rect 25884 9178 25912 10066
rect 26344 9994 26372 10202
rect 26332 9988 26384 9994
rect 26332 9930 26384 9936
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 25976 9382 26004 9590
rect 26332 9580 26384 9586
rect 26160 9540 26332 9568
rect 26160 9450 26188 9540
rect 26332 9522 26384 9528
rect 26148 9444 26200 9450
rect 26148 9386 26200 9392
rect 26240 9444 26292 9450
rect 26240 9386 26292 9392
rect 25964 9376 26016 9382
rect 25964 9318 26016 9324
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25976 9110 26004 9318
rect 25964 9104 26016 9110
rect 25964 9046 26016 9052
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25240 8362 25268 8842
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25608 8498 25636 8774
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25792 8362 25820 8774
rect 26160 8634 26188 9386
rect 26252 9110 26280 9386
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26240 9104 26292 9110
rect 26240 9046 26292 9052
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25780 8356 25832 8362
rect 25780 8298 25832 8304
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24308 7948 24360 7954
rect 24308 7890 24360 7896
rect 25240 7818 25268 8298
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25608 8022 25636 8230
rect 25596 8016 25648 8022
rect 25596 7958 25648 7964
rect 26252 7886 26280 9046
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26344 8430 26372 8978
rect 26436 8906 26464 9318
rect 26528 9110 26556 19887
rect 27988 19858 28040 19864
rect 28000 19718 28028 19858
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27988 19712 28040 19718
rect 27988 19654 28040 19660
rect 26984 19612 27292 19621
rect 26984 19610 26990 19612
rect 27046 19610 27070 19612
rect 27126 19610 27150 19612
rect 27206 19610 27230 19612
rect 27286 19610 27292 19612
rect 27046 19558 27048 19610
rect 27228 19558 27230 19610
rect 26984 19556 26990 19558
rect 27046 19556 27070 19558
rect 27126 19556 27150 19558
rect 27206 19556 27230 19558
rect 27286 19556 27292 19558
rect 26984 19547 27292 19556
rect 27448 19310 27476 19654
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26976 19304 27028 19310
rect 26976 19246 27028 19252
rect 27436 19304 27488 19310
rect 27436 19246 27488 19252
rect 26712 18834 26740 19246
rect 26792 19236 26844 19242
rect 26792 19178 26844 19184
rect 26804 18834 26832 19178
rect 26896 18970 26924 19246
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 26700 18828 26752 18834
rect 26700 18770 26752 18776
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 26804 18222 26832 18770
rect 26988 18612 27016 19246
rect 27644 19068 27952 19077
rect 27644 19066 27650 19068
rect 27706 19066 27730 19068
rect 27786 19066 27810 19068
rect 27866 19066 27890 19068
rect 27946 19066 27952 19068
rect 27706 19014 27708 19066
rect 27888 19014 27890 19066
rect 27644 19012 27650 19014
rect 27706 19012 27730 19014
rect 27786 19012 27810 19014
rect 27866 19012 27890 19014
rect 27946 19012 27952 19014
rect 27644 19003 27952 19012
rect 27436 18964 27488 18970
rect 27436 18906 27488 18912
rect 26896 18584 27016 18612
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 26620 17814 26648 18158
rect 26608 17808 26660 17814
rect 26608 17750 26660 17756
rect 26896 16998 26924 18584
rect 26984 18524 27292 18533
rect 26984 18522 26990 18524
rect 27046 18522 27070 18524
rect 27126 18522 27150 18524
rect 27206 18522 27230 18524
rect 27286 18522 27292 18524
rect 27046 18470 27048 18522
rect 27228 18470 27230 18522
rect 26984 18468 26990 18470
rect 27046 18468 27070 18470
rect 27126 18468 27150 18470
rect 27206 18468 27230 18470
rect 27286 18468 27292 18470
rect 26984 18459 27292 18468
rect 27448 18154 27476 18906
rect 28000 18902 28028 19654
rect 28092 19514 28120 20742
rect 29196 20058 29224 21422
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 30484 21010 30512 21286
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 29276 20936 29328 20942
rect 29276 20878 29328 20884
rect 29288 20398 29316 20878
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29380 20602 29408 20742
rect 29368 20596 29420 20602
rect 29368 20538 29420 20544
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 28816 19916 28868 19922
rect 28816 19858 28868 19864
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28828 19378 28856 19858
rect 28816 19372 28868 19378
rect 28816 19314 28868 19320
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 27988 18896 28040 18902
rect 27526 18864 27582 18873
rect 27988 18838 28040 18844
rect 27526 18799 27528 18808
rect 27580 18799 27582 18808
rect 27712 18828 27764 18834
rect 27528 18770 27580 18776
rect 27712 18770 27764 18776
rect 27804 18828 27856 18834
rect 27804 18770 27856 18776
rect 28080 18828 28132 18834
rect 28080 18770 28132 18776
rect 28632 18828 28684 18834
rect 28632 18770 28684 18776
rect 27724 18426 27752 18770
rect 27816 18630 27844 18770
rect 27804 18624 27856 18630
rect 27804 18566 27856 18572
rect 28092 18426 28120 18770
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 28080 18420 28132 18426
rect 28080 18362 28132 18368
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 28356 18352 28408 18358
rect 28356 18294 28408 18300
rect 27632 18170 27660 18294
rect 28368 18222 28396 18294
rect 27540 18154 27660 18170
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 28644 18154 28672 18770
rect 29104 18698 29132 19246
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29092 18692 29144 18698
rect 29092 18634 29144 18640
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 27436 18148 27488 18154
rect 27436 18090 27488 18096
rect 27540 18148 27672 18154
rect 27540 18142 27620 18148
rect 27540 17762 27568 18142
rect 27620 18090 27672 18096
rect 28632 18148 28684 18154
rect 28632 18090 28684 18096
rect 28078 18048 28134 18057
rect 27644 17980 27952 17989
rect 28078 17983 28134 17992
rect 27644 17978 27650 17980
rect 27706 17978 27730 17980
rect 27786 17978 27810 17980
rect 27866 17978 27890 17980
rect 27946 17978 27952 17980
rect 27706 17926 27708 17978
rect 27888 17926 27890 17978
rect 27644 17924 27650 17926
rect 27706 17924 27730 17926
rect 27786 17924 27810 17926
rect 27866 17924 27890 17926
rect 27946 17924 27952 17926
rect 27644 17915 27952 17924
rect 27540 17734 27660 17762
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 26984 17436 27292 17445
rect 26984 17434 26990 17436
rect 27046 17434 27070 17436
rect 27126 17434 27150 17436
rect 27206 17434 27230 17436
rect 27286 17434 27292 17436
rect 27046 17382 27048 17434
rect 27228 17382 27230 17434
rect 26984 17380 26990 17382
rect 27046 17380 27070 17382
rect 27126 17380 27150 17382
rect 27206 17380 27230 17382
rect 27286 17380 27292 17382
rect 26984 17371 27292 17380
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26606 16824 26662 16833
rect 26606 16759 26662 16768
rect 26620 16114 26648 16759
rect 26792 16652 26844 16658
rect 26712 16612 26792 16640
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26608 15972 26660 15978
rect 26608 15914 26660 15920
rect 26620 15638 26648 15914
rect 26608 15632 26660 15638
rect 26608 15574 26660 15580
rect 26712 15162 26740 16612
rect 26896 16640 26924 16934
rect 27448 16658 27476 17274
rect 26844 16612 26924 16640
rect 27436 16652 27488 16658
rect 26792 16594 26844 16600
rect 27436 16594 27488 16600
rect 26984 16348 27292 16357
rect 26984 16346 26990 16348
rect 27046 16346 27070 16348
rect 27126 16346 27150 16348
rect 27206 16346 27230 16348
rect 27286 16346 27292 16348
rect 27046 16294 27048 16346
rect 27228 16294 27230 16346
rect 26984 16292 26990 16294
rect 27046 16292 27070 16294
rect 27126 16292 27150 16294
rect 27206 16292 27230 16294
rect 27286 16292 27292 16294
rect 26984 16283 27292 16292
rect 26792 16176 26844 16182
rect 26792 16118 26844 16124
rect 26700 15156 26752 15162
rect 26620 15116 26700 15144
rect 26620 14550 26648 15116
rect 26700 15098 26752 15104
rect 26804 15094 26832 16118
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 26984 15260 27292 15269
rect 26984 15258 26990 15260
rect 27046 15258 27070 15260
rect 27126 15258 27150 15260
rect 27206 15258 27230 15260
rect 27286 15258 27292 15260
rect 27046 15206 27048 15258
rect 27228 15206 27230 15258
rect 26984 15204 26990 15206
rect 27046 15204 27070 15206
rect 27126 15204 27150 15206
rect 27206 15204 27230 15206
rect 27286 15204 27292 15206
rect 26984 15195 27292 15204
rect 26792 15088 26844 15094
rect 26792 15030 26844 15036
rect 27160 15088 27212 15094
rect 27160 15030 27212 15036
rect 26700 15020 26752 15026
rect 26700 14962 26752 14968
rect 26608 14544 26660 14550
rect 26608 14486 26660 14492
rect 26712 14074 26740 14962
rect 26804 14482 26832 15030
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26700 14068 26752 14074
rect 26700 14010 26752 14016
rect 26804 13530 26832 14282
rect 26896 14074 26924 14894
rect 27172 14618 27200 15030
rect 27252 14816 27304 14822
rect 27252 14758 27304 14764
rect 27160 14612 27212 14618
rect 27160 14554 27212 14560
rect 27172 14482 27200 14554
rect 27264 14482 27292 14758
rect 26976 14476 27028 14482
rect 26976 14418 27028 14424
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27252 14476 27304 14482
rect 27252 14418 27304 14424
rect 26988 14385 27016 14418
rect 26974 14376 27030 14385
rect 26974 14311 27030 14320
rect 26984 14172 27292 14181
rect 26984 14170 26990 14172
rect 27046 14170 27070 14172
rect 27126 14170 27150 14172
rect 27206 14170 27230 14172
rect 27286 14170 27292 14172
rect 27046 14118 27048 14170
rect 27228 14118 27230 14170
rect 26984 14116 26990 14118
rect 27046 14116 27070 14118
rect 27126 14116 27150 14118
rect 27206 14116 27230 14118
rect 27286 14116 27292 14118
rect 26984 14107 27292 14116
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 27356 13870 27384 15914
rect 27448 15094 27476 16594
rect 27540 16454 27568 17614
rect 27632 17270 27660 17734
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 27632 17066 27660 17206
rect 27620 17060 27672 17066
rect 27620 17002 27672 17008
rect 27644 16892 27952 16901
rect 27644 16890 27650 16892
rect 27706 16890 27730 16892
rect 27786 16890 27810 16892
rect 27866 16890 27890 16892
rect 27946 16890 27952 16892
rect 27706 16838 27708 16890
rect 27888 16838 27890 16890
rect 27644 16836 27650 16838
rect 27706 16836 27730 16838
rect 27786 16836 27810 16838
rect 27866 16836 27890 16838
rect 27946 16836 27952 16838
rect 27644 16827 27952 16836
rect 28000 16658 28028 17478
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27988 16448 28040 16454
rect 27988 16390 28040 16396
rect 27644 15804 27952 15813
rect 27644 15802 27650 15804
rect 27706 15802 27730 15804
rect 27786 15802 27810 15804
rect 27866 15802 27890 15804
rect 27946 15802 27952 15804
rect 27706 15750 27708 15802
rect 27888 15750 27890 15802
rect 27644 15748 27650 15750
rect 27706 15748 27730 15750
rect 27786 15748 27810 15750
rect 27866 15748 27890 15750
rect 27946 15748 27952 15750
rect 27644 15739 27952 15748
rect 28000 15570 28028 16390
rect 27988 15564 28040 15570
rect 27988 15506 28040 15512
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 28000 14958 28028 15506
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27988 14952 28040 14958
rect 27988 14894 28040 14900
rect 27448 14618 27476 14894
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27540 14482 27568 14758
rect 27644 14716 27952 14725
rect 27644 14714 27650 14716
rect 27706 14714 27730 14716
rect 27786 14714 27810 14716
rect 27866 14714 27890 14716
rect 27946 14714 27952 14716
rect 27706 14662 27708 14714
rect 27888 14662 27890 14714
rect 27644 14660 27650 14662
rect 27706 14660 27730 14662
rect 27786 14660 27810 14662
rect 27866 14660 27890 14662
rect 27946 14660 27952 14662
rect 27644 14651 27952 14660
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27804 14476 27856 14482
rect 27804 14418 27856 14424
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27724 13938 27752 14214
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27816 13870 27844 14418
rect 27896 14408 27948 14414
rect 27896 14350 27948 14356
rect 27908 13870 27936 14350
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27896 13864 27948 13870
rect 27896 13806 27948 13812
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26988 13394 27016 13670
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26984 13084 27292 13093
rect 26984 13082 26990 13084
rect 27046 13082 27070 13084
rect 27126 13082 27150 13084
rect 27206 13082 27230 13084
rect 27286 13082 27292 13084
rect 27046 13030 27048 13082
rect 27228 13030 27230 13082
rect 26984 13028 26990 13030
rect 27046 13028 27070 13030
rect 27126 13028 27150 13030
rect 27206 13028 27230 13030
rect 27286 13028 27292 13030
rect 26984 13019 27292 13028
rect 27356 12374 27384 13806
rect 27644 13628 27952 13637
rect 27644 13626 27650 13628
rect 27706 13626 27730 13628
rect 27786 13626 27810 13628
rect 27866 13626 27890 13628
rect 27946 13626 27952 13628
rect 27706 13574 27708 13626
rect 27888 13574 27890 13626
rect 27644 13572 27650 13574
rect 27706 13572 27730 13574
rect 27786 13572 27810 13574
rect 27866 13572 27890 13574
rect 27946 13572 27952 13574
rect 27644 13563 27952 13572
rect 28000 13462 28028 14282
rect 27988 13456 28040 13462
rect 27988 13398 28040 13404
rect 27644 12540 27952 12549
rect 27644 12538 27650 12540
rect 27706 12538 27730 12540
rect 27786 12538 27810 12540
rect 27866 12538 27890 12540
rect 27946 12538 27952 12540
rect 27706 12486 27708 12538
rect 27888 12486 27890 12538
rect 27644 12484 27650 12486
rect 27706 12484 27730 12486
rect 27786 12484 27810 12486
rect 27866 12484 27890 12486
rect 27946 12484 27952 12486
rect 27644 12475 27952 12484
rect 27344 12368 27396 12374
rect 27344 12310 27396 12316
rect 26984 11996 27292 12005
rect 26984 11994 26990 11996
rect 27046 11994 27070 11996
rect 27126 11994 27150 11996
rect 27206 11994 27230 11996
rect 27286 11994 27292 11996
rect 27046 11942 27048 11994
rect 27228 11942 27230 11994
rect 26984 11940 26990 11942
rect 27046 11940 27070 11942
rect 27126 11940 27150 11942
rect 27206 11940 27230 11942
rect 27286 11940 27292 11942
rect 26984 11931 27292 11940
rect 27356 11762 27384 12310
rect 28092 11898 28120 17983
rect 28172 17876 28224 17882
rect 28172 17818 28224 17824
rect 28184 17338 28212 17818
rect 28540 17808 28592 17814
rect 28540 17750 28592 17756
rect 28356 17604 28408 17610
rect 28356 17546 28408 17552
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 28184 17134 28212 17274
rect 28264 17264 28316 17270
rect 28264 17206 28316 17212
rect 28172 17128 28224 17134
rect 28172 17070 28224 17076
rect 28172 16992 28224 16998
rect 28172 16934 28224 16940
rect 28184 16046 28212 16934
rect 28172 16040 28224 16046
rect 28172 15982 28224 15988
rect 28276 15706 28304 17206
rect 28368 17134 28396 17546
rect 28552 17338 28580 17750
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 28356 17128 28408 17134
rect 28356 17070 28408 17076
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 28276 14634 28304 15642
rect 28448 15564 28500 15570
rect 28552 15552 28580 17274
rect 28644 16250 28672 17614
rect 28632 16244 28684 16250
rect 28632 16186 28684 16192
rect 28500 15524 28580 15552
rect 28448 15506 28500 15512
rect 28356 15088 28408 15094
rect 28356 15030 28408 15036
rect 28184 14606 28304 14634
rect 28184 13394 28212 14606
rect 28262 14512 28318 14521
rect 28368 14482 28396 15030
rect 28460 14890 28488 15506
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28448 14884 28500 14890
rect 28448 14826 28500 14832
rect 28262 14447 28264 14456
rect 28316 14447 28318 14456
rect 28356 14476 28408 14482
rect 28264 14418 28316 14424
rect 28356 14418 28408 14424
rect 28368 14385 28396 14418
rect 28354 14376 28410 14385
rect 28354 14311 28410 14320
rect 28262 13968 28318 13977
rect 28262 13903 28318 13912
rect 28276 13870 28304 13903
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 28460 12850 28488 14826
rect 28552 14482 28580 15302
rect 28632 14952 28684 14958
rect 28632 14894 28684 14900
rect 28644 14482 28672 14894
rect 28540 14476 28592 14482
rect 28540 14418 28592 14424
rect 28632 14476 28684 14482
rect 28632 14418 28684 14424
rect 28644 13530 28672 14418
rect 28828 13734 28856 18566
rect 29104 18442 29132 18634
rect 29012 18414 29132 18442
rect 28908 18148 28960 18154
rect 28908 18090 28960 18096
rect 28920 17270 28948 18090
rect 29012 17882 29040 18414
rect 29196 18358 29224 18702
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 29184 18352 29236 18358
rect 29184 18294 29236 18300
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 29012 17134 29040 17478
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 29104 17082 29132 18294
rect 29288 17882 29316 20334
rect 29460 20324 29512 20330
rect 29460 20266 29512 20272
rect 29472 20058 29500 20266
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29644 20256 29696 20262
rect 29644 20198 29696 20204
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29564 19922 29592 20198
rect 29656 19990 29684 20198
rect 29644 19984 29696 19990
rect 29644 19926 29696 19932
rect 29552 19916 29604 19922
rect 29552 19858 29604 19864
rect 29368 19848 29420 19854
rect 29368 19790 29420 19796
rect 29380 19530 29408 19790
rect 29380 19502 29592 19530
rect 29380 19310 29408 19502
rect 29460 19440 29512 19446
rect 29460 19382 29512 19388
rect 29472 19310 29500 19382
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29460 19304 29512 19310
rect 29460 19246 29512 19252
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29380 18970 29408 19110
rect 29472 18970 29500 19246
rect 29564 18970 29592 19502
rect 29368 18964 29420 18970
rect 29368 18906 29420 18912
rect 29460 18964 29512 18970
rect 29460 18906 29512 18912
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29472 18834 29500 18906
rect 29460 18828 29512 18834
rect 29460 18770 29512 18776
rect 29472 18714 29500 18770
rect 29380 18686 29500 18714
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29380 17882 29408 18686
rect 29564 18426 29592 18702
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29656 18290 29684 19926
rect 29828 19916 29880 19922
rect 29828 19858 29880 19864
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29748 19174 29776 19654
rect 29840 19514 29868 19858
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 29828 19508 29880 19514
rect 29828 19450 29880 19456
rect 29932 19446 29960 19654
rect 29920 19440 29972 19446
rect 29920 19382 29972 19388
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 30288 19304 30340 19310
rect 30288 19246 30340 19252
rect 30380 19304 30432 19310
rect 30380 19246 30432 19252
rect 29736 19168 29788 19174
rect 29736 19110 29788 19116
rect 29840 18970 29868 19246
rect 29920 19236 29972 19242
rect 29920 19178 29972 19184
rect 29932 18970 29960 19178
rect 29736 18964 29788 18970
rect 29736 18906 29788 18912
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 29920 18964 29972 18970
rect 29920 18906 29972 18912
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29460 18216 29512 18222
rect 29460 18158 29512 18164
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29368 17876 29420 17882
rect 29368 17818 29420 17824
rect 29380 17202 29408 17818
rect 29472 17728 29500 18158
rect 29564 17898 29592 18226
rect 29656 18154 29684 18226
rect 29644 18148 29696 18154
rect 29644 18090 29696 18096
rect 29564 17870 29684 17898
rect 29552 17740 29604 17746
rect 29472 17700 29552 17728
rect 29472 17338 29500 17700
rect 29552 17682 29604 17688
rect 29656 17678 29684 17870
rect 29644 17672 29696 17678
rect 29644 17614 29696 17620
rect 29552 17604 29604 17610
rect 29552 17546 29604 17552
rect 29460 17332 29512 17338
rect 29460 17274 29512 17280
rect 29368 17196 29420 17202
rect 29368 17138 29420 17144
rect 29104 17054 29224 17082
rect 29092 16992 29144 16998
rect 29092 16934 29144 16940
rect 29104 16726 29132 16934
rect 29092 16720 29144 16726
rect 29092 16662 29144 16668
rect 29196 16130 29224 17054
rect 29472 16726 29500 17274
rect 29460 16720 29512 16726
rect 29460 16662 29512 16668
rect 29368 16652 29420 16658
rect 29368 16594 29420 16600
rect 29104 16102 29224 16130
rect 29104 16046 29132 16102
rect 29380 16046 29408 16594
rect 29564 16454 29592 17546
rect 29656 16590 29684 17614
rect 29644 16584 29696 16590
rect 29644 16526 29696 16532
rect 29552 16448 29604 16454
rect 29552 16390 29604 16396
rect 29564 16114 29592 16390
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29092 16040 29144 16046
rect 29276 16040 29328 16046
rect 29092 15982 29144 15988
rect 29196 16000 29276 16028
rect 29104 15706 29132 15982
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 29196 15570 29224 16000
rect 29276 15982 29328 15988
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29288 15570 29316 15642
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29276 15564 29328 15570
rect 29276 15506 29328 15512
rect 29012 15162 29040 15506
rect 29104 15434 29132 15506
rect 29092 15428 29144 15434
rect 29092 15370 29144 15376
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29012 14414 29040 14962
rect 29104 14822 29132 15370
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 29196 14550 29224 15506
rect 29288 15094 29316 15506
rect 29276 15088 29328 15094
rect 29276 15030 29328 15036
rect 29276 14816 29328 14822
rect 29276 14758 29328 14764
rect 29184 14544 29236 14550
rect 29184 14486 29236 14492
rect 29196 14414 29224 14486
rect 29000 14408 29052 14414
rect 29000 14350 29052 14356
rect 29184 14408 29236 14414
rect 29184 14350 29236 14356
rect 29288 14346 29316 14758
rect 29380 14618 29408 15982
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29472 15162 29500 15506
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 29564 14958 29592 16050
rect 29748 15026 29776 18906
rect 30208 18873 30236 19246
rect 30300 18902 30328 19246
rect 30392 18970 30420 19246
rect 30656 19168 30708 19174
rect 30656 19110 30708 19116
rect 30380 18964 30432 18970
rect 30380 18906 30432 18912
rect 30288 18896 30340 18902
rect 30194 18864 30250 18873
rect 30104 18828 30156 18834
rect 30288 18838 30340 18844
rect 30194 18799 30196 18808
rect 30104 18770 30156 18776
rect 30248 18799 30250 18808
rect 30196 18770 30248 18776
rect 30116 18426 30144 18770
rect 30668 18698 30696 19110
rect 30472 18692 30524 18698
rect 30472 18634 30524 18640
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30288 16788 30340 16794
rect 30288 16730 30340 16736
rect 29920 16720 29972 16726
rect 29920 16662 29972 16668
rect 29932 16046 29960 16662
rect 30300 16590 30328 16730
rect 30288 16584 30340 16590
rect 30288 16526 30340 16532
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29920 15904 29972 15910
rect 29920 15846 29972 15852
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29736 15020 29788 15026
rect 29736 14962 29788 14968
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29368 14612 29420 14618
rect 29368 14554 29420 14560
rect 29276 14340 29328 14346
rect 29276 14282 29328 14288
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 28816 13728 28868 13734
rect 28816 13670 28868 13676
rect 28632 13524 28684 13530
rect 28632 13466 28684 13472
rect 28448 12844 28500 12850
rect 28448 12786 28500 12792
rect 28828 12714 28856 13670
rect 28908 13388 28960 13394
rect 28908 13330 28960 13336
rect 28816 12708 28868 12714
rect 28816 12650 28868 12656
rect 28920 12306 28948 13330
rect 29012 12782 29040 14214
rect 29104 13870 29132 14214
rect 29288 14074 29316 14282
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 29196 12986 29224 13942
rect 29288 13258 29316 14010
rect 29380 13870 29408 14554
rect 29656 14414 29684 14962
rect 29932 14890 29960 15846
rect 30484 14958 30512 18634
rect 30656 17536 30708 17542
rect 30656 17478 30708 17484
rect 30668 17202 30696 17478
rect 30748 17332 30800 17338
rect 30748 17274 30800 17280
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30760 16658 30788 17274
rect 31024 17128 31076 17134
rect 31024 17070 31076 17076
rect 30564 16652 30616 16658
rect 30564 16594 30616 16600
rect 30748 16652 30800 16658
rect 30748 16594 30800 16600
rect 30576 16250 30604 16594
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30564 15088 30616 15094
rect 30564 15030 30616 15036
rect 30472 14952 30524 14958
rect 30472 14894 30524 14900
rect 29920 14884 29972 14890
rect 29920 14826 29972 14832
rect 30196 14884 30248 14890
rect 30196 14826 30248 14832
rect 29828 14816 29880 14822
rect 29828 14758 29880 14764
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29460 13932 29512 13938
rect 29460 13874 29512 13880
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 29472 13462 29500 13874
rect 29840 13870 29868 14758
rect 29552 13864 29604 13870
rect 29552 13806 29604 13812
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29564 13530 29592 13806
rect 29932 13802 29960 14826
rect 30104 14272 30156 14278
rect 30104 14214 30156 14220
rect 29920 13796 29972 13802
rect 29920 13738 29972 13744
rect 29552 13524 29604 13530
rect 29552 13466 29604 13472
rect 29460 13456 29512 13462
rect 29460 13398 29512 13404
rect 29276 13252 29328 13258
rect 29276 13194 29328 13200
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 30116 12850 30144 14214
rect 30208 13977 30236 14826
rect 30576 14482 30604 15030
rect 30668 14958 30696 15302
rect 30656 14952 30708 14958
rect 30656 14894 30708 14900
rect 30840 14952 30892 14958
rect 30840 14894 30892 14900
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30484 14074 30512 14418
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30194 13968 30250 13977
rect 30194 13903 30250 13912
rect 30852 13530 30880 14894
rect 30932 14612 30984 14618
rect 30932 14554 30984 14560
rect 30944 14074 30972 14554
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 30944 13326 30972 14010
rect 31036 13870 31064 17070
rect 31024 13864 31076 13870
rect 31024 13806 31076 13812
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 31036 12306 31064 13806
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31128 13394 31156 13670
rect 31116 13388 31168 13394
rect 31116 13330 31168 13336
rect 28908 12300 28960 12306
rect 28908 12242 28960 12248
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 31024 12300 31076 12306
rect 31024 12242 31076 12248
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 28184 11694 28212 12038
rect 28828 11898 28856 12174
rect 29184 12096 29236 12102
rect 29184 12038 29236 12044
rect 28816 11892 28868 11898
rect 28816 11834 28868 11840
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 26884 11688 26936 11694
rect 28172 11688 28224 11694
rect 26884 11630 26936 11636
rect 27066 11656 27122 11665
rect 26804 11354 26832 11630
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 26620 9518 26648 9590
rect 26712 9518 26740 9658
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26804 9466 26832 10066
rect 26896 9654 26924 11630
rect 28172 11630 28224 11636
rect 27066 11591 27068 11600
rect 27120 11591 27122 11600
rect 27528 11620 27580 11626
rect 27068 11562 27120 11568
rect 27528 11562 27580 11568
rect 27540 11200 27568 11562
rect 27644 11452 27952 11461
rect 27644 11450 27650 11452
rect 27706 11450 27730 11452
rect 27786 11450 27810 11452
rect 27866 11450 27890 11452
rect 27946 11450 27952 11452
rect 27706 11398 27708 11450
rect 27888 11398 27890 11450
rect 27644 11396 27650 11398
rect 27706 11396 27730 11398
rect 27786 11396 27810 11398
rect 27866 11396 27890 11398
rect 27946 11396 27952 11398
rect 27644 11387 27952 11396
rect 28184 11218 28212 11630
rect 28540 11552 28592 11558
rect 28540 11494 28592 11500
rect 28172 11212 28224 11218
rect 27540 11172 27660 11200
rect 27632 11082 27660 11172
rect 28172 11154 28224 11160
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 28552 11014 28580 11494
rect 28828 11354 28856 11834
rect 29196 11762 29224 12038
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 29092 11620 29144 11626
rect 29092 11562 29144 11568
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 29104 11218 29132 11562
rect 28908 11212 28960 11218
rect 28908 11154 28960 11160
rect 29092 11212 29144 11218
rect 29092 11154 29144 11160
rect 28540 11008 28592 11014
rect 28540 10950 28592 10956
rect 26984 10908 27292 10917
rect 26984 10906 26990 10908
rect 27046 10906 27070 10908
rect 27126 10906 27150 10908
rect 27206 10906 27230 10908
rect 27286 10906 27292 10908
rect 27046 10854 27048 10906
rect 27228 10854 27230 10906
rect 26984 10852 26990 10854
rect 27046 10852 27070 10854
rect 27126 10852 27150 10854
rect 27206 10852 27230 10854
rect 27286 10852 27292 10854
rect 26984 10843 27292 10852
rect 28920 10606 28948 11154
rect 29564 11082 29592 12242
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 29736 12096 29788 12102
rect 29736 12038 29788 12044
rect 29920 12096 29972 12102
rect 29920 12038 29972 12044
rect 29748 11694 29776 12038
rect 29736 11688 29788 11694
rect 29736 11630 29788 11636
rect 29932 11286 29960 12038
rect 30748 11552 30800 11558
rect 30748 11494 30800 11500
rect 29920 11280 29972 11286
rect 29920 11222 29972 11228
rect 30760 11218 30788 11494
rect 30012 11212 30064 11218
rect 30012 11154 30064 11160
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 29552 11076 29604 11082
rect 29552 11018 29604 11024
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 29012 10674 29040 10950
rect 29564 10742 29592 11018
rect 30024 10810 30052 11154
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 28908 10600 28960 10606
rect 28908 10542 28960 10548
rect 28632 10464 28684 10470
rect 28632 10406 28684 10412
rect 27644 10364 27952 10373
rect 27644 10362 27650 10364
rect 27706 10362 27730 10364
rect 27786 10362 27810 10364
rect 27866 10362 27890 10364
rect 27946 10362 27952 10364
rect 27706 10310 27708 10362
rect 27888 10310 27890 10362
rect 27644 10308 27650 10310
rect 27706 10308 27730 10310
rect 27786 10308 27810 10310
rect 27866 10308 27890 10310
rect 27946 10308 27952 10310
rect 27644 10299 27952 10308
rect 28644 10130 28672 10406
rect 28632 10124 28684 10130
rect 28632 10066 28684 10072
rect 28816 10124 28868 10130
rect 28816 10066 28868 10072
rect 26984 9820 27292 9829
rect 26984 9818 26990 9820
rect 27046 9818 27070 9820
rect 27126 9818 27150 9820
rect 27206 9818 27230 9820
rect 27286 9818 27292 9820
rect 27046 9766 27048 9818
rect 27228 9766 27230 9818
rect 26984 9764 26990 9766
rect 27046 9764 27070 9766
rect 27126 9764 27150 9766
rect 27206 9764 27230 9766
rect 27286 9764 27292 9766
rect 26984 9755 27292 9764
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 26884 9512 26936 9518
rect 26804 9460 26884 9466
rect 26804 9454 26936 9460
rect 26620 9382 26648 9454
rect 26608 9376 26660 9382
rect 26608 9318 26660 9324
rect 26712 9178 26740 9454
rect 26804 9438 26924 9454
rect 27080 9450 27108 9590
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27068 9444 27120 9450
rect 27068 9386 27120 9392
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26516 9104 26568 9110
rect 26516 9046 26568 9052
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26792 8832 26844 8838
rect 26792 8774 26844 8780
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26804 7954 26832 8774
rect 26984 8732 27292 8741
rect 26984 8730 26990 8732
rect 27046 8730 27070 8732
rect 27126 8730 27150 8732
rect 27206 8730 27230 8732
rect 27286 8730 27292 8732
rect 27046 8678 27048 8730
rect 27228 8678 27230 8730
rect 26984 8676 26990 8678
rect 27046 8676 27070 8678
rect 27126 8676 27150 8678
rect 27206 8676 27230 8678
rect 27286 8676 27292 8678
rect 26984 8667 27292 8676
rect 27356 8430 27384 9522
rect 28092 9518 28120 9590
rect 28184 9518 28212 9658
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 28172 9512 28224 9518
rect 28172 9454 28224 9460
rect 28092 9382 28120 9454
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 27644 9276 27952 9285
rect 27644 9274 27650 9276
rect 27706 9274 27730 9276
rect 27786 9274 27810 9276
rect 27866 9274 27890 9276
rect 27946 9274 27952 9276
rect 27706 9222 27708 9274
rect 27888 9222 27890 9274
rect 27644 9220 27650 9222
rect 27706 9220 27730 9222
rect 27786 9220 27810 9222
rect 27866 9220 27890 9222
rect 27946 9220 27952 9222
rect 27644 9211 27952 9220
rect 28184 9042 28212 9454
rect 28448 9444 28500 9450
rect 28448 9386 28500 9392
rect 28460 9178 28488 9386
rect 28828 9382 28856 10066
rect 28920 10062 28948 10542
rect 30116 10266 30144 10610
rect 30760 10538 30788 11154
rect 30944 10810 30972 12174
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 30748 10532 30800 10538
rect 30748 10474 30800 10480
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 30288 10260 30340 10266
rect 30288 10202 30340 10208
rect 30196 10124 30248 10130
rect 30196 10066 30248 10072
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28448 9172 28500 9178
rect 28448 9114 28500 9120
rect 28172 9036 28224 9042
rect 28172 8978 28224 8984
rect 28184 8634 28212 8978
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28828 8430 28856 9318
rect 29012 8498 29040 9590
rect 30116 9518 30144 9862
rect 30208 9586 30236 10066
rect 30196 9580 30248 9586
rect 30196 9522 30248 9528
rect 30300 9518 30328 10202
rect 31036 10130 31064 12242
rect 31116 11688 31168 11694
rect 31116 11630 31168 11636
rect 31128 11354 31156 11630
rect 31116 11348 31168 11354
rect 31116 11290 31168 11296
rect 31128 10606 31156 11290
rect 31300 11008 31352 11014
rect 31300 10950 31352 10956
rect 31312 10606 31340 10950
rect 31116 10600 31168 10606
rect 31116 10542 31168 10548
rect 31300 10600 31352 10606
rect 31300 10542 31352 10548
rect 31024 10124 31076 10130
rect 31024 10066 31076 10072
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 30104 9512 30156 9518
rect 30104 9454 30156 9460
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 29104 9110 29132 9318
rect 29932 9178 29960 9454
rect 29920 9172 29972 9178
rect 29920 9114 29972 9120
rect 29092 9104 29144 9110
rect 29092 9046 29144 9052
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 30024 8634 30052 8978
rect 30012 8628 30064 8634
rect 30012 8570 30064 8576
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 27356 7954 27384 8366
rect 27528 8356 27580 8362
rect 27528 8298 27580 8304
rect 27540 8090 27568 8298
rect 27644 8188 27952 8197
rect 27644 8186 27650 8188
rect 27706 8186 27730 8188
rect 27786 8186 27810 8188
rect 27866 8186 27890 8188
rect 27946 8186 27952 8188
rect 27706 8134 27708 8186
rect 27888 8134 27890 8186
rect 27644 8132 27650 8134
rect 27706 8132 27730 8134
rect 27786 8132 27810 8134
rect 27866 8132 27890 8134
rect 27946 8132 27952 8134
rect 27644 8123 27952 8132
rect 28000 8090 28028 8366
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 25228 7812 25280 7818
rect 25228 7754 25280 7760
rect 26984 7644 27292 7653
rect 26984 7642 26990 7644
rect 27046 7642 27070 7644
rect 27126 7642 27150 7644
rect 27206 7642 27230 7644
rect 27286 7642 27292 7644
rect 27046 7590 27048 7642
rect 27228 7590 27230 7642
rect 26984 7588 26990 7590
rect 27046 7588 27070 7590
rect 27126 7588 27150 7590
rect 27206 7588 27230 7590
rect 27286 7588 27292 7590
rect 26984 7579 27292 7588
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 27356 7342 27384 7890
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 27344 7336 27396 7342
rect 27344 7278 27396 7284
rect 30380 7336 30432 7342
rect 30380 7278 30432 7284
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22480 5166 22508 6190
rect 23400 6186 23428 6598
rect 24872 6390 24900 7278
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 26252 7018 26280 7142
rect 26068 6990 26280 7018
rect 26068 6662 26096 6990
rect 26436 6866 26464 7142
rect 26240 6860 26292 6866
rect 26240 6802 26292 6808
rect 26424 6860 26476 6866
rect 26976 6860 27028 6866
rect 26424 6802 26476 6808
rect 26896 6820 26976 6848
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 26056 6656 26108 6662
rect 26056 6598 26108 6604
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 23388 6180 23440 6186
rect 23388 6122 23440 6128
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 22664 5370 22692 5714
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22756 5234 22784 5714
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22008 5102 22060 5108
rect 22112 5120 22324 5148
rect 22468 5160 22520 5166
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21652 4826 21680 4966
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21100 4010 21128 4626
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21560 4282 21588 4422
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21560 4078 21588 4218
rect 21652 4146 21680 4762
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21088 4004 21140 4010
rect 21088 3946 21140 3952
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19720 2514 19748 3334
rect 19812 2582 19840 3538
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20272 2990 20300 3334
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20364 2774 20392 3538
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 19870 2748 20178 2757
rect 19870 2746 19876 2748
rect 19932 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20178 2748
rect 19932 2694 19934 2746
rect 20114 2694 20116 2746
rect 19870 2692 19876 2694
rect 19932 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20178 2694
rect 19870 2683 20178 2692
rect 20272 2746 20392 2774
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 18248 1970 18276 2450
rect 19210 2204 19518 2213
rect 19210 2202 19216 2204
rect 19272 2202 19296 2204
rect 19352 2202 19376 2204
rect 19432 2202 19456 2204
rect 19512 2202 19518 2204
rect 19272 2150 19274 2202
rect 19454 2150 19456 2202
rect 19210 2148 19216 2150
rect 19272 2148 19296 2150
rect 19352 2148 19376 2150
rect 19432 2148 19456 2150
rect 19512 2148 19518 2150
rect 19210 2139 19518 2148
rect 19708 2032 19760 2038
rect 19708 1974 19760 1980
rect 18236 1964 18288 1970
rect 18236 1906 18288 1912
rect 17776 1896 17828 1902
rect 17776 1838 17828 1844
rect 17788 1766 17816 1838
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 17776 1760 17828 1766
rect 17776 1702 17828 1708
rect 18328 1760 18380 1766
rect 18328 1702 18380 1708
rect 19432 1760 19484 1766
rect 19432 1702 19484 1708
rect 16764 1556 16816 1562
rect 16764 1498 16816 1504
rect 17604 1494 17632 1702
rect 17592 1488 17644 1494
rect 17592 1430 17644 1436
rect 16488 1420 16540 1426
rect 16488 1362 16540 1368
rect 18340 1358 18368 1702
rect 19444 1426 19472 1702
rect 19720 1562 19748 1974
rect 19812 1970 19840 2518
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19996 2106 20024 2450
rect 20272 2106 20300 2746
rect 19984 2100 20036 2106
rect 19984 2042 20036 2048
rect 20260 2100 20312 2106
rect 20260 2042 20312 2048
rect 19800 1964 19852 1970
rect 19800 1906 19852 1912
rect 19870 1660 20178 1669
rect 19870 1658 19876 1660
rect 19932 1658 19956 1660
rect 20012 1658 20036 1660
rect 20092 1658 20116 1660
rect 20172 1658 20178 1660
rect 19932 1606 19934 1658
rect 20114 1606 20116 1658
rect 19870 1604 19876 1606
rect 19932 1604 19956 1606
rect 20012 1604 20036 1606
rect 20092 1604 20116 1606
rect 20172 1604 20178 1606
rect 19870 1595 20178 1604
rect 19708 1556 19760 1562
rect 19708 1498 19760 1504
rect 20272 1494 20300 2042
rect 20640 2038 20668 3334
rect 21928 3058 21956 3470
rect 22112 3398 22140 5120
rect 22468 5102 22520 5108
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 23020 5092 23072 5098
rect 23020 5034 23072 5040
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22112 3194 22140 3334
rect 22204 3194 22232 4014
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22388 3058 22416 5034
rect 23032 4486 23060 5034
rect 23124 4690 23152 5510
rect 23400 5234 23428 5850
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23676 5166 23704 6190
rect 24964 5778 24992 6190
rect 25596 6180 25648 6186
rect 25596 6122 25648 6128
rect 25608 5914 25636 6122
rect 25596 5908 25648 5914
rect 25596 5850 25648 5856
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 26068 5574 26096 6598
rect 26160 6458 26188 6734
rect 26252 6458 26280 6802
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26344 6202 26372 6598
rect 26252 6174 26372 6202
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 26252 5642 26280 6174
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26344 5710 26372 6054
rect 26436 5846 26464 6190
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 26712 5914 26740 6054
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26424 5840 26476 5846
rect 26424 5782 26476 5788
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26240 5636 26292 5642
rect 26240 5578 26292 5584
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4758 23612 4966
rect 23572 4752 23624 4758
rect 23572 4694 23624 4700
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 22664 4146 22692 4422
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 23032 4078 23060 4422
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23676 4010 23704 5102
rect 23952 4078 23980 5510
rect 26252 5234 26280 5578
rect 26344 5234 26372 5646
rect 26896 5234 26924 6820
rect 26976 6802 27028 6808
rect 26984 6556 27292 6565
rect 26984 6554 26990 6556
rect 27046 6554 27070 6556
rect 27126 6554 27150 6556
rect 27206 6554 27230 6556
rect 27286 6554 27292 6556
rect 27046 6502 27048 6554
rect 27228 6502 27230 6554
rect 26984 6500 26990 6502
rect 27046 6500 27070 6502
rect 27126 6500 27150 6502
rect 27206 6500 27230 6502
rect 27286 6500 27292 6502
rect 26984 6491 27292 6500
rect 27252 6384 27304 6390
rect 27252 6326 27304 6332
rect 27264 5556 27292 6326
rect 27356 5846 27384 7278
rect 27528 7268 27580 7274
rect 27528 7210 27580 7216
rect 27540 6730 27568 7210
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 27644 7100 27952 7109
rect 27644 7098 27650 7100
rect 27706 7098 27730 7100
rect 27786 7098 27810 7100
rect 27866 7098 27890 7100
rect 27946 7098 27952 7100
rect 27706 7046 27708 7098
rect 27888 7046 27890 7098
rect 27644 7044 27650 7046
rect 27706 7044 27730 7046
rect 27786 7044 27810 7046
rect 27866 7044 27890 7046
rect 27946 7044 27952 7046
rect 27644 7035 27952 7044
rect 29104 6934 29132 7142
rect 29092 6928 29144 6934
rect 29092 6870 29144 6876
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 28908 6860 28960 6866
rect 28908 6802 28960 6808
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 27528 6724 27580 6730
rect 27528 6666 27580 6672
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27448 6322 27476 6598
rect 27988 6384 28040 6390
rect 27988 6326 28040 6332
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27436 6180 27488 6186
rect 27436 6122 27488 6128
rect 27344 5840 27396 5846
rect 27344 5782 27396 5788
rect 27264 5528 27384 5556
rect 26984 5468 27292 5477
rect 26984 5466 26990 5468
rect 27046 5466 27070 5468
rect 27126 5466 27150 5468
rect 27206 5466 27230 5468
rect 27286 5466 27292 5468
rect 27046 5414 27048 5466
rect 27228 5414 27230 5466
rect 26984 5412 26990 5414
rect 27046 5412 27070 5414
rect 27126 5412 27150 5414
rect 27206 5412 27230 5414
rect 27286 5412 27292 5414
rect 26984 5403 27292 5412
rect 27356 5234 27384 5528
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26332 5228 26384 5234
rect 26332 5170 26384 5176
rect 26608 5228 26660 5234
rect 26608 5170 26660 5176
rect 26884 5228 26936 5234
rect 26884 5170 26936 5176
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 23676 2990 23704 3946
rect 24872 3194 24900 4150
rect 25056 4078 25084 5170
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25424 4826 25452 4966
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 25688 4548 25740 4554
rect 25688 4490 25740 4496
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25332 4282 25360 4422
rect 25320 4276 25372 4282
rect 25320 4218 25372 4224
rect 25700 4146 25728 4490
rect 25792 4282 25820 4558
rect 26620 4282 26648 5170
rect 27448 5166 27476 6122
rect 27540 5710 27568 6258
rect 28000 6254 28028 6326
rect 28092 6254 28120 6802
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 27988 6248 28040 6254
rect 27988 6190 28040 6196
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 27644 6012 27952 6021
rect 27644 6010 27650 6012
rect 27706 6010 27730 6012
rect 27786 6010 27810 6012
rect 27866 6010 27890 6012
rect 27946 6010 27952 6012
rect 27706 5958 27708 6010
rect 27888 5958 27890 6010
rect 27644 5956 27650 5958
rect 27706 5956 27730 5958
rect 27786 5956 27810 5958
rect 27866 5956 27890 5958
rect 27946 5956 27952 5958
rect 27644 5947 27952 5956
rect 28000 5914 28028 6190
rect 28092 6118 28120 6190
rect 28080 6112 28132 6118
rect 28080 6054 28132 6060
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 28092 5778 28120 6054
rect 28080 5772 28132 5778
rect 28080 5714 28132 5720
rect 28368 5710 28396 6666
rect 28920 6662 28948 6802
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 29288 5846 29316 6802
rect 30012 6656 30064 6662
rect 30012 6598 30064 6604
rect 29920 6180 29972 6186
rect 29920 6122 29972 6128
rect 29932 5914 29960 6122
rect 30024 6118 30052 6598
rect 30012 6112 30064 6118
rect 30012 6054 30064 6060
rect 29920 5908 29972 5914
rect 29920 5850 29972 5856
rect 29276 5840 29328 5846
rect 29276 5782 29328 5788
rect 30392 5778 30420 7278
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 30484 5914 30512 6190
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 30380 5772 30432 5778
rect 30380 5714 30432 5720
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 29092 5704 29144 5710
rect 30472 5704 30524 5710
rect 29144 5664 29224 5692
rect 29092 5646 29144 5652
rect 28080 5568 28132 5574
rect 28080 5510 28132 5516
rect 27436 5160 27488 5166
rect 27436 5102 27488 5108
rect 27644 4924 27952 4933
rect 27644 4922 27650 4924
rect 27706 4922 27730 4924
rect 27786 4922 27810 4924
rect 27866 4922 27890 4924
rect 27946 4922 27952 4924
rect 27706 4870 27708 4922
rect 27888 4870 27890 4922
rect 27644 4868 27650 4870
rect 27706 4868 27730 4870
rect 27786 4868 27810 4870
rect 27866 4868 27890 4870
rect 27946 4868 27952 4870
rect 27644 4859 27952 4868
rect 28092 4826 28120 5510
rect 28908 5092 28960 5098
rect 28908 5034 28960 5040
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 28172 4752 28224 4758
rect 28172 4694 28224 4700
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 26984 4380 27292 4389
rect 26984 4378 26990 4380
rect 27046 4378 27070 4380
rect 27126 4378 27150 4380
rect 27206 4378 27230 4380
rect 27286 4378 27292 4380
rect 27046 4326 27048 4378
rect 27228 4326 27230 4378
rect 26984 4324 26990 4326
rect 27046 4324 27070 4326
rect 27126 4324 27150 4326
rect 27206 4324 27230 4326
rect 27286 4324 27292 4326
rect 26984 4315 27292 4324
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 26608 4276 26660 4282
rect 26608 4218 26660 4224
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 25056 3942 25084 4014
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 25056 3058 25084 3878
rect 26620 3398 26648 4218
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 26976 4072 27028 4078
rect 26976 4014 27028 4020
rect 26988 3738 27016 4014
rect 26976 3732 27028 3738
rect 26976 3674 27028 3680
rect 27264 3482 27292 4082
rect 27644 3836 27952 3845
rect 27644 3834 27650 3836
rect 27706 3834 27730 3836
rect 27786 3834 27810 3836
rect 27866 3834 27890 3836
rect 27946 3834 27952 3836
rect 27706 3782 27708 3834
rect 27888 3782 27890 3834
rect 27644 3780 27650 3782
rect 27706 3780 27730 3782
rect 27786 3780 27810 3782
rect 27866 3780 27890 3782
rect 27946 3780 27952 3782
rect 27644 3771 27952 3780
rect 27264 3454 27384 3482
rect 25596 3392 25648 3398
rect 25596 3334 25648 3340
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 25608 3126 25636 3334
rect 26984 3292 27292 3301
rect 26984 3290 26990 3292
rect 27046 3290 27070 3292
rect 27126 3290 27150 3292
rect 27206 3290 27230 3292
rect 27286 3290 27292 3292
rect 27046 3238 27048 3290
rect 27228 3238 27230 3290
rect 26984 3236 26990 3238
rect 27046 3236 27070 3238
rect 27126 3236 27150 3238
rect 27206 3236 27230 3238
rect 27286 3236 27292 3238
rect 26984 3227 27292 3236
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 25596 3120 25648 3126
rect 25596 3062 25648 3068
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 21008 2514 21036 2926
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21652 2514 21680 2790
rect 20996 2508 21048 2514
rect 20996 2450 21048 2456
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 20812 2100 20864 2106
rect 20812 2042 20864 2048
rect 20628 2032 20680 2038
rect 20628 1974 20680 1980
rect 20260 1488 20312 1494
rect 20260 1430 20312 1436
rect 19432 1420 19484 1426
rect 19432 1362 19484 1368
rect 18328 1352 18380 1358
rect 18328 1294 18380 1300
rect 19210 1116 19518 1125
rect 19210 1114 19216 1116
rect 19272 1114 19296 1116
rect 19352 1114 19376 1116
rect 19432 1114 19456 1116
rect 19512 1114 19518 1116
rect 19272 1062 19274 1114
rect 19454 1062 19456 1114
rect 19210 1060 19216 1062
rect 19272 1060 19296 1062
rect 19352 1060 19376 1062
rect 19432 1060 19456 1062
rect 19512 1060 19518 1062
rect 19210 1051 19518 1060
rect 13820 876 13872 882
rect 13820 818 13872 824
rect 20824 814 20852 2042
rect 21008 1902 21036 2450
rect 22020 2446 22048 2926
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 21456 2440 21508 2446
rect 21454 2408 21456 2417
rect 22008 2440 22060 2446
rect 21508 2408 21510 2417
rect 22008 2382 22060 2388
rect 22098 2408 22154 2417
rect 21454 2343 21510 2352
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 20996 1896 21048 1902
rect 20996 1838 21048 1844
rect 21008 1562 21036 1838
rect 21284 1834 21312 2246
rect 21272 1828 21324 1834
rect 21272 1770 21324 1776
rect 20996 1556 21048 1562
rect 20996 1498 21048 1504
rect 21376 1426 21404 2246
rect 22020 2106 22048 2382
rect 22098 2343 22100 2352
rect 22152 2343 22154 2352
rect 22100 2314 22152 2320
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 21456 2032 21508 2038
rect 21456 1974 21508 1980
rect 21468 1834 21496 1974
rect 22008 1896 22060 1902
rect 22112 1884 22140 2314
rect 22204 1902 22232 2790
rect 23676 2650 23704 2926
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22296 2106 22324 2382
rect 22376 2304 22428 2310
rect 22376 2246 22428 2252
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 22060 1856 22140 1884
rect 22192 1896 22244 1902
rect 22008 1838 22060 1844
rect 22192 1838 22244 1844
rect 21456 1828 21508 1834
rect 21456 1770 21508 1776
rect 21732 1828 21784 1834
rect 21732 1770 21784 1776
rect 21744 1562 21772 1770
rect 22204 1562 22232 1838
rect 21732 1556 21784 1562
rect 21732 1498 21784 1504
rect 22192 1556 22244 1562
rect 22192 1498 22244 1504
rect 22296 1494 22324 2042
rect 22284 1488 22336 1494
rect 22284 1430 22336 1436
rect 21364 1420 21416 1426
rect 21364 1362 21416 1368
rect 21548 1420 21600 1426
rect 21548 1362 21600 1368
rect 21560 1018 21588 1362
rect 21548 1012 21600 1018
rect 21548 954 21600 960
rect 22388 814 22416 2246
rect 22664 2106 22692 2450
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 23204 1896 23256 1902
rect 23204 1838 23256 1844
rect 23216 1562 23244 1838
rect 23204 1556 23256 1562
rect 23204 1498 23256 1504
rect 23676 1426 23704 2586
rect 23768 2514 23796 2790
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 23860 2038 23888 2450
rect 24136 2106 24164 2518
rect 25240 2514 25268 2926
rect 25228 2508 25280 2514
rect 25148 2468 25228 2496
rect 24400 2304 24452 2310
rect 24400 2246 24452 2252
rect 24412 2106 24440 2246
rect 24124 2100 24176 2106
rect 24124 2042 24176 2048
rect 24400 2100 24452 2106
rect 24400 2042 24452 2048
rect 23756 2032 23808 2038
rect 23756 1974 23808 1980
rect 23848 2032 23900 2038
rect 23848 1974 23900 1980
rect 23940 2032 23992 2038
rect 23940 1974 23992 1980
rect 23768 1494 23796 1974
rect 23952 1834 23980 1974
rect 24412 1902 24440 2042
rect 25148 1902 25176 2468
rect 25228 2450 25280 2456
rect 25332 2394 25360 2926
rect 26252 2514 26280 2926
rect 26528 2582 26556 2994
rect 26700 2984 26752 2990
rect 26698 2952 26700 2961
rect 26792 2984 26844 2990
rect 26752 2952 26754 2961
rect 26792 2926 26844 2932
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 26698 2887 26754 2896
rect 26700 2848 26752 2854
rect 26700 2790 26752 2796
rect 26516 2576 26568 2582
rect 26516 2518 26568 2524
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 25332 2378 25544 2394
rect 25320 2372 25556 2378
rect 25372 2366 25504 2372
rect 25320 2314 25372 2320
rect 25504 2314 25556 2320
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 25240 1902 25268 2246
rect 25332 2106 25360 2314
rect 25320 2100 25372 2106
rect 25320 2042 25372 2048
rect 25792 1902 25820 2450
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 2106 25912 2246
rect 25872 2100 25924 2106
rect 25872 2042 25924 2048
rect 25884 1902 25912 2042
rect 26148 2032 26200 2038
rect 26148 1974 26200 1980
rect 24400 1896 24452 1902
rect 24400 1838 24452 1844
rect 25136 1896 25188 1902
rect 25136 1838 25188 1844
rect 25228 1896 25280 1902
rect 25228 1838 25280 1844
rect 25780 1896 25832 1902
rect 25780 1838 25832 1844
rect 25872 1896 25924 1902
rect 25872 1838 25924 1844
rect 23940 1828 23992 1834
rect 23940 1770 23992 1776
rect 25148 1562 25176 1838
rect 25596 1828 25648 1834
rect 25596 1770 25648 1776
rect 25412 1760 25464 1766
rect 25412 1702 25464 1708
rect 25136 1556 25188 1562
rect 25136 1498 25188 1504
rect 23756 1488 23808 1494
rect 23756 1430 23808 1436
rect 25424 1426 25452 1702
rect 25608 1562 25636 1770
rect 26160 1766 26188 1974
rect 26148 1760 26200 1766
rect 26148 1702 26200 1708
rect 25596 1556 25648 1562
rect 25596 1498 25648 1504
rect 23664 1420 23716 1426
rect 23664 1362 23716 1368
rect 25412 1420 25464 1426
rect 25412 1362 25464 1368
rect 23676 814 23704 1362
rect 26252 1358 26280 2450
rect 26528 1970 26556 2518
rect 26516 1964 26568 1970
rect 26516 1906 26568 1912
rect 26516 1760 26568 1766
rect 26516 1702 26568 1708
rect 26528 1426 26556 1702
rect 26712 1494 26740 2790
rect 26804 2582 26832 2926
rect 27080 2854 27108 2926
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 26792 2576 26844 2582
rect 26792 2518 26844 2524
rect 26896 2106 26924 2790
rect 27172 2514 27200 3130
rect 27356 2922 27384 3454
rect 27436 3392 27488 3398
rect 27436 3334 27488 3340
rect 27448 3058 27476 3334
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27344 2916 27396 2922
rect 27344 2858 27396 2864
rect 27436 2916 27488 2922
rect 27436 2858 27488 2864
rect 27356 2774 27384 2858
rect 27264 2746 27384 2774
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 27264 2378 27292 2746
rect 27448 2650 27476 2858
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 27344 2508 27396 2514
rect 27344 2450 27396 2456
rect 27252 2372 27304 2378
rect 27252 2314 27304 2320
rect 26984 2204 27292 2213
rect 26984 2202 26990 2204
rect 27046 2202 27070 2204
rect 27126 2202 27150 2204
rect 27206 2202 27230 2204
rect 27286 2202 27292 2204
rect 27046 2150 27048 2202
rect 27228 2150 27230 2202
rect 26984 2148 26990 2150
rect 27046 2148 27070 2150
rect 27126 2148 27150 2150
rect 27206 2148 27230 2150
rect 27286 2148 27292 2150
rect 26984 2139 27292 2148
rect 27356 2106 27384 2450
rect 26884 2100 26936 2106
rect 26884 2042 26936 2048
rect 27344 2100 27396 2106
rect 27344 2042 27396 2048
rect 26700 1488 26752 1494
rect 26700 1430 26752 1436
rect 26896 1426 26924 2042
rect 27068 1896 27120 1902
rect 27068 1838 27120 1844
rect 27080 1562 27108 1838
rect 27068 1556 27120 1562
rect 27068 1498 27120 1504
rect 27448 1426 27476 2586
rect 27540 2378 27568 3062
rect 28000 3058 28028 4558
rect 28092 4214 28120 4626
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 28184 4146 28212 4694
rect 28736 4690 28764 4966
rect 28724 4684 28776 4690
rect 28724 4626 28776 4632
rect 28264 4548 28316 4554
rect 28264 4490 28316 4496
rect 28276 4146 28304 4490
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 28184 3738 28212 4082
rect 28172 3732 28224 3738
rect 28172 3674 28224 3680
rect 28552 3670 28580 4422
rect 28816 3936 28868 3942
rect 28816 3878 28868 3884
rect 28828 3670 28856 3878
rect 28540 3664 28592 3670
rect 28540 3606 28592 3612
rect 28816 3664 28868 3670
rect 28816 3606 28868 3612
rect 28920 3602 28948 5034
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 29012 4826 29040 4966
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29012 3738 29040 4558
rect 29092 4548 29144 4554
rect 29092 4490 29144 4496
rect 29104 4282 29132 4490
rect 29196 4486 29224 5664
rect 30472 5646 30524 5652
rect 29644 5568 29696 5574
rect 29644 5510 29696 5516
rect 29656 5166 29684 5510
rect 30484 5166 30512 5646
rect 30656 5636 30708 5642
rect 30656 5578 30708 5584
rect 30564 5296 30616 5302
rect 30564 5238 30616 5244
rect 29368 5160 29420 5166
rect 29368 5102 29420 5108
rect 29460 5160 29512 5166
rect 29460 5102 29512 5108
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 30472 5160 30524 5166
rect 30472 5102 30524 5108
rect 29380 4826 29408 5102
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 29184 4480 29236 4486
rect 29184 4422 29236 4428
rect 29380 4282 29408 4762
rect 29472 4282 29500 5102
rect 29092 4276 29144 4282
rect 29092 4218 29144 4224
rect 29368 4276 29420 4282
rect 29368 4218 29420 4224
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 29104 3602 29132 4218
rect 29656 3942 29684 5102
rect 30576 4078 30604 5238
rect 30668 5166 30696 5578
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 30564 4072 30616 4078
rect 30564 4014 30616 4020
rect 30932 4072 30984 4078
rect 30932 4014 30984 4020
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 30944 2990 30972 4014
rect 28816 2984 28868 2990
rect 28814 2952 28816 2961
rect 29092 2984 29144 2990
rect 28868 2952 28870 2961
rect 28814 2887 28870 2896
rect 29012 2944 29092 2972
rect 28828 2854 28856 2887
rect 29012 2854 29040 2944
rect 29092 2926 29144 2932
rect 30932 2984 30984 2990
rect 30932 2926 30984 2932
rect 28816 2848 28868 2854
rect 28816 2790 28868 2796
rect 29000 2848 29052 2854
rect 29000 2790 29052 2796
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 29368 2848 29420 2854
rect 29368 2790 29420 2796
rect 27644 2748 27952 2757
rect 27644 2746 27650 2748
rect 27706 2746 27730 2748
rect 27786 2746 27810 2748
rect 27866 2746 27890 2748
rect 27946 2746 27952 2748
rect 27706 2694 27708 2746
rect 27888 2694 27890 2746
rect 27644 2692 27650 2694
rect 27706 2692 27730 2694
rect 27786 2692 27810 2694
rect 27866 2692 27890 2694
rect 27946 2692 27952 2694
rect 27644 2683 27952 2692
rect 29104 2582 29132 2790
rect 29092 2576 29144 2582
rect 29092 2518 29144 2524
rect 29380 2514 29408 2790
rect 29368 2508 29420 2514
rect 29368 2450 29420 2456
rect 27528 2372 27580 2378
rect 27528 2314 27580 2320
rect 28448 1896 28500 1902
rect 28448 1838 28500 1844
rect 27988 1828 28040 1834
rect 27988 1770 28040 1776
rect 27644 1660 27952 1669
rect 27644 1658 27650 1660
rect 27706 1658 27730 1660
rect 27786 1658 27810 1660
rect 27866 1658 27890 1660
rect 27946 1658 27952 1660
rect 27706 1606 27708 1658
rect 27888 1606 27890 1658
rect 27644 1604 27650 1606
rect 27706 1604 27730 1606
rect 27786 1604 27810 1606
rect 27866 1604 27890 1606
rect 27946 1604 27952 1606
rect 27644 1595 27952 1604
rect 26516 1420 26568 1426
rect 26516 1362 26568 1368
rect 26884 1420 26936 1426
rect 26884 1362 26936 1368
rect 27436 1420 27488 1426
rect 27436 1362 27488 1368
rect 26240 1352 26292 1358
rect 26240 1294 26292 1300
rect 25596 1216 25648 1222
rect 25596 1158 25648 1164
rect 25608 814 25636 1158
rect 26252 1018 26280 1294
rect 28000 1290 28028 1770
rect 28460 1562 28488 1838
rect 28448 1556 28500 1562
rect 28448 1498 28500 1504
rect 27988 1284 28040 1290
rect 27988 1226 28040 1232
rect 26984 1116 27292 1125
rect 26984 1114 26990 1116
rect 27046 1114 27070 1116
rect 27126 1114 27150 1116
rect 27206 1114 27230 1116
rect 27286 1114 27292 1116
rect 27046 1062 27048 1114
rect 27228 1062 27230 1114
rect 26984 1060 26990 1062
rect 27046 1060 27070 1062
rect 27126 1060 27150 1062
rect 27206 1060 27230 1062
rect 27286 1060 27292 1062
rect 26984 1051 27292 1060
rect 26240 1012 26292 1018
rect 26240 954 26292 960
rect 9956 808 10008 814
rect 9956 750 10008 756
rect 10692 808 10744 814
rect 10692 750 10744 756
rect 11980 808 12032 814
rect 11980 750 12032 756
rect 20812 808 20864 814
rect 20812 750 20864 756
rect 22376 808 22428 814
rect 22376 750 22428 756
rect 23664 808 23716 814
rect 23664 750 23716 756
rect 25596 808 25648 814
rect 25596 750 25648 756
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 12096 572 12404 581
rect 12096 570 12102 572
rect 12158 570 12182 572
rect 12238 570 12262 572
rect 12318 570 12342 572
rect 12398 570 12404 572
rect 12158 518 12160 570
rect 12340 518 12342 570
rect 12096 516 12102 518
rect 12158 516 12182 518
rect 12238 516 12262 518
rect 12318 516 12342 518
rect 12398 516 12404 518
rect 12096 507 12404 516
rect 19870 572 20178 581
rect 19870 570 19876 572
rect 19932 570 19956 572
rect 20012 570 20036 572
rect 20092 570 20116 572
rect 20172 570 20178 572
rect 19932 518 19934 570
rect 20114 518 20116 570
rect 19870 516 19876 518
rect 19932 516 19956 518
rect 20012 516 20036 518
rect 20092 516 20116 518
rect 20172 516 20178 518
rect 19870 507 20178 516
rect 27644 572 27952 581
rect 27644 570 27650 572
rect 27706 570 27730 572
rect 27786 570 27810 572
rect 27866 570 27890 572
rect 27946 570 27952 572
rect 27706 518 27708 570
rect 27888 518 27890 570
rect 27644 516 27650 518
rect 27706 516 27730 518
rect 27786 516 27810 518
rect 27866 516 27890 518
rect 27946 516 27952 518
rect 27644 507 27952 516
<< via2 >>
rect 11794 21936 11850 21992
rect 12254 21936 12310 21992
rect 23846 21936 23902 21992
rect 24950 21936 25006 21992
rect 25502 21936 25558 21992
rect 26054 21936 26110 21992
rect 27526 21936 27582 21992
rect 28262 21936 28318 21992
rect 8666 21800 8722 21856
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 6458 21684 6514 21720
rect 6458 21664 6460 21684
rect 6460 21664 6512 21684
rect 6512 21664 6514 21684
rect 7286 21684 7342 21720
rect 7286 21664 7288 21684
rect 7288 21664 7340 21684
rect 7340 21664 7342 21684
rect 8390 21684 8446 21720
rect 11442 21786 11498 21788
rect 11522 21786 11578 21788
rect 11602 21786 11658 21788
rect 11682 21786 11738 21788
rect 11442 21734 11488 21786
rect 11488 21734 11498 21786
rect 11522 21734 11552 21786
rect 11552 21734 11564 21786
rect 11564 21734 11578 21786
rect 11602 21734 11616 21786
rect 11616 21734 11628 21786
rect 11628 21734 11658 21786
rect 11682 21734 11692 21786
rect 11692 21734 11738 21786
rect 11442 21732 11498 21734
rect 11522 21732 11578 21734
rect 11602 21732 11658 21734
rect 11682 21732 11738 21734
rect 8390 21664 8392 21684
rect 8392 21664 8444 21684
rect 8444 21664 8446 21684
rect 9954 21684 10010 21720
rect 9954 21664 9956 21684
rect 9956 21664 10008 21684
rect 10008 21664 10010 21684
rect 10322 21684 10378 21720
rect 21638 21800 21694 21856
rect 19216 21786 19272 21788
rect 19296 21786 19352 21788
rect 19376 21786 19432 21788
rect 19456 21786 19512 21788
rect 19216 21734 19262 21786
rect 19262 21734 19272 21786
rect 19296 21734 19326 21786
rect 19326 21734 19338 21786
rect 19338 21734 19352 21786
rect 19376 21734 19390 21786
rect 19390 21734 19402 21786
rect 19402 21734 19432 21786
rect 19456 21734 19466 21786
rect 19466 21734 19512 21786
rect 19216 21732 19272 21734
rect 19296 21732 19352 21734
rect 19376 21732 19432 21734
rect 19456 21732 19512 21734
rect 10322 21664 10324 21684
rect 10324 21664 10376 21684
rect 10376 21664 10378 21684
rect 12806 21684 12862 21720
rect 12806 21664 12808 21684
rect 12808 21664 12860 21684
rect 12860 21664 12862 21684
rect 1950 15000 2006 15056
rect 11702 21528 11758 21584
rect 16670 21528 16726 21584
rect 19430 21528 19486 21584
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 6274 21140 6330 21176
rect 6274 21120 6276 21140
rect 6276 21120 6328 21140
rect 6328 21120 6330 21140
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 3974 18808 4030 18864
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 4250 18808 4306 18864
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 3422 17040 3478 17096
rect 8482 21140 8538 21176
rect 8482 21120 8484 21140
rect 8484 21120 8536 21140
rect 8536 21120 8538 21140
rect 6366 19252 6368 19272
rect 6368 19252 6420 19272
rect 6420 19252 6422 19272
rect 6366 19216 6422 19252
rect 6642 19236 6698 19272
rect 6642 19216 6644 19236
rect 6644 19216 6696 19236
rect 6696 19216 6698 19236
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 3698 15408 3754 15464
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 5262 15408 5318 15464
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 3790 11736 3846 11792
rect 4894 14456 4950 14512
rect 4066 11600 4122 11656
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 3238 9868 3240 9888
rect 3240 9868 3292 9888
rect 3292 9868 3294 9888
rect 3238 9832 3294 9868
rect 3238 9696 3294 9752
rect 3146 9444 3202 9480
rect 3146 9424 3148 9444
rect 3148 9424 3200 9444
rect 3200 9424 3202 9444
rect 3054 7928 3110 7984
rect 2134 6296 2190 6352
rect 2502 6432 2558 6488
rect 2594 6196 2596 6216
rect 2596 6196 2648 6216
rect 2648 6196 2650 6216
rect 2594 6160 2650 6196
rect 3790 9988 3846 10024
rect 3790 9968 3792 9988
rect 3792 9968 3844 9988
rect 3844 9968 3846 9988
rect 4066 9968 4122 10024
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 3606 9560 3662 9616
rect 4066 9632 4122 9688
rect 3974 9424 4030 9480
rect 3698 9036 3754 9072
rect 3698 9016 3700 9036
rect 3700 9016 3752 9036
rect 3752 9016 3754 9036
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 3882 7284 3884 7304
rect 3884 7284 3936 7304
rect 3936 7284 3938 7304
rect 3238 6332 3240 6352
rect 3240 6332 3292 6352
rect 3292 6332 3294 6352
rect 3238 6296 3294 6332
rect 3882 7248 3938 7284
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 3514 6432 3570 6488
rect 4434 11736 4490 11792
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 4434 7384 4490 7440
rect 3422 6196 3424 6216
rect 3424 6196 3476 6216
rect 3476 6196 3478 6216
rect 3422 6160 3478 6196
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 8574 20596 8630 20632
rect 8574 20576 8576 20596
rect 8576 20576 8628 20596
rect 8628 20576 8630 20596
rect 9402 17040 9458 17096
rect 7378 15000 7434 15056
rect 5262 11192 5318 11248
rect 6550 10124 6606 10160
rect 6550 10104 6552 10124
rect 6552 10104 6604 10124
rect 6604 10104 6606 10124
rect 6090 6604 6092 6624
rect 6092 6604 6144 6624
rect 6144 6604 6146 6624
rect 6090 6568 6146 6604
rect 9494 15952 9550 16008
rect 24398 21800 24454 21856
rect 26514 21800 26570 21856
rect 26990 21786 27046 21788
rect 27070 21786 27126 21788
rect 27150 21786 27206 21788
rect 27230 21786 27286 21788
rect 26990 21734 27036 21786
rect 27036 21734 27046 21786
rect 27070 21734 27100 21786
rect 27100 21734 27112 21786
rect 27112 21734 27126 21786
rect 27150 21734 27164 21786
rect 27164 21734 27176 21786
rect 27176 21734 27206 21786
rect 27230 21734 27240 21786
rect 27240 21734 27286 21786
rect 26990 21732 27046 21734
rect 27070 21732 27126 21734
rect 27150 21732 27206 21734
rect 27230 21732 27286 21734
rect 12102 21242 12158 21244
rect 12182 21242 12238 21244
rect 12262 21242 12318 21244
rect 12342 21242 12398 21244
rect 12102 21190 12148 21242
rect 12148 21190 12158 21242
rect 12182 21190 12212 21242
rect 12212 21190 12224 21242
rect 12224 21190 12238 21242
rect 12262 21190 12276 21242
rect 12276 21190 12288 21242
rect 12288 21190 12318 21242
rect 12342 21190 12352 21242
rect 12352 21190 12398 21242
rect 12102 21188 12158 21190
rect 12182 21188 12238 21190
rect 12262 21188 12318 21190
rect 12342 21188 12398 21190
rect 13818 21140 13874 21176
rect 13818 21120 13820 21140
rect 13820 21120 13872 21140
rect 13872 21120 13874 21140
rect 10506 20712 10562 20768
rect 11442 20698 11498 20700
rect 11522 20698 11578 20700
rect 11602 20698 11658 20700
rect 11682 20698 11738 20700
rect 11442 20646 11488 20698
rect 11488 20646 11498 20698
rect 11522 20646 11552 20698
rect 11552 20646 11564 20698
rect 11564 20646 11578 20698
rect 11602 20646 11616 20698
rect 11616 20646 11628 20698
rect 11628 20646 11658 20698
rect 11682 20646 11692 20698
rect 11692 20646 11738 20698
rect 11442 20644 11498 20646
rect 11522 20644 11578 20646
rect 11602 20644 11658 20646
rect 11682 20644 11738 20646
rect 12898 20576 12954 20632
rect 15474 21004 15530 21040
rect 15474 20984 15476 21004
rect 15476 20984 15528 21004
rect 15528 20984 15530 21004
rect 13818 20576 13874 20632
rect 12102 20154 12158 20156
rect 12182 20154 12238 20156
rect 12262 20154 12318 20156
rect 12342 20154 12398 20156
rect 12102 20102 12148 20154
rect 12148 20102 12158 20154
rect 12182 20102 12212 20154
rect 12212 20102 12224 20154
rect 12224 20102 12238 20154
rect 12262 20102 12276 20154
rect 12276 20102 12288 20154
rect 12288 20102 12318 20154
rect 12342 20102 12352 20154
rect 12352 20102 12398 20154
rect 12102 20100 12158 20102
rect 12182 20100 12238 20102
rect 12262 20100 12318 20102
rect 12342 20100 12398 20102
rect 10046 18164 10048 18184
rect 10048 18164 10100 18184
rect 10100 18164 10102 18184
rect 10046 18128 10102 18164
rect 10138 17720 10194 17776
rect 10506 18264 10562 18320
rect 11442 19610 11498 19612
rect 11522 19610 11578 19612
rect 11602 19610 11658 19612
rect 11682 19610 11738 19612
rect 11442 19558 11488 19610
rect 11488 19558 11498 19610
rect 11522 19558 11552 19610
rect 11552 19558 11564 19610
rect 11564 19558 11578 19610
rect 11602 19558 11616 19610
rect 11616 19558 11628 19610
rect 11628 19558 11658 19610
rect 11682 19558 11692 19610
rect 11692 19558 11738 19610
rect 11442 19556 11498 19558
rect 11522 19556 11578 19558
rect 11602 19556 11658 19558
rect 11682 19556 11738 19558
rect 11442 18522 11498 18524
rect 11522 18522 11578 18524
rect 11602 18522 11658 18524
rect 11682 18522 11738 18524
rect 11442 18470 11488 18522
rect 11488 18470 11498 18522
rect 11522 18470 11552 18522
rect 11552 18470 11564 18522
rect 11564 18470 11578 18522
rect 11602 18470 11616 18522
rect 11616 18470 11628 18522
rect 11628 18470 11658 18522
rect 11682 18470 11692 18522
rect 11692 18470 11738 18522
rect 11442 18468 11498 18470
rect 11522 18468 11578 18470
rect 11602 18468 11658 18470
rect 11682 18468 11738 18470
rect 10230 15428 10286 15464
rect 10230 15408 10232 15428
rect 10232 15408 10284 15428
rect 10284 15408 10286 15428
rect 10782 15988 10784 16008
rect 10784 15988 10836 16008
rect 10836 15988 10838 16008
rect 10782 15952 10838 15988
rect 12102 19066 12158 19068
rect 12182 19066 12238 19068
rect 12262 19066 12318 19068
rect 12342 19066 12398 19068
rect 12102 19014 12148 19066
rect 12148 19014 12158 19066
rect 12182 19014 12212 19066
rect 12212 19014 12224 19066
rect 12224 19014 12238 19066
rect 12262 19014 12276 19066
rect 12276 19014 12288 19066
rect 12288 19014 12318 19066
rect 12342 19014 12352 19066
rect 12352 19014 12398 19066
rect 12102 19012 12158 19014
rect 12182 19012 12238 19014
rect 12262 19012 12318 19014
rect 12342 19012 12398 19014
rect 11886 18672 11942 18728
rect 12102 17978 12158 17980
rect 12182 17978 12238 17980
rect 12262 17978 12318 17980
rect 12342 17978 12398 17980
rect 12102 17926 12148 17978
rect 12148 17926 12158 17978
rect 12182 17926 12212 17978
rect 12212 17926 12224 17978
rect 12224 17926 12238 17978
rect 12262 17926 12276 17978
rect 12276 17926 12288 17978
rect 12288 17926 12318 17978
rect 12342 17926 12352 17978
rect 12352 17926 12398 17978
rect 12102 17924 12158 17926
rect 12182 17924 12238 17926
rect 12262 17924 12318 17926
rect 12342 17924 12398 17926
rect 13266 17876 13322 17912
rect 13266 17856 13268 17876
rect 13268 17856 13320 17876
rect 13320 17856 13322 17876
rect 11978 17720 12034 17776
rect 11794 17584 11850 17640
rect 11442 17434 11498 17436
rect 11522 17434 11578 17436
rect 11602 17434 11658 17436
rect 11682 17434 11738 17436
rect 11442 17382 11488 17434
rect 11488 17382 11498 17434
rect 11522 17382 11552 17434
rect 11552 17382 11564 17434
rect 11564 17382 11578 17434
rect 11602 17382 11616 17434
rect 11616 17382 11628 17434
rect 11628 17382 11658 17434
rect 11682 17382 11692 17434
rect 11692 17382 11738 17434
rect 11442 17380 11498 17382
rect 11522 17380 11578 17382
rect 11602 17380 11658 17382
rect 11682 17380 11738 17382
rect 11442 16346 11498 16348
rect 11522 16346 11578 16348
rect 11602 16346 11658 16348
rect 11682 16346 11738 16348
rect 11442 16294 11488 16346
rect 11488 16294 11498 16346
rect 11522 16294 11552 16346
rect 11552 16294 11564 16346
rect 11564 16294 11578 16346
rect 11602 16294 11616 16346
rect 11616 16294 11628 16346
rect 11628 16294 11658 16346
rect 11682 16294 11692 16346
rect 11692 16294 11738 16346
rect 11442 16292 11498 16294
rect 11522 16292 11578 16294
rect 11602 16292 11658 16294
rect 11682 16292 11738 16294
rect 11442 15258 11498 15260
rect 11522 15258 11578 15260
rect 11602 15258 11658 15260
rect 11682 15258 11738 15260
rect 11442 15206 11488 15258
rect 11488 15206 11498 15258
rect 11522 15206 11552 15258
rect 11552 15206 11564 15258
rect 11564 15206 11578 15258
rect 11602 15206 11616 15258
rect 11616 15206 11628 15258
rect 11628 15206 11658 15258
rect 11682 15206 11692 15258
rect 11692 15206 11738 15258
rect 11442 15204 11498 15206
rect 11522 15204 11578 15206
rect 11602 15204 11658 15206
rect 11682 15204 11738 15206
rect 11242 14864 11298 14920
rect 7286 9036 7342 9072
rect 7286 9016 7288 9036
rect 7288 9016 7340 9036
rect 7340 9016 7342 9036
rect 8114 11600 8170 11656
rect 10598 12860 10600 12880
rect 10600 12860 10652 12880
rect 10652 12860 10654 12880
rect 10598 12824 10654 12860
rect 8574 10104 8630 10160
rect 7378 7928 7434 7984
rect 6274 6432 6330 6488
rect 6918 6432 6974 6488
rect 6826 6180 6882 6216
rect 6826 6160 6828 6180
rect 6828 6160 6880 6180
rect 6880 6160 6882 6180
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 7470 6568 7526 6624
rect 10046 11892 10102 11928
rect 10046 11872 10048 11892
rect 10048 11872 10100 11892
rect 10100 11872 10102 11892
rect 8390 7248 8446 7304
rect 11442 14170 11498 14172
rect 11522 14170 11578 14172
rect 11602 14170 11658 14172
rect 11682 14170 11738 14172
rect 11442 14118 11488 14170
rect 11488 14118 11498 14170
rect 11522 14118 11552 14170
rect 11552 14118 11564 14170
rect 11564 14118 11578 14170
rect 11602 14118 11616 14170
rect 11616 14118 11628 14170
rect 11628 14118 11658 14170
rect 11682 14118 11692 14170
rect 11692 14118 11738 14170
rect 11442 14116 11498 14118
rect 11522 14116 11578 14118
rect 11602 14116 11658 14118
rect 11682 14116 11738 14118
rect 12102 16890 12158 16892
rect 12182 16890 12238 16892
rect 12262 16890 12318 16892
rect 12342 16890 12398 16892
rect 12102 16838 12148 16890
rect 12148 16838 12158 16890
rect 12182 16838 12212 16890
rect 12212 16838 12224 16890
rect 12224 16838 12238 16890
rect 12262 16838 12276 16890
rect 12276 16838 12288 16890
rect 12288 16838 12318 16890
rect 12342 16838 12352 16890
rect 12352 16838 12398 16890
rect 12102 16836 12158 16838
rect 12182 16836 12238 16838
rect 12262 16836 12318 16838
rect 12342 16836 12398 16838
rect 12102 15802 12158 15804
rect 12182 15802 12238 15804
rect 12262 15802 12318 15804
rect 12342 15802 12398 15804
rect 12102 15750 12148 15802
rect 12148 15750 12158 15802
rect 12182 15750 12212 15802
rect 12212 15750 12224 15802
rect 12224 15750 12238 15802
rect 12262 15750 12276 15802
rect 12276 15750 12288 15802
rect 12288 15750 12318 15802
rect 12342 15750 12352 15802
rect 12352 15750 12398 15802
rect 12102 15748 12158 15750
rect 12182 15748 12238 15750
rect 12262 15748 12318 15750
rect 12342 15748 12398 15750
rect 12622 14864 12678 14920
rect 12102 14714 12158 14716
rect 12182 14714 12238 14716
rect 12262 14714 12318 14716
rect 12342 14714 12398 14716
rect 12102 14662 12148 14714
rect 12148 14662 12158 14714
rect 12182 14662 12212 14714
rect 12212 14662 12224 14714
rect 12224 14662 12238 14714
rect 12262 14662 12276 14714
rect 12276 14662 12288 14714
rect 12288 14662 12318 14714
rect 12342 14662 12352 14714
rect 12352 14662 12398 14714
rect 12102 14660 12158 14662
rect 12182 14660 12238 14662
rect 12262 14660 12318 14662
rect 12342 14660 12398 14662
rect 11442 13082 11498 13084
rect 11522 13082 11578 13084
rect 11602 13082 11658 13084
rect 11682 13082 11738 13084
rect 11442 13030 11488 13082
rect 11488 13030 11498 13082
rect 11522 13030 11552 13082
rect 11552 13030 11564 13082
rect 11564 13030 11578 13082
rect 11602 13030 11616 13082
rect 11616 13030 11628 13082
rect 11628 13030 11658 13082
rect 11682 13030 11692 13082
rect 11692 13030 11738 13082
rect 11442 13028 11498 13030
rect 11522 13028 11578 13030
rect 11602 13028 11658 13030
rect 11682 13028 11738 13030
rect 11442 11994 11498 11996
rect 11522 11994 11578 11996
rect 11602 11994 11658 11996
rect 11682 11994 11738 11996
rect 11442 11942 11488 11994
rect 11488 11942 11498 11994
rect 11522 11942 11552 11994
rect 11552 11942 11564 11994
rect 11564 11942 11578 11994
rect 11602 11942 11616 11994
rect 11616 11942 11628 11994
rect 11628 11942 11658 11994
rect 11682 11942 11692 11994
rect 11692 11942 11738 11994
rect 11442 11940 11498 11942
rect 11522 11940 11578 11942
rect 11602 11940 11658 11942
rect 11682 11940 11738 11942
rect 11442 10906 11498 10908
rect 11522 10906 11578 10908
rect 11602 10906 11658 10908
rect 11682 10906 11738 10908
rect 11442 10854 11488 10906
rect 11488 10854 11498 10906
rect 11522 10854 11552 10906
rect 11552 10854 11564 10906
rect 11564 10854 11578 10906
rect 11602 10854 11616 10906
rect 11616 10854 11628 10906
rect 11628 10854 11658 10906
rect 11682 10854 11692 10906
rect 11692 10854 11738 10906
rect 11442 10852 11498 10854
rect 11522 10852 11578 10854
rect 11602 10852 11658 10854
rect 11682 10852 11738 10854
rect 13818 17740 13874 17776
rect 13818 17720 13820 17740
rect 13820 17720 13872 17740
rect 13872 17720 13874 17740
rect 14922 18400 14978 18456
rect 15290 18420 15346 18456
rect 15290 18400 15292 18420
rect 15292 18400 15344 18420
rect 15344 18400 15346 18420
rect 12102 13626 12158 13628
rect 12182 13626 12238 13628
rect 12262 13626 12318 13628
rect 12342 13626 12398 13628
rect 12102 13574 12148 13626
rect 12148 13574 12158 13626
rect 12182 13574 12212 13626
rect 12212 13574 12224 13626
rect 12224 13574 12238 13626
rect 12262 13574 12276 13626
rect 12276 13574 12288 13626
rect 12288 13574 12318 13626
rect 12342 13574 12352 13626
rect 12352 13574 12398 13626
rect 12102 13572 12158 13574
rect 12182 13572 12238 13574
rect 12262 13572 12318 13574
rect 12342 13572 12398 13574
rect 12102 12538 12158 12540
rect 12182 12538 12238 12540
rect 12262 12538 12318 12540
rect 12342 12538 12398 12540
rect 12102 12486 12148 12538
rect 12148 12486 12158 12538
rect 12182 12486 12212 12538
rect 12212 12486 12224 12538
rect 12224 12486 12238 12538
rect 12262 12486 12276 12538
rect 12276 12486 12288 12538
rect 12288 12486 12318 12538
rect 12342 12486 12352 12538
rect 12352 12486 12398 12538
rect 12102 12484 12158 12486
rect 12182 12484 12238 12486
rect 12262 12484 12318 12486
rect 12342 12484 12398 12486
rect 11978 11600 12034 11656
rect 12102 11450 12158 11452
rect 12182 11450 12238 11452
rect 12262 11450 12318 11452
rect 12342 11450 12398 11452
rect 12102 11398 12148 11450
rect 12148 11398 12158 11450
rect 12182 11398 12212 11450
rect 12212 11398 12224 11450
rect 12224 11398 12238 11450
rect 12262 11398 12276 11450
rect 12276 11398 12288 11450
rect 12288 11398 12318 11450
rect 12342 11398 12352 11450
rect 12352 11398 12398 11450
rect 12102 11396 12158 11398
rect 12182 11396 12238 11398
rect 12262 11396 12318 11398
rect 12342 11396 12398 11398
rect 13266 14612 13322 14648
rect 13266 14592 13268 14612
rect 13268 14592 13320 14612
rect 13320 14592 13322 14612
rect 14186 15544 14242 15600
rect 15658 19080 15714 19136
rect 15566 17720 15622 17776
rect 16302 19916 16358 19952
rect 16762 20848 16818 20904
rect 16946 20712 17002 20768
rect 16302 19896 16304 19916
rect 16304 19896 16356 19916
rect 16356 19896 16358 19916
rect 16302 18536 16358 18592
rect 16302 17992 16358 18048
rect 11442 9818 11498 9820
rect 11522 9818 11578 9820
rect 11602 9818 11658 9820
rect 11682 9818 11738 9820
rect 11442 9766 11488 9818
rect 11488 9766 11498 9818
rect 11522 9766 11552 9818
rect 11552 9766 11564 9818
rect 11564 9766 11578 9818
rect 11602 9766 11616 9818
rect 11616 9766 11628 9818
rect 11628 9766 11658 9818
rect 11682 9766 11692 9818
rect 11692 9766 11738 9818
rect 11442 9764 11498 9766
rect 11522 9764 11578 9766
rect 11602 9764 11658 9766
rect 11682 9764 11738 9766
rect 9862 7948 9918 7984
rect 9862 7928 9864 7948
rect 9864 7928 9916 7948
rect 9916 7928 9918 7948
rect 10138 7928 10194 7984
rect 10598 7928 10654 7984
rect 10322 7792 10378 7848
rect 6182 3596 6238 3632
rect 6182 3576 6184 3596
rect 6184 3576 6236 3596
rect 6236 3576 6238 3596
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 8666 3612 8668 3632
rect 8668 3612 8720 3632
rect 8720 3612 8722 3632
rect 8666 3576 8722 3612
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 11442 8730 11498 8732
rect 11522 8730 11578 8732
rect 11602 8730 11658 8732
rect 11682 8730 11738 8732
rect 11442 8678 11488 8730
rect 11488 8678 11498 8730
rect 11522 8678 11552 8730
rect 11552 8678 11564 8730
rect 11564 8678 11578 8730
rect 11602 8678 11616 8730
rect 11616 8678 11628 8730
rect 11628 8678 11658 8730
rect 11682 8678 11692 8730
rect 11692 8678 11738 8730
rect 11442 8676 11498 8678
rect 11522 8676 11578 8678
rect 11602 8676 11658 8678
rect 11682 8676 11738 8678
rect 11442 7642 11498 7644
rect 11522 7642 11578 7644
rect 11602 7642 11658 7644
rect 11682 7642 11738 7644
rect 11442 7590 11488 7642
rect 11488 7590 11498 7642
rect 11522 7590 11552 7642
rect 11552 7590 11564 7642
rect 11564 7590 11578 7642
rect 11602 7590 11616 7642
rect 11616 7590 11628 7642
rect 11628 7590 11658 7642
rect 11682 7590 11692 7642
rect 11692 7590 11738 7642
rect 11442 7588 11498 7590
rect 11522 7588 11578 7590
rect 11602 7588 11658 7590
rect 11682 7588 11738 7590
rect 12102 10362 12158 10364
rect 12182 10362 12238 10364
rect 12262 10362 12318 10364
rect 12342 10362 12398 10364
rect 12102 10310 12148 10362
rect 12148 10310 12158 10362
rect 12182 10310 12212 10362
rect 12212 10310 12224 10362
rect 12224 10310 12238 10362
rect 12262 10310 12276 10362
rect 12276 10310 12288 10362
rect 12288 10310 12318 10362
rect 12342 10310 12352 10362
rect 12352 10310 12398 10362
rect 12102 10308 12158 10310
rect 12182 10308 12238 10310
rect 12262 10308 12318 10310
rect 12342 10308 12398 10310
rect 12070 10140 12072 10160
rect 12072 10140 12124 10160
rect 12124 10140 12126 10160
rect 12070 10104 12126 10140
rect 12346 9968 12402 10024
rect 12102 9274 12158 9276
rect 12182 9274 12238 9276
rect 12262 9274 12318 9276
rect 12342 9274 12398 9276
rect 12102 9222 12148 9274
rect 12148 9222 12158 9274
rect 12182 9222 12212 9274
rect 12212 9222 12224 9274
rect 12224 9222 12238 9274
rect 12262 9222 12276 9274
rect 12276 9222 12288 9274
rect 12288 9222 12318 9274
rect 12342 9222 12352 9274
rect 12352 9222 12398 9274
rect 12102 9220 12158 9222
rect 12182 9220 12238 9222
rect 12262 9220 12318 9222
rect 12342 9220 12398 9222
rect 11886 9052 11888 9072
rect 11888 9052 11940 9072
rect 11940 9052 11942 9072
rect 11886 9016 11942 9052
rect 14094 11328 14150 11384
rect 12806 9016 12862 9072
rect 12102 8186 12158 8188
rect 12182 8186 12238 8188
rect 12262 8186 12318 8188
rect 12342 8186 12398 8188
rect 12102 8134 12148 8186
rect 12148 8134 12158 8186
rect 12182 8134 12212 8186
rect 12212 8134 12224 8186
rect 12224 8134 12238 8186
rect 12262 8134 12276 8186
rect 12276 8134 12288 8186
rect 12288 8134 12318 8186
rect 12342 8134 12352 8186
rect 12352 8134 12398 8186
rect 12102 8132 12158 8134
rect 12182 8132 12238 8134
rect 12262 8132 12318 8134
rect 12342 8132 12398 8134
rect 10966 5752 11022 5808
rect 11794 7284 11796 7304
rect 11796 7284 11848 7304
rect 11848 7284 11850 7304
rect 11794 7248 11850 7284
rect 12102 7098 12158 7100
rect 12182 7098 12238 7100
rect 12262 7098 12318 7100
rect 12342 7098 12398 7100
rect 12102 7046 12148 7098
rect 12148 7046 12158 7098
rect 12182 7046 12212 7098
rect 12212 7046 12224 7098
rect 12224 7046 12238 7098
rect 12262 7046 12276 7098
rect 12276 7046 12288 7098
rect 12288 7046 12318 7098
rect 12342 7046 12352 7098
rect 12352 7046 12398 7098
rect 12102 7044 12158 7046
rect 12182 7044 12238 7046
rect 12262 7044 12318 7046
rect 12342 7044 12398 7046
rect 11442 6554 11498 6556
rect 11522 6554 11578 6556
rect 11602 6554 11658 6556
rect 11682 6554 11738 6556
rect 11442 6502 11488 6554
rect 11488 6502 11498 6554
rect 11522 6502 11552 6554
rect 11552 6502 11564 6554
rect 11564 6502 11578 6554
rect 11602 6502 11616 6554
rect 11616 6502 11628 6554
rect 11628 6502 11658 6554
rect 11682 6502 11692 6554
rect 11692 6502 11738 6554
rect 11442 6500 11498 6502
rect 11522 6500 11578 6502
rect 11602 6500 11658 6502
rect 11682 6500 11738 6502
rect 11442 5466 11498 5468
rect 11522 5466 11578 5468
rect 11602 5466 11658 5468
rect 11682 5466 11738 5468
rect 11442 5414 11488 5466
rect 11488 5414 11498 5466
rect 11522 5414 11552 5466
rect 11552 5414 11564 5466
rect 11564 5414 11578 5466
rect 11602 5414 11616 5466
rect 11616 5414 11628 5466
rect 11628 5414 11658 5466
rect 11682 5414 11692 5466
rect 11692 5414 11738 5466
rect 11442 5412 11498 5414
rect 11522 5412 11578 5414
rect 11602 5412 11658 5414
rect 11682 5412 11738 5414
rect 11442 4378 11498 4380
rect 11522 4378 11578 4380
rect 11602 4378 11658 4380
rect 11682 4378 11738 4380
rect 11442 4326 11488 4378
rect 11488 4326 11498 4378
rect 11522 4326 11552 4378
rect 11552 4326 11564 4378
rect 11564 4326 11578 4378
rect 11602 4326 11616 4378
rect 11616 4326 11628 4378
rect 11628 4326 11658 4378
rect 11682 4326 11692 4378
rect 11692 4326 11738 4378
rect 11442 4324 11498 4326
rect 11522 4324 11578 4326
rect 11602 4324 11658 4326
rect 11682 4324 11738 4326
rect 10690 2760 10746 2816
rect 11442 3290 11498 3292
rect 11522 3290 11578 3292
rect 11602 3290 11658 3292
rect 11682 3290 11738 3292
rect 11442 3238 11488 3290
rect 11488 3238 11498 3290
rect 11522 3238 11552 3290
rect 11552 3238 11564 3290
rect 11564 3238 11578 3290
rect 11602 3238 11616 3290
rect 11616 3238 11628 3290
rect 11628 3238 11658 3290
rect 11682 3238 11692 3290
rect 11692 3238 11738 3290
rect 11442 3236 11498 3238
rect 11522 3236 11578 3238
rect 11602 3236 11658 3238
rect 11682 3236 11738 3238
rect 11518 2796 11520 2816
rect 11520 2796 11572 2816
rect 11572 2796 11574 2816
rect 11518 2760 11574 2796
rect 11702 2388 11704 2408
rect 11704 2388 11756 2408
rect 11756 2388 11758 2408
rect 11702 2352 11758 2388
rect 11442 2202 11498 2204
rect 11522 2202 11578 2204
rect 11602 2202 11658 2204
rect 11682 2202 11738 2204
rect 11442 2150 11488 2202
rect 11488 2150 11498 2202
rect 11522 2150 11552 2202
rect 11552 2150 11564 2202
rect 11564 2150 11578 2202
rect 11602 2150 11616 2202
rect 11616 2150 11628 2202
rect 11628 2150 11658 2202
rect 11682 2150 11692 2202
rect 11692 2150 11738 2202
rect 11442 2148 11498 2150
rect 11522 2148 11578 2150
rect 11602 2148 11658 2150
rect 11682 2148 11738 2150
rect 13082 7112 13138 7168
rect 13082 6160 13138 6216
rect 12102 6010 12158 6012
rect 12182 6010 12238 6012
rect 12262 6010 12318 6012
rect 12342 6010 12398 6012
rect 12102 5958 12148 6010
rect 12148 5958 12158 6010
rect 12182 5958 12212 6010
rect 12212 5958 12224 6010
rect 12224 5958 12238 6010
rect 12262 5958 12276 6010
rect 12276 5958 12288 6010
rect 12288 5958 12318 6010
rect 12342 5958 12352 6010
rect 12352 5958 12398 6010
rect 12102 5956 12158 5958
rect 12182 5956 12238 5958
rect 12262 5956 12318 5958
rect 12342 5956 12398 5958
rect 12162 5772 12218 5808
rect 12162 5752 12164 5772
rect 12164 5752 12216 5772
rect 12216 5752 12218 5772
rect 12898 5616 12954 5672
rect 12102 4922 12158 4924
rect 12182 4922 12238 4924
rect 12262 4922 12318 4924
rect 12342 4922 12398 4924
rect 12102 4870 12148 4922
rect 12148 4870 12158 4922
rect 12182 4870 12212 4922
rect 12212 4870 12224 4922
rect 12224 4870 12238 4922
rect 12262 4870 12276 4922
rect 12276 4870 12288 4922
rect 12288 4870 12318 4922
rect 12342 4870 12352 4922
rect 12352 4870 12398 4922
rect 12102 4868 12158 4870
rect 12182 4868 12238 4870
rect 12262 4868 12318 4870
rect 12342 4868 12398 4870
rect 12102 3834 12158 3836
rect 12182 3834 12238 3836
rect 12262 3834 12318 3836
rect 12342 3834 12398 3836
rect 12102 3782 12148 3834
rect 12148 3782 12158 3834
rect 12182 3782 12212 3834
rect 12212 3782 12224 3834
rect 12224 3782 12238 3834
rect 12262 3782 12276 3834
rect 12276 3782 12288 3834
rect 12288 3782 12318 3834
rect 12342 3782 12352 3834
rect 12352 3782 12398 3834
rect 12102 3780 12158 3782
rect 12182 3780 12238 3782
rect 12262 3780 12318 3782
rect 12342 3780 12398 3782
rect 17682 20712 17738 20768
rect 17590 19932 17592 19952
rect 17592 19932 17644 19952
rect 17644 19932 17646 19952
rect 17590 19896 17646 19932
rect 16670 19080 16726 19136
rect 16946 19236 17002 19272
rect 17130 19252 17132 19272
rect 17132 19252 17184 19272
rect 17184 19252 17186 19272
rect 16946 19216 16948 19236
rect 16948 19216 17000 19236
rect 17000 19216 17002 19236
rect 17130 19216 17186 19252
rect 17038 19080 17094 19136
rect 17038 18944 17094 19000
rect 16946 18828 17002 18864
rect 16946 18808 16948 18828
rect 16948 18808 17000 18828
rect 17000 18808 17002 18828
rect 16670 17332 16726 17368
rect 16670 17312 16672 17332
rect 16672 17312 16724 17332
rect 16724 17312 16726 17332
rect 18234 20848 18290 20904
rect 19246 21412 19302 21448
rect 19246 21392 19248 21412
rect 19248 21392 19300 21412
rect 19300 21392 19302 21412
rect 18050 20476 18052 20496
rect 18052 20476 18104 20496
rect 18104 20476 18106 20496
rect 18050 20440 18106 20476
rect 18326 20340 18328 20360
rect 18328 20340 18380 20360
rect 18380 20340 18382 20360
rect 17222 18400 17278 18456
rect 17498 18536 17554 18592
rect 17498 18400 17554 18456
rect 17038 17856 17094 17912
rect 17130 17720 17186 17776
rect 16210 14476 16266 14512
rect 16210 14456 16212 14476
rect 16212 14456 16264 14476
rect 16264 14456 16266 14476
rect 15934 12824 15990 12880
rect 16302 12824 16358 12880
rect 16486 12824 16542 12880
rect 16302 10104 16358 10160
rect 16026 9968 16082 10024
rect 15566 9036 15622 9072
rect 15566 9016 15568 9036
rect 15568 9016 15620 9036
rect 15620 9016 15622 9036
rect 14922 7520 14978 7576
rect 14002 5772 14058 5808
rect 14002 5752 14004 5772
rect 14004 5752 14056 5772
rect 14056 5752 14058 5772
rect 14186 5752 14242 5808
rect 13542 5616 13598 5672
rect 13818 5208 13874 5264
rect 15014 7384 15070 7440
rect 15566 7792 15622 7848
rect 15658 7148 15660 7168
rect 15660 7148 15712 7168
rect 15712 7148 15714 7168
rect 15658 7112 15714 7148
rect 14738 5616 14794 5672
rect 15750 5752 15806 5808
rect 15198 5616 15254 5672
rect 11886 2760 11942 2816
rect 12102 2746 12158 2748
rect 12182 2746 12238 2748
rect 12262 2746 12318 2748
rect 12342 2746 12398 2748
rect 12102 2694 12148 2746
rect 12148 2694 12158 2746
rect 12182 2694 12212 2746
rect 12212 2694 12224 2746
rect 12224 2694 12238 2746
rect 12262 2694 12276 2746
rect 12276 2694 12288 2746
rect 12288 2694 12318 2746
rect 12342 2694 12352 2746
rect 12352 2694 12398 2746
rect 12102 2692 12158 2694
rect 12182 2692 12238 2694
rect 12262 2692 12318 2694
rect 12342 2692 12398 2694
rect 12102 1658 12158 1660
rect 12182 1658 12238 1660
rect 12262 1658 12318 1660
rect 12342 1658 12398 1660
rect 12102 1606 12148 1658
rect 12148 1606 12158 1658
rect 12182 1606 12212 1658
rect 12212 1606 12224 1658
rect 12224 1606 12238 1658
rect 12262 1606 12276 1658
rect 12276 1606 12288 1658
rect 12288 1606 12318 1658
rect 12342 1606 12352 1658
rect 12352 1606 12398 1658
rect 12102 1604 12158 1606
rect 12182 1604 12238 1606
rect 12262 1604 12318 1606
rect 12342 1604 12398 1606
rect 11442 1114 11498 1116
rect 11522 1114 11578 1116
rect 11602 1114 11658 1116
rect 11682 1114 11738 1116
rect 11442 1062 11488 1114
rect 11488 1062 11498 1114
rect 11522 1062 11552 1114
rect 11552 1062 11564 1114
rect 11564 1062 11578 1114
rect 11602 1062 11616 1114
rect 11616 1062 11628 1114
rect 11628 1062 11658 1114
rect 11682 1062 11692 1114
rect 11692 1062 11738 1114
rect 11442 1060 11498 1062
rect 11522 1060 11578 1062
rect 11602 1060 11658 1062
rect 11682 1060 11738 1062
rect 16302 7520 16358 7576
rect 16578 7248 16634 7304
rect 16118 5208 16174 5264
rect 17590 15000 17646 15056
rect 17866 16632 17922 16688
rect 18326 20304 18382 20340
rect 18878 20304 18934 20360
rect 19216 20698 19272 20700
rect 19296 20698 19352 20700
rect 19376 20698 19432 20700
rect 19456 20698 19512 20700
rect 19216 20646 19262 20698
rect 19262 20646 19272 20698
rect 19296 20646 19326 20698
rect 19326 20646 19338 20698
rect 19338 20646 19352 20698
rect 19376 20646 19390 20698
rect 19390 20646 19402 20698
rect 19402 20646 19432 20698
rect 19456 20646 19466 20698
rect 19466 20646 19512 20698
rect 19216 20644 19272 20646
rect 19296 20644 19352 20646
rect 19376 20644 19432 20646
rect 19456 20644 19512 20646
rect 19062 20440 19118 20496
rect 19876 21242 19932 21244
rect 19956 21242 20012 21244
rect 20036 21242 20092 21244
rect 20116 21242 20172 21244
rect 19876 21190 19922 21242
rect 19922 21190 19932 21242
rect 19956 21190 19986 21242
rect 19986 21190 19998 21242
rect 19998 21190 20012 21242
rect 20036 21190 20050 21242
rect 20050 21190 20062 21242
rect 20062 21190 20092 21242
rect 20116 21190 20126 21242
rect 20126 21190 20172 21242
rect 19876 21188 19932 21190
rect 19956 21188 20012 21190
rect 20036 21188 20092 21190
rect 20116 21188 20172 21190
rect 18510 19760 18566 19816
rect 19062 19780 19118 19816
rect 19062 19760 19064 19780
rect 19064 19760 19116 19780
rect 19116 19760 19118 19780
rect 19216 19610 19272 19612
rect 19296 19610 19352 19612
rect 19376 19610 19432 19612
rect 19456 19610 19512 19612
rect 19216 19558 19262 19610
rect 19262 19558 19272 19610
rect 19296 19558 19326 19610
rect 19326 19558 19338 19610
rect 19338 19558 19352 19610
rect 19376 19558 19390 19610
rect 19390 19558 19402 19610
rect 19402 19558 19432 19610
rect 19456 19558 19466 19610
rect 19466 19558 19512 19610
rect 19216 19556 19272 19558
rect 19296 19556 19352 19558
rect 19376 19556 19432 19558
rect 19456 19556 19512 19558
rect 19876 20154 19932 20156
rect 19956 20154 20012 20156
rect 20036 20154 20092 20156
rect 20116 20154 20172 20156
rect 19876 20102 19922 20154
rect 19922 20102 19932 20154
rect 19956 20102 19986 20154
rect 19986 20102 19998 20154
rect 19998 20102 20012 20154
rect 20036 20102 20050 20154
rect 20050 20102 20062 20154
rect 20062 20102 20092 20154
rect 20116 20102 20126 20154
rect 20126 20102 20172 20154
rect 19876 20100 19932 20102
rect 19956 20100 20012 20102
rect 20036 20100 20092 20102
rect 20116 20100 20172 20102
rect 20350 20052 20406 20088
rect 20350 20032 20352 20052
rect 20352 20032 20404 20052
rect 20404 20032 20406 20052
rect 19154 19252 19156 19272
rect 19156 19252 19208 19272
rect 19208 19252 19210 19272
rect 18510 18944 18566 19000
rect 18234 17992 18290 18048
rect 19154 19216 19210 19252
rect 19216 18522 19272 18524
rect 19296 18522 19352 18524
rect 19376 18522 19432 18524
rect 19456 18522 19512 18524
rect 19216 18470 19262 18522
rect 19262 18470 19272 18522
rect 19296 18470 19326 18522
rect 19326 18470 19338 18522
rect 19338 18470 19352 18522
rect 19376 18470 19390 18522
rect 19390 18470 19402 18522
rect 19402 18470 19432 18522
rect 19456 18470 19466 18522
rect 19466 18470 19512 18522
rect 19216 18468 19272 18470
rect 19296 18468 19352 18470
rect 19376 18468 19432 18470
rect 19456 18468 19512 18470
rect 18050 14592 18106 14648
rect 19216 17434 19272 17436
rect 19296 17434 19352 17436
rect 19376 17434 19432 17436
rect 19456 17434 19512 17436
rect 19216 17382 19262 17434
rect 19262 17382 19272 17434
rect 19296 17382 19326 17434
rect 19326 17382 19338 17434
rect 19338 17382 19352 17434
rect 19376 17382 19390 17434
rect 19390 17382 19402 17434
rect 19402 17382 19432 17434
rect 19456 17382 19466 17434
rect 19466 17382 19512 17434
rect 19216 17380 19272 17382
rect 19296 17380 19352 17382
rect 19376 17380 19432 17382
rect 19456 17380 19512 17382
rect 19216 16346 19272 16348
rect 19296 16346 19352 16348
rect 19376 16346 19432 16348
rect 19456 16346 19512 16348
rect 19216 16294 19262 16346
rect 19262 16294 19272 16346
rect 19296 16294 19326 16346
rect 19326 16294 19338 16346
rect 19338 16294 19352 16346
rect 19376 16294 19390 16346
rect 19390 16294 19402 16346
rect 19402 16294 19432 16346
rect 19456 16294 19466 16346
rect 19466 16294 19512 16346
rect 19216 16292 19272 16294
rect 19296 16292 19352 16294
rect 19376 16292 19432 16294
rect 19456 16292 19512 16294
rect 20258 19080 20314 19136
rect 19876 19066 19932 19068
rect 19956 19066 20012 19068
rect 20036 19066 20092 19068
rect 20116 19066 20172 19068
rect 19876 19014 19922 19066
rect 19922 19014 19932 19066
rect 19956 19014 19986 19066
rect 19986 19014 19998 19066
rect 19998 19014 20012 19066
rect 20036 19014 20050 19066
rect 20050 19014 20062 19066
rect 20062 19014 20092 19066
rect 20116 19014 20126 19066
rect 20126 19014 20172 19066
rect 19876 19012 19932 19014
rect 19956 19012 20012 19014
rect 20036 19012 20092 19014
rect 20116 19012 20172 19014
rect 20258 18536 20314 18592
rect 20074 18400 20130 18456
rect 20718 18536 20774 18592
rect 20442 17992 20498 18048
rect 19876 17978 19932 17980
rect 19956 17978 20012 17980
rect 20036 17978 20092 17980
rect 20116 17978 20172 17980
rect 19876 17926 19922 17978
rect 19922 17926 19932 17978
rect 19956 17926 19986 17978
rect 19986 17926 19998 17978
rect 19998 17926 20012 17978
rect 20036 17926 20050 17978
rect 20050 17926 20062 17978
rect 20062 17926 20092 17978
rect 20116 17926 20126 17978
rect 20126 17926 20172 17978
rect 19876 17924 19932 17926
rect 19956 17924 20012 17926
rect 20036 17924 20092 17926
rect 20116 17924 20172 17926
rect 19876 16890 19932 16892
rect 19956 16890 20012 16892
rect 20036 16890 20092 16892
rect 20116 16890 20172 16892
rect 19876 16838 19922 16890
rect 19922 16838 19932 16890
rect 19956 16838 19986 16890
rect 19986 16838 19998 16890
rect 19998 16838 20012 16890
rect 20036 16838 20050 16890
rect 20050 16838 20062 16890
rect 20062 16838 20092 16890
rect 20116 16838 20126 16890
rect 20126 16838 20172 16890
rect 19876 16836 19932 16838
rect 19956 16836 20012 16838
rect 20036 16836 20092 16838
rect 20116 16836 20172 16838
rect 20442 16768 20498 16824
rect 20166 16632 20222 16688
rect 20442 16632 20498 16688
rect 19216 15258 19272 15260
rect 19296 15258 19352 15260
rect 19376 15258 19432 15260
rect 19456 15258 19512 15260
rect 19216 15206 19262 15258
rect 19262 15206 19272 15258
rect 19296 15206 19326 15258
rect 19326 15206 19338 15258
rect 19338 15206 19352 15258
rect 19376 15206 19390 15258
rect 19390 15206 19402 15258
rect 19402 15206 19432 15258
rect 19456 15206 19466 15258
rect 19466 15206 19512 15258
rect 19216 15204 19272 15206
rect 19296 15204 19352 15206
rect 19376 15204 19432 15206
rect 19456 15204 19512 15206
rect 17682 11328 17738 11384
rect 17774 11192 17830 11248
rect 19216 14170 19272 14172
rect 19296 14170 19352 14172
rect 19376 14170 19432 14172
rect 19456 14170 19512 14172
rect 19216 14118 19262 14170
rect 19262 14118 19272 14170
rect 19296 14118 19326 14170
rect 19326 14118 19338 14170
rect 19338 14118 19352 14170
rect 19376 14118 19390 14170
rect 19390 14118 19402 14170
rect 19402 14118 19432 14170
rect 19456 14118 19466 14170
rect 19466 14118 19512 14170
rect 19216 14116 19272 14118
rect 19296 14116 19352 14118
rect 19376 14116 19432 14118
rect 19456 14116 19512 14118
rect 20258 15816 20314 15872
rect 19876 15802 19932 15804
rect 19956 15802 20012 15804
rect 20036 15802 20092 15804
rect 20116 15802 20172 15804
rect 19876 15750 19922 15802
rect 19922 15750 19932 15802
rect 19956 15750 19986 15802
rect 19986 15750 19998 15802
rect 19998 15750 20012 15802
rect 20036 15750 20050 15802
rect 20050 15750 20062 15802
rect 20062 15750 20092 15802
rect 20116 15750 20126 15802
rect 20126 15750 20172 15802
rect 19876 15748 19932 15750
rect 19956 15748 20012 15750
rect 20036 15748 20092 15750
rect 20116 15748 20172 15750
rect 19876 14714 19932 14716
rect 19956 14714 20012 14716
rect 20036 14714 20092 14716
rect 20116 14714 20172 14716
rect 19876 14662 19922 14714
rect 19922 14662 19932 14714
rect 19956 14662 19986 14714
rect 19986 14662 19998 14714
rect 19998 14662 20012 14714
rect 20036 14662 20050 14714
rect 20050 14662 20062 14714
rect 20062 14662 20092 14714
rect 20116 14662 20126 14714
rect 20126 14662 20172 14714
rect 19876 14660 19932 14662
rect 19956 14660 20012 14662
rect 20036 14660 20092 14662
rect 20116 14660 20172 14662
rect 19890 14184 19946 14240
rect 19876 13626 19932 13628
rect 19956 13626 20012 13628
rect 20036 13626 20092 13628
rect 20116 13626 20172 13628
rect 19876 13574 19922 13626
rect 19922 13574 19932 13626
rect 19956 13574 19986 13626
rect 19986 13574 19998 13626
rect 19998 13574 20012 13626
rect 20036 13574 20050 13626
rect 20050 13574 20062 13626
rect 20062 13574 20092 13626
rect 20116 13574 20126 13626
rect 20126 13574 20172 13626
rect 19876 13572 19932 13574
rect 19956 13572 20012 13574
rect 20036 13572 20092 13574
rect 20116 13572 20172 13574
rect 19982 13368 20038 13424
rect 19216 13082 19272 13084
rect 19296 13082 19352 13084
rect 19376 13082 19432 13084
rect 19456 13082 19512 13084
rect 19216 13030 19262 13082
rect 19262 13030 19272 13082
rect 19296 13030 19326 13082
rect 19326 13030 19338 13082
rect 19338 13030 19352 13082
rect 19376 13030 19390 13082
rect 19390 13030 19402 13082
rect 19402 13030 19432 13082
rect 19456 13030 19466 13082
rect 19466 13030 19512 13082
rect 19216 13028 19272 13030
rect 19296 13028 19352 13030
rect 19376 13028 19432 13030
rect 19456 13028 19512 13030
rect 20718 16768 20774 16824
rect 20626 16632 20682 16688
rect 22926 20848 22982 20904
rect 22098 19760 22154 19816
rect 21454 18808 21510 18864
rect 20810 15988 20812 16008
rect 20812 15988 20864 16008
rect 20864 15988 20866 16008
rect 20810 15952 20866 15988
rect 20810 15680 20866 15736
rect 19876 12538 19932 12540
rect 19956 12538 20012 12540
rect 20036 12538 20092 12540
rect 20116 12538 20172 12540
rect 19876 12486 19922 12538
rect 19922 12486 19932 12538
rect 19956 12486 19986 12538
rect 19986 12486 19998 12538
rect 19998 12486 20012 12538
rect 20036 12486 20050 12538
rect 20050 12486 20062 12538
rect 20062 12486 20092 12538
rect 20116 12486 20126 12538
rect 20126 12486 20172 12538
rect 19876 12484 19932 12486
rect 19956 12484 20012 12486
rect 20036 12484 20092 12486
rect 20116 12484 20172 12486
rect 21086 15408 21142 15464
rect 20902 15000 20958 15056
rect 21270 17604 21326 17640
rect 21270 17584 21272 17604
rect 21272 17584 21324 17604
rect 21324 17584 21326 17604
rect 22282 19624 22338 19680
rect 22742 19796 22744 19816
rect 22744 19796 22796 19816
rect 22796 19796 22798 19816
rect 22742 19760 22798 19796
rect 23110 20032 23166 20088
rect 22926 19624 22982 19680
rect 23018 19116 23020 19136
rect 23020 19116 23072 19136
rect 23072 19116 23074 19136
rect 23018 19080 23074 19116
rect 22926 18400 22982 18456
rect 22466 18264 22522 18320
rect 21914 18128 21970 18184
rect 22466 17992 22522 18048
rect 21178 14864 21234 14920
rect 15014 2352 15070 2408
rect 19216 11994 19272 11996
rect 19296 11994 19352 11996
rect 19376 11994 19432 11996
rect 19456 11994 19512 11996
rect 19216 11942 19262 11994
rect 19262 11942 19272 11994
rect 19296 11942 19326 11994
rect 19326 11942 19338 11994
rect 19338 11942 19352 11994
rect 19376 11942 19390 11994
rect 19390 11942 19402 11994
rect 19402 11942 19432 11994
rect 19456 11942 19466 11994
rect 19466 11942 19512 11994
rect 19216 11940 19272 11942
rect 19296 11940 19352 11942
rect 19376 11940 19432 11942
rect 19456 11940 19512 11942
rect 19876 11450 19932 11452
rect 19956 11450 20012 11452
rect 20036 11450 20092 11452
rect 20116 11450 20172 11452
rect 19876 11398 19922 11450
rect 19922 11398 19932 11450
rect 19956 11398 19986 11450
rect 19986 11398 19998 11450
rect 19998 11398 20012 11450
rect 20036 11398 20050 11450
rect 20050 11398 20062 11450
rect 20062 11398 20092 11450
rect 20116 11398 20126 11450
rect 20126 11398 20172 11450
rect 19876 11396 19932 11398
rect 19956 11396 20012 11398
rect 20036 11396 20092 11398
rect 20116 11396 20172 11398
rect 19216 10906 19272 10908
rect 19296 10906 19352 10908
rect 19376 10906 19432 10908
rect 19456 10906 19512 10908
rect 19216 10854 19262 10906
rect 19262 10854 19272 10906
rect 19296 10854 19326 10906
rect 19326 10854 19338 10906
rect 19338 10854 19352 10906
rect 19376 10854 19390 10906
rect 19390 10854 19402 10906
rect 19402 10854 19432 10906
rect 19456 10854 19466 10906
rect 19466 10854 19512 10906
rect 19216 10852 19272 10854
rect 19296 10852 19352 10854
rect 19376 10852 19432 10854
rect 19456 10852 19512 10854
rect 19216 9818 19272 9820
rect 19296 9818 19352 9820
rect 19376 9818 19432 9820
rect 19456 9818 19512 9820
rect 19216 9766 19262 9818
rect 19262 9766 19272 9818
rect 19296 9766 19326 9818
rect 19326 9766 19338 9818
rect 19338 9766 19352 9818
rect 19376 9766 19390 9818
rect 19390 9766 19402 9818
rect 19402 9766 19432 9818
rect 19456 9766 19466 9818
rect 19466 9766 19512 9818
rect 19216 9764 19272 9766
rect 19296 9764 19352 9766
rect 19376 9764 19432 9766
rect 19456 9764 19512 9766
rect 19216 8730 19272 8732
rect 19296 8730 19352 8732
rect 19376 8730 19432 8732
rect 19456 8730 19512 8732
rect 19216 8678 19262 8730
rect 19262 8678 19272 8730
rect 19296 8678 19326 8730
rect 19326 8678 19338 8730
rect 19338 8678 19352 8730
rect 19376 8678 19390 8730
rect 19390 8678 19402 8730
rect 19402 8678 19432 8730
rect 19456 8678 19466 8730
rect 19466 8678 19512 8730
rect 19216 8676 19272 8678
rect 19296 8676 19352 8678
rect 19376 8676 19432 8678
rect 19456 8676 19512 8678
rect 19216 7642 19272 7644
rect 19296 7642 19352 7644
rect 19376 7642 19432 7644
rect 19456 7642 19512 7644
rect 19216 7590 19262 7642
rect 19262 7590 19272 7642
rect 19296 7590 19326 7642
rect 19326 7590 19338 7642
rect 19338 7590 19352 7642
rect 19376 7590 19390 7642
rect 19390 7590 19402 7642
rect 19402 7590 19432 7642
rect 19456 7590 19466 7642
rect 19466 7590 19512 7642
rect 19216 7588 19272 7590
rect 19296 7588 19352 7590
rect 19376 7588 19432 7590
rect 19456 7588 19512 7590
rect 19216 6554 19272 6556
rect 19296 6554 19352 6556
rect 19376 6554 19432 6556
rect 19456 6554 19512 6556
rect 19216 6502 19262 6554
rect 19262 6502 19272 6554
rect 19296 6502 19326 6554
rect 19326 6502 19338 6554
rect 19338 6502 19352 6554
rect 19376 6502 19390 6554
rect 19390 6502 19402 6554
rect 19402 6502 19432 6554
rect 19456 6502 19466 6554
rect 19466 6502 19512 6554
rect 19216 6500 19272 6502
rect 19296 6500 19352 6502
rect 19376 6500 19432 6502
rect 19456 6500 19512 6502
rect 21638 15816 21694 15872
rect 22098 16088 22154 16144
rect 22466 16768 22522 16824
rect 21822 15564 21878 15600
rect 21822 15544 21824 15564
rect 21824 15544 21876 15564
rect 21876 15544 21878 15564
rect 22742 16088 22798 16144
rect 21730 14184 21786 14240
rect 22098 14184 22154 14240
rect 19876 10362 19932 10364
rect 19956 10362 20012 10364
rect 20036 10362 20092 10364
rect 20116 10362 20172 10364
rect 19876 10310 19922 10362
rect 19922 10310 19932 10362
rect 19956 10310 19986 10362
rect 19986 10310 19998 10362
rect 19998 10310 20012 10362
rect 20036 10310 20050 10362
rect 20050 10310 20062 10362
rect 20062 10310 20092 10362
rect 20116 10310 20126 10362
rect 20126 10310 20172 10362
rect 19876 10308 19932 10310
rect 19956 10308 20012 10310
rect 20036 10308 20092 10310
rect 20116 10308 20172 10310
rect 19876 9274 19932 9276
rect 19956 9274 20012 9276
rect 20036 9274 20092 9276
rect 20116 9274 20172 9276
rect 19876 9222 19922 9274
rect 19922 9222 19932 9274
rect 19956 9222 19986 9274
rect 19986 9222 19998 9274
rect 19998 9222 20012 9274
rect 20036 9222 20050 9274
rect 20050 9222 20062 9274
rect 20062 9222 20092 9274
rect 20116 9222 20126 9274
rect 20126 9222 20172 9274
rect 19876 9220 19932 9222
rect 19956 9220 20012 9222
rect 20036 9220 20092 9222
rect 20116 9220 20172 9222
rect 19876 8186 19932 8188
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 19876 8134 19922 8186
rect 19922 8134 19932 8186
rect 19956 8134 19986 8186
rect 19986 8134 19998 8186
rect 19998 8134 20012 8186
rect 20036 8134 20050 8186
rect 20050 8134 20062 8186
rect 20062 8134 20092 8186
rect 20116 8134 20126 8186
rect 20126 8134 20172 8186
rect 19876 8132 19932 8134
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 19876 7098 19932 7100
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 19876 7046 19922 7098
rect 19922 7046 19932 7098
rect 19956 7046 19986 7098
rect 19986 7046 19998 7098
rect 19998 7046 20012 7098
rect 20036 7046 20050 7098
rect 20050 7046 20062 7098
rect 20062 7046 20092 7098
rect 20116 7046 20126 7098
rect 20126 7046 20172 7098
rect 19876 7044 19932 7046
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20626 7284 20628 7304
rect 20628 7284 20680 7304
rect 20680 7284 20682 7304
rect 20626 7248 20682 7284
rect 19216 5466 19272 5468
rect 19296 5466 19352 5468
rect 19376 5466 19432 5468
rect 19456 5466 19512 5468
rect 19216 5414 19262 5466
rect 19262 5414 19272 5466
rect 19296 5414 19326 5466
rect 19326 5414 19338 5466
rect 19338 5414 19352 5466
rect 19376 5414 19390 5466
rect 19390 5414 19402 5466
rect 19402 5414 19432 5466
rect 19456 5414 19466 5466
rect 19466 5414 19512 5466
rect 19216 5412 19272 5414
rect 19296 5412 19352 5414
rect 19376 5412 19432 5414
rect 19456 5412 19512 5414
rect 22926 15952 22982 16008
rect 22650 14456 22706 14512
rect 22558 13912 22614 13968
rect 24674 18672 24730 18728
rect 24398 16632 24454 16688
rect 24582 15680 24638 15736
rect 28998 21800 29054 21856
rect 27650 21242 27706 21244
rect 27730 21242 27786 21244
rect 27810 21242 27866 21244
rect 27890 21242 27946 21244
rect 27650 21190 27696 21242
rect 27696 21190 27706 21242
rect 27730 21190 27760 21242
rect 27760 21190 27772 21242
rect 27772 21190 27786 21242
rect 27810 21190 27824 21242
rect 27824 21190 27836 21242
rect 27836 21190 27866 21242
rect 27890 21190 27900 21242
rect 27900 21190 27946 21242
rect 27650 21188 27706 21190
rect 27730 21188 27786 21190
rect 27810 21188 27866 21190
rect 27890 21188 27946 21190
rect 26990 20698 27046 20700
rect 27070 20698 27126 20700
rect 27150 20698 27206 20700
rect 27230 20698 27286 20700
rect 26990 20646 27036 20698
rect 27036 20646 27046 20698
rect 27070 20646 27100 20698
rect 27100 20646 27112 20698
rect 27112 20646 27126 20698
rect 27150 20646 27164 20698
rect 27164 20646 27176 20698
rect 27176 20646 27206 20698
rect 27230 20646 27240 20698
rect 27240 20646 27286 20698
rect 26990 20644 27046 20646
rect 27070 20644 27126 20646
rect 27150 20644 27206 20646
rect 27230 20644 27286 20646
rect 27650 20154 27706 20156
rect 27730 20154 27786 20156
rect 27810 20154 27866 20156
rect 27890 20154 27946 20156
rect 27650 20102 27696 20154
rect 27696 20102 27706 20154
rect 27730 20102 27760 20154
rect 27760 20102 27772 20154
rect 27772 20102 27786 20154
rect 27810 20102 27824 20154
rect 27824 20102 27836 20154
rect 27836 20102 27866 20154
rect 27890 20102 27900 20154
rect 27900 20102 27946 20154
rect 27650 20100 27706 20102
rect 27730 20100 27786 20102
rect 27810 20100 27866 20102
rect 27890 20100 27946 20102
rect 26514 19896 26570 19952
rect 27526 19932 27528 19952
rect 27528 19932 27580 19952
rect 27580 19932 27582 19952
rect 27526 19896 27582 19932
rect 25318 18128 25374 18184
rect 24398 14320 24454 14376
rect 25870 17992 25926 18048
rect 26146 16768 26202 16824
rect 26238 14320 26294 14376
rect 19876 6010 19932 6012
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 19876 5958 19922 6010
rect 19922 5958 19932 6010
rect 19956 5958 19986 6010
rect 19986 5958 19998 6010
rect 19998 5958 20012 6010
rect 20036 5958 20050 6010
rect 20050 5958 20062 6010
rect 20062 5958 20092 6010
rect 20116 5958 20126 6010
rect 20126 5958 20172 6010
rect 19876 5956 19932 5958
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 19876 4922 19932 4924
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 19876 4870 19922 4922
rect 19922 4870 19932 4922
rect 19956 4870 19986 4922
rect 19986 4870 19998 4922
rect 19998 4870 20012 4922
rect 20036 4870 20050 4922
rect 20050 4870 20062 4922
rect 20062 4870 20092 4922
rect 20116 4870 20126 4922
rect 20126 4870 20172 4922
rect 19876 4868 19932 4870
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 19216 4378 19272 4380
rect 19296 4378 19352 4380
rect 19376 4378 19432 4380
rect 19456 4378 19512 4380
rect 19216 4326 19262 4378
rect 19262 4326 19272 4378
rect 19296 4326 19326 4378
rect 19326 4326 19338 4378
rect 19338 4326 19352 4378
rect 19376 4326 19390 4378
rect 19390 4326 19402 4378
rect 19402 4326 19432 4378
rect 19456 4326 19466 4378
rect 19466 4326 19512 4378
rect 19216 4324 19272 4326
rect 19296 4324 19352 4326
rect 19376 4324 19432 4326
rect 19456 4324 19512 4326
rect 19216 3290 19272 3292
rect 19296 3290 19352 3292
rect 19376 3290 19432 3292
rect 19456 3290 19512 3292
rect 19216 3238 19262 3290
rect 19262 3238 19272 3290
rect 19296 3238 19326 3290
rect 19326 3238 19338 3290
rect 19338 3238 19352 3290
rect 19376 3238 19390 3290
rect 19390 3238 19402 3290
rect 19402 3238 19432 3290
rect 19456 3238 19466 3290
rect 19466 3238 19512 3290
rect 19216 3236 19272 3238
rect 19296 3236 19352 3238
rect 19376 3236 19432 3238
rect 19456 3236 19512 3238
rect 19876 3834 19932 3836
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 19876 3782 19922 3834
rect 19922 3782 19932 3834
rect 19956 3782 19986 3834
rect 19986 3782 19998 3834
rect 19998 3782 20012 3834
rect 20036 3782 20050 3834
rect 20050 3782 20062 3834
rect 20062 3782 20092 3834
rect 20116 3782 20126 3834
rect 20126 3782 20172 3834
rect 19876 3780 19932 3782
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 26990 19610 27046 19612
rect 27070 19610 27126 19612
rect 27150 19610 27206 19612
rect 27230 19610 27286 19612
rect 26990 19558 27036 19610
rect 27036 19558 27046 19610
rect 27070 19558 27100 19610
rect 27100 19558 27112 19610
rect 27112 19558 27126 19610
rect 27150 19558 27164 19610
rect 27164 19558 27176 19610
rect 27176 19558 27206 19610
rect 27230 19558 27240 19610
rect 27240 19558 27286 19610
rect 26990 19556 27046 19558
rect 27070 19556 27126 19558
rect 27150 19556 27206 19558
rect 27230 19556 27286 19558
rect 27650 19066 27706 19068
rect 27730 19066 27786 19068
rect 27810 19066 27866 19068
rect 27890 19066 27946 19068
rect 27650 19014 27696 19066
rect 27696 19014 27706 19066
rect 27730 19014 27760 19066
rect 27760 19014 27772 19066
rect 27772 19014 27786 19066
rect 27810 19014 27824 19066
rect 27824 19014 27836 19066
rect 27836 19014 27866 19066
rect 27890 19014 27900 19066
rect 27900 19014 27946 19066
rect 27650 19012 27706 19014
rect 27730 19012 27786 19014
rect 27810 19012 27866 19014
rect 27890 19012 27946 19014
rect 26990 18522 27046 18524
rect 27070 18522 27126 18524
rect 27150 18522 27206 18524
rect 27230 18522 27286 18524
rect 26990 18470 27036 18522
rect 27036 18470 27046 18522
rect 27070 18470 27100 18522
rect 27100 18470 27112 18522
rect 27112 18470 27126 18522
rect 27150 18470 27164 18522
rect 27164 18470 27176 18522
rect 27176 18470 27206 18522
rect 27230 18470 27240 18522
rect 27240 18470 27286 18522
rect 26990 18468 27046 18470
rect 27070 18468 27126 18470
rect 27150 18468 27206 18470
rect 27230 18468 27286 18470
rect 27526 18828 27582 18864
rect 27526 18808 27528 18828
rect 27528 18808 27580 18828
rect 27580 18808 27582 18828
rect 28078 17992 28134 18048
rect 27650 17978 27706 17980
rect 27730 17978 27786 17980
rect 27810 17978 27866 17980
rect 27890 17978 27946 17980
rect 27650 17926 27696 17978
rect 27696 17926 27706 17978
rect 27730 17926 27760 17978
rect 27760 17926 27772 17978
rect 27772 17926 27786 17978
rect 27810 17926 27824 17978
rect 27824 17926 27836 17978
rect 27836 17926 27866 17978
rect 27890 17926 27900 17978
rect 27900 17926 27946 17978
rect 27650 17924 27706 17926
rect 27730 17924 27786 17926
rect 27810 17924 27866 17926
rect 27890 17924 27946 17926
rect 26990 17434 27046 17436
rect 27070 17434 27126 17436
rect 27150 17434 27206 17436
rect 27230 17434 27286 17436
rect 26990 17382 27036 17434
rect 27036 17382 27046 17434
rect 27070 17382 27100 17434
rect 27100 17382 27112 17434
rect 27112 17382 27126 17434
rect 27150 17382 27164 17434
rect 27164 17382 27176 17434
rect 27176 17382 27206 17434
rect 27230 17382 27240 17434
rect 27240 17382 27286 17434
rect 26990 17380 27046 17382
rect 27070 17380 27126 17382
rect 27150 17380 27206 17382
rect 27230 17380 27286 17382
rect 26606 16768 26662 16824
rect 26990 16346 27046 16348
rect 27070 16346 27126 16348
rect 27150 16346 27206 16348
rect 27230 16346 27286 16348
rect 26990 16294 27036 16346
rect 27036 16294 27046 16346
rect 27070 16294 27100 16346
rect 27100 16294 27112 16346
rect 27112 16294 27126 16346
rect 27150 16294 27164 16346
rect 27164 16294 27176 16346
rect 27176 16294 27206 16346
rect 27230 16294 27240 16346
rect 27240 16294 27286 16346
rect 26990 16292 27046 16294
rect 27070 16292 27126 16294
rect 27150 16292 27206 16294
rect 27230 16292 27286 16294
rect 26990 15258 27046 15260
rect 27070 15258 27126 15260
rect 27150 15258 27206 15260
rect 27230 15258 27286 15260
rect 26990 15206 27036 15258
rect 27036 15206 27046 15258
rect 27070 15206 27100 15258
rect 27100 15206 27112 15258
rect 27112 15206 27126 15258
rect 27150 15206 27164 15258
rect 27164 15206 27176 15258
rect 27176 15206 27206 15258
rect 27230 15206 27240 15258
rect 27240 15206 27286 15258
rect 26990 15204 27046 15206
rect 27070 15204 27126 15206
rect 27150 15204 27206 15206
rect 27230 15204 27286 15206
rect 26974 14320 27030 14376
rect 26990 14170 27046 14172
rect 27070 14170 27126 14172
rect 27150 14170 27206 14172
rect 27230 14170 27286 14172
rect 26990 14118 27036 14170
rect 27036 14118 27046 14170
rect 27070 14118 27100 14170
rect 27100 14118 27112 14170
rect 27112 14118 27126 14170
rect 27150 14118 27164 14170
rect 27164 14118 27176 14170
rect 27176 14118 27206 14170
rect 27230 14118 27240 14170
rect 27240 14118 27286 14170
rect 26990 14116 27046 14118
rect 27070 14116 27126 14118
rect 27150 14116 27206 14118
rect 27230 14116 27286 14118
rect 27650 16890 27706 16892
rect 27730 16890 27786 16892
rect 27810 16890 27866 16892
rect 27890 16890 27946 16892
rect 27650 16838 27696 16890
rect 27696 16838 27706 16890
rect 27730 16838 27760 16890
rect 27760 16838 27772 16890
rect 27772 16838 27786 16890
rect 27810 16838 27824 16890
rect 27824 16838 27836 16890
rect 27836 16838 27866 16890
rect 27890 16838 27900 16890
rect 27900 16838 27946 16890
rect 27650 16836 27706 16838
rect 27730 16836 27786 16838
rect 27810 16836 27866 16838
rect 27890 16836 27946 16838
rect 27650 15802 27706 15804
rect 27730 15802 27786 15804
rect 27810 15802 27866 15804
rect 27890 15802 27946 15804
rect 27650 15750 27696 15802
rect 27696 15750 27706 15802
rect 27730 15750 27760 15802
rect 27760 15750 27772 15802
rect 27772 15750 27786 15802
rect 27810 15750 27824 15802
rect 27824 15750 27836 15802
rect 27836 15750 27866 15802
rect 27890 15750 27900 15802
rect 27900 15750 27946 15802
rect 27650 15748 27706 15750
rect 27730 15748 27786 15750
rect 27810 15748 27866 15750
rect 27890 15748 27946 15750
rect 27650 14714 27706 14716
rect 27730 14714 27786 14716
rect 27810 14714 27866 14716
rect 27890 14714 27946 14716
rect 27650 14662 27696 14714
rect 27696 14662 27706 14714
rect 27730 14662 27760 14714
rect 27760 14662 27772 14714
rect 27772 14662 27786 14714
rect 27810 14662 27824 14714
rect 27824 14662 27836 14714
rect 27836 14662 27866 14714
rect 27890 14662 27900 14714
rect 27900 14662 27946 14714
rect 27650 14660 27706 14662
rect 27730 14660 27786 14662
rect 27810 14660 27866 14662
rect 27890 14660 27946 14662
rect 26990 13082 27046 13084
rect 27070 13082 27126 13084
rect 27150 13082 27206 13084
rect 27230 13082 27286 13084
rect 26990 13030 27036 13082
rect 27036 13030 27046 13082
rect 27070 13030 27100 13082
rect 27100 13030 27112 13082
rect 27112 13030 27126 13082
rect 27150 13030 27164 13082
rect 27164 13030 27176 13082
rect 27176 13030 27206 13082
rect 27230 13030 27240 13082
rect 27240 13030 27286 13082
rect 26990 13028 27046 13030
rect 27070 13028 27126 13030
rect 27150 13028 27206 13030
rect 27230 13028 27286 13030
rect 27650 13626 27706 13628
rect 27730 13626 27786 13628
rect 27810 13626 27866 13628
rect 27890 13626 27946 13628
rect 27650 13574 27696 13626
rect 27696 13574 27706 13626
rect 27730 13574 27760 13626
rect 27760 13574 27772 13626
rect 27772 13574 27786 13626
rect 27810 13574 27824 13626
rect 27824 13574 27836 13626
rect 27836 13574 27866 13626
rect 27890 13574 27900 13626
rect 27900 13574 27946 13626
rect 27650 13572 27706 13574
rect 27730 13572 27786 13574
rect 27810 13572 27866 13574
rect 27890 13572 27946 13574
rect 27650 12538 27706 12540
rect 27730 12538 27786 12540
rect 27810 12538 27866 12540
rect 27890 12538 27946 12540
rect 27650 12486 27696 12538
rect 27696 12486 27706 12538
rect 27730 12486 27760 12538
rect 27760 12486 27772 12538
rect 27772 12486 27786 12538
rect 27810 12486 27824 12538
rect 27824 12486 27836 12538
rect 27836 12486 27866 12538
rect 27890 12486 27900 12538
rect 27900 12486 27946 12538
rect 27650 12484 27706 12486
rect 27730 12484 27786 12486
rect 27810 12484 27866 12486
rect 27890 12484 27946 12486
rect 26990 11994 27046 11996
rect 27070 11994 27126 11996
rect 27150 11994 27206 11996
rect 27230 11994 27286 11996
rect 26990 11942 27036 11994
rect 27036 11942 27046 11994
rect 27070 11942 27100 11994
rect 27100 11942 27112 11994
rect 27112 11942 27126 11994
rect 27150 11942 27164 11994
rect 27164 11942 27176 11994
rect 27176 11942 27206 11994
rect 27230 11942 27240 11994
rect 27240 11942 27286 11994
rect 26990 11940 27046 11942
rect 27070 11940 27126 11942
rect 27150 11940 27206 11942
rect 27230 11940 27286 11942
rect 28262 14476 28318 14512
rect 28262 14456 28264 14476
rect 28264 14456 28316 14476
rect 28316 14456 28318 14476
rect 28354 14320 28410 14376
rect 28262 13912 28318 13968
rect 30194 18828 30250 18864
rect 30194 18808 30196 18828
rect 30196 18808 30248 18828
rect 30248 18808 30250 18828
rect 30194 13912 30250 13968
rect 27066 11620 27122 11656
rect 27066 11600 27068 11620
rect 27068 11600 27120 11620
rect 27120 11600 27122 11620
rect 27650 11450 27706 11452
rect 27730 11450 27786 11452
rect 27810 11450 27866 11452
rect 27890 11450 27946 11452
rect 27650 11398 27696 11450
rect 27696 11398 27706 11450
rect 27730 11398 27760 11450
rect 27760 11398 27772 11450
rect 27772 11398 27786 11450
rect 27810 11398 27824 11450
rect 27824 11398 27836 11450
rect 27836 11398 27866 11450
rect 27890 11398 27900 11450
rect 27900 11398 27946 11450
rect 27650 11396 27706 11398
rect 27730 11396 27786 11398
rect 27810 11396 27866 11398
rect 27890 11396 27946 11398
rect 26990 10906 27046 10908
rect 27070 10906 27126 10908
rect 27150 10906 27206 10908
rect 27230 10906 27286 10908
rect 26990 10854 27036 10906
rect 27036 10854 27046 10906
rect 27070 10854 27100 10906
rect 27100 10854 27112 10906
rect 27112 10854 27126 10906
rect 27150 10854 27164 10906
rect 27164 10854 27176 10906
rect 27176 10854 27206 10906
rect 27230 10854 27240 10906
rect 27240 10854 27286 10906
rect 26990 10852 27046 10854
rect 27070 10852 27126 10854
rect 27150 10852 27206 10854
rect 27230 10852 27286 10854
rect 27650 10362 27706 10364
rect 27730 10362 27786 10364
rect 27810 10362 27866 10364
rect 27890 10362 27946 10364
rect 27650 10310 27696 10362
rect 27696 10310 27706 10362
rect 27730 10310 27760 10362
rect 27760 10310 27772 10362
rect 27772 10310 27786 10362
rect 27810 10310 27824 10362
rect 27824 10310 27836 10362
rect 27836 10310 27866 10362
rect 27890 10310 27900 10362
rect 27900 10310 27946 10362
rect 27650 10308 27706 10310
rect 27730 10308 27786 10310
rect 27810 10308 27866 10310
rect 27890 10308 27946 10310
rect 26990 9818 27046 9820
rect 27070 9818 27126 9820
rect 27150 9818 27206 9820
rect 27230 9818 27286 9820
rect 26990 9766 27036 9818
rect 27036 9766 27046 9818
rect 27070 9766 27100 9818
rect 27100 9766 27112 9818
rect 27112 9766 27126 9818
rect 27150 9766 27164 9818
rect 27164 9766 27176 9818
rect 27176 9766 27206 9818
rect 27230 9766 27240 9818
rect 27240 9766 27286 9818
rect 26990 9764 27046 9766
rect 27070 9764 27126 9766
rect 27150 9764 27206 9766
rect 27230 9764 27286 9766
rect 26990 8730 27046 8732
rect 27070 8730 27126 8732
rect 27150 8730 27206 8732
rect 27230 8730 27286 8732
rect 26990 8678 27036 8730
rect 27036 8678 27046 8730
rect 27070 8678 27100 8730
rect 27100 8678 27112 8730
rect 27112 8678 27126 8730
rect 27150 8678 27164 8730
rect 27164 8678 27176 8730
rect 27176 8678 27206 8730
rect 27230 8678 27240 8730
rect 27240 8678 27286 8730
rect 26990 8676 27046 8678
rect 27070 8676 27126 8678
rect 27150 8676 27206 8678
rect 27230 8676 27286 8678
rect 27650 9274 27706 9276
rect 27730 9274 27786 9276
rect 27810 9274 27866 9276
rect 27890 9274 27946 9276
rect 27650 9222 27696 9274
rect 27696 9222 27706 9274
rect 27730 9222 27760 9274
rect 27760 9222 27772 9274
rect 27772 9222 27786 9274
rect 27810 9222 27824 9274
rect 27824 9222 27836 9274
rect 27836 9222 27866 9274
rect 27890 9222 27900 9274
rect 27900 9222 27946 9274
rect 27650 9220 27706 9222
rect 27730 9220 27786 9222
rect 27810 9220 27866 9222
rect 27890 9220 27946 9222
rect 27650 8186 27706 8188
rect 27730 8186 27786 8188
rect 27810 8186 27866 8188
rect 27890 8186 27946 8188
rect 27650 8134 27696 8186
rect 27696 8134 27706 8186
rect 27730 8134 27760 8186
rect 27760 8134 27772 8186
rect 27772 8134 27786 8186
rect 27810 8134 27824 8186
rect 27824 8134 27836 8186
rect 27836 8134 27866 8186
rect 27890 8134 27900 8186
rect 27900 8134 27946 8186
rect 27650 8132 27706 8134
rect 27730 8132 27786 8134
rect 27810 8132 27866 8134
rect 27890 8132 27946 8134
rect 26990 7642 27046 7644
rect 27070 7642 27126 7644
rect 27150 7642 27206 7644
rect 27230 7642 27286 7644
rect 26990 7590 27036 7642
rect 27036 7590 27046 7642
rect 27070 7590 27100 7642
rect 27100 7590 27112 7642
rect 27112 7590 27126 7642
rect 27150 7590 27164 7642
rect 27164 7590 27176 7642
rect 27176 7590 27206 7642
rect 27230 7590 27240 7642
rect 27240 7590 27286 7642
rect 26990 7588 27046 7590
rect 27070 7588 27126 7590
rect 27150 7588 27206 7590
rect 27230 7588 27286 7590
rect 19876 2746 19932 2748
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 19876 2694 19922 2746
rect 19922 2694 19932 2746
rect 19956 2694 19986 2746
rect 19986 2694 19998 2746
rect 19998 2694 20012 2746
rect 20036 2694 20050 2746
rect 20050 2694 20062 2746
rect 20062 2694 20092 2746
rect 20116 2694 20126 2746
rect 20126 2694 20172 2746
rect 19876 2692 19932 2694
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 19216 2202 19272 2204
rect 19296 2202 19352 2204
rect 19376 2202 19432 2204
rect 19456 2202 19512 2204
rect 19216 2150 19262 2202
rect 19262 2150 19272 2202
rect 19296 2150 19326 2202
rect 19326 2150 19338 2202
rect 19338 2150 19352 2202
rect 19376 2150 19390 2202
rect 19390 2150 19402 2202
rect 19402 2150 19432 2202
rect 19456 2150 19466 2202
rect 19466 2150 19512 2202
rect 19216 2148 19272 2150
rect 19296 2148 19352 2150
rect 19376 2148 19432 2150
rect 19456 2148 19512 2150
rect 19876 1658 19932 1660
rect 19956 1658 20012 1660
rect 20036 1658 20092 1660
rect 20116 1658 20172 1660
rect 19876 1606 19922 1658
rect 19922 1606 19932 1658
rect 19956 1606 19986 1658
rect 19986 1606 19998 1658
rect 19998 1606 20012 1658
rect 20036 1606 20050 1658
rect 20050 1606 20062 1658
rect 20062 1606 20092 1658
rect 20116 1606 20126 1658
rect 20126 1606 20172 1658
rect 19876 1604 19932 1606
rect 19956 1604 20012 1606
rect 20036 1604 20092 1606
rect 20116 1604 20172 1606
rect 26990 6554 27046 6556
rect 27070 6554 27126 6556
rect 27150 6554 27206 6556
rect 27230 6554 27286 6556
rect 26990 6502 27036 6554
rect 27036 6502 27046 6554
rect 27070 6502 27100 6554
rect 27100 6502 27112 6554
rect 27112 6502 27126 6554
rect 27150 6502 27164 6554
rect 27164 6502 27176 6554
rect 27176 6502 27206 6554
rect 27230 6502 27240 6554
rect 27240 6502 27286 6554
rect 26990 6500 27046 6502
rect 27070 6500 27126 6502
rect 27150 6500 27206 6502
rect 27230 6500 27286 6502
rect 27650 7098 27706 7100
rect 27730 7098 27786 7100
rect 27810 7098 27866 7100
rect 27890 7098 27946 7100
rect 27650 7046 27696 7098
rect 27696 7046 27706 7098
rect 27730 7046 27760 7098
rect 27760 7046 27772 7098
rect 27772 7046 27786 7098
rect 27810 7046 27824 7098
rect 27824 7046 27836 7098
rect 27836 7046 27866 7098
rect 27890 7046 27900 7098
rect 27900 7046 27946 7098
rect 27650 7044 27706 7046
rect 27730 7044 27786 7046
rect 27810 7044 27866 7046
rect 27890 7044 27946 7046
rect 26990 5466 27046 5468
rect 27070 5466 27126 5468
rect 27150 5466 27206 5468
rect 27230 5466 27286 5468
rect 26990 5414 27036 5466
rect 27036 5414 27046 5466
rect 27070 5414 27100 5466
rect 27100 5414 27112 5466
rect 27112 5414 27126 5466
rect 27150 5414 27164 5466
rect 27164 5414 27176 5466
rect 27176 5414 27206 5466
rect 27230 5414 27240 5466
rect 27240 5414 27286 5466
rect 26990 5412 27046 5414
rect 27070 5412 27126 5414
rect 27150 5412 27206 5414
rect 27230 5412 27286 5414
rect 27650 6010 27706 6012
rect 27730 6010 27786 6012
rect 27810 6010 27866 6012
rect 27890 6010 27946 6012
rect 27650 5958 27696 6010
rect 27696 5958 27706 6010
rect 27730 5958 27760 6010
rect 27760 5958 27772 6010
rect 27772 5958 27786 6010
rect 27810 5958 27824 6010
rect 27824 5958 27836 6010
rect 27836 5958 27866 6010
rect 27890 5958 27900 6010
rect 27900 5958 27946 6010
rect 27650 5956 27706 5958
rect 27730 5956 27786 5958
rect 27810 5956 27866 5958
rect 27890 5956 27946 5958
rect 27650 4922 27706 4924
rect 27730 4922 27786 4924
rect 27810 4922 27866 4924
rect 27890 4922 27946 4924
rect 27650 4870 27696 4922
rect 27696 4870 27706 4922
rect 27730 4870 27760 4922
rect 27760 4870 27772 4922
rect 27772 4870 27786 4922
rect 27810 4870 27824 4922
rect 27824 4870 27836 4922
rect 27836 4870 27866 4922
rect 27890 4870 27900 4922
rect 27900 4870 27946 4922
rect 27650 4868 27706 4870
rect 27730 4868 27786 4870
rect 27810 4868 27866 4870
rect 27890 4868 27946 4870
rect 26990 4378 27046 4380
rect 27070 4378 27126 4380
rect 27150 4378 27206 4380
rect 27230 4378 27286 4380
rect 26990 4326 27036 4378
rect 27036 4326 27046 4378
rect 27070 4326 27100 4378
rect 27100 4326 27112 4378
rect 27112 4326 27126 4378
rect 27150 4326 27164 4378
rect 27164 4326 27176 4378
rect 27176 4326 27206 4378
rect 27230 4326 27240 4378
rect 27240 4326 27286 4378
rect 26990 4324 27046 4326
rect 27070 4324 27126 4326
rect 27150 4324 27206 4326
rect 27230 4324 27286 4326
rect 27650 3834 27706 3836
rect 27730 3834 27786 3836
rect 27810 3834 27866 3836
rect 27890 3834 27946 3836
rect 27650 3782 27696 3834
rect 27696 3782 27706 3834
rect 27730 3782 27760 3834
rect 27760 3782 27772 3834
rect 27772 3782 27786 3834
rect 27810 3782 27824 3834
rect 27824 3782 27836 3834
rect 27836 3782 27866 3834
rect 27890 3782 27900 3834
rect 27900 3782 27946 3834
rect 27650 3780 27706 3782
rect 27730 3780 27786 3782
rect 27810 3780 27866 3782
rect 27890 3780 27946 3782
rect 26990 3290 27046 3292
rect 27070 3290 27126 3292
rect 27150 3290 27206 3292
rect 27230 3290 27286 3292
rect 26990 3238 27036 3290
rect 27036 3238 27046 3290
rect 27070 3238 27100 3290
rect 27100 3238 27112 3290
rect 27112 3238 27126 3290
rect 27150 3238 27164 3290
rect 27164 3238 27176 3290
rect 27176 3238 27206 3290
rect 27230 3238 27240 3290
rect 27240 3238 27286 3290
rect 26990 3236 27046 3238
rect 27070 3236 27126 3238
rect 27150 3236 27206 3238
rect 27230 3236 27286 3238
rect 19216 1114 19272 1116
rect 19296 1114 19352 1116
rect 19376 1114 19432 1116
rect 19456 1114 19512 1116
rect 19216 1062 19262 1114
rect 19262 1062 19272 1114
rect 19296 1062 19326 1114
rect 19326 1062 19338 1114
rect 19338 1062 19352 1114
rect 19376 1062 19390 1114
rect 19390 1062 19402 1114
rect 19402 1062 19432 1114
rect 19456 1062 19466 1114
rect 19466 1062 19512 1114
rect 19216 1060 19272 1062
rect 19296 1060 19352 1062
rect 19376 1060 19432 1062
rect 19456 1060 19512 1062
rect 21454 2388 21456 2408
rect 21456 2388 21508 2408
rect 21508 2388 21510 2408
rect 21454 2352 21510 2388
rect 22098 2372 22154 2408
rect 22098 2352 22100 2372
rect 22100 2352 22152 2372
rect 22152 2352 22154 2372
rect 26698 2932 26700 2952
rect 26700 2932 26752 2952
rect 26752 2932 26754 2952
rect 26698 2896 26754 2932
rect 26990 2202 27046 2204
rect 27070 2202 27126 2204
rect 27150 2202 27206 2204
rect 27230 2202 27286 2204
rect 26990 2150 27036 2202
rect 27036 2150 27046 2202
rect 27070 2150 27100 2202
rect 27100 2150 27112 2202
rect 27112 2150 27126 2202
rect 27150 2150 27164 2202
rect 27164 2150 27176 2202
rect 27176 2150 27206 2202
rect 27230 2150 27240 2202
rect 27240 2150 27286 2202
rect 26990 2148 27046 2150
rect 27070 2148 27126 2150
rect 27150 2148 27206 2150
rect 27230 2148 27286 2150
rect 28814 2932 28816 2952
rect 28816 2932 28868 2952
rect 28868 2932 28870 2952
rect 28814 2896 28870 2932
rect 27650 2746 27706 2748
rect 27730 2746 27786 2748
rect 27810 2746 27866 2748
rect 27890 2746 27946 2748
rect 27650 2694 27696 2746
rect 27696 2694 27706 2746
rect 27730 2694 27760 2746
rect 27760 2694 27772 2746
rect 27772 2694 27786 2746
rect 27810 2694 27824 2746
rect 27824 2694 27836 2746
rect 27836 2694 27866 2746
rect 27890 2694 27900 2746
rect 27900 2694 27946 2746
rect 27650 2692 27706 2694
rect 27730 2692 27786 2694
rect 27810 2692 27866 2694
rect 27890 2692 27946 2694
rect 27650 1658 27706 1660
rect 27730 1658 27786 1660
rect 27810 1658 27866 1660
rect 27890 1658 27946 1660
rect 27650 1606 27696 1658
rect 27696 1606 27706 1658
rect 27730 1606 27760 1658
rect 27760 1606 27772 1658
rect 27772 1606 27786 1658
rect 27810 1606 27824 1658
rect 27824 1606 27836 1658
rect 27836 1606 27866 1658
rect 27890 1606 27900 1658
rect 27900 1606 27946 1658
rect 27650 1604 27706 1606
rect 27730 1604 27786 1606
rect 27810 1604 27866 1606
rect 27890 1604 27946 1606
rect 26990 1114 27046 1116
rect 27070 1114 27126 1116
rect 27150 1114 27206 1116
rect 27230 1114 27286 1116
rect 26990 1062 27036 1114
rect 27036 1062 27046 1114
rect 27070 1062 27100 1114
rect 27100 1062 27112 1114
rect 27112 1062 27126 1114
rect 27150 1062 27164 1114
rect 27164 1062 27176 1114
rect 27176 1062 27206 1114
rect 27230 1062 27240 1114
rect 27240 1062 27286 1114
rect 26990 1060 27046 1062
rect 27070 1060 27126 1062
rect 27150 1060 27206 1062
rect 27230 1060 27286 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 12102 570 12158 572
rect 12182 570 12238 572
rect 12262 570 12318 572
rect 12342 570 12398 572
rect 12102 518 12148 570
rect 12148 518 12158 570
rect 12182 518 12212 570
rect 12212 518 12224 570
rect 12224 518 12238 570
rect 12262 518 12276 570
rect 12276 518 12288 570
rect 12288 518 12318 570
rect 12342 518 12352 570
rect 12352 518 12398 570
rect 12102 516 12158 518
rect 12182 516 12238 518
rect 12262 516 12318 518
rect 12342 516 12398 518
rect 19876 570 19932 572
rect 19956 570 20012 572
rect 20036 570 20092 572
rect 20116 570 20172 572
rect 19876 518 19922 570
rect 19922 518 19932 570
rect 19956 518 19986 570
rect 19986 518 19998 570
rect 19998 518 20012 570
rect 20036 518 20050 570
rect 20050 518 20062 570
rect 20062 518 20092 570
rect 20116 518 20126 570
rect 20126 518 20172 570
rect 19876 516 19932 518
rect 19956 516 20012 518
rect 20036 516 20092 518
rect 20116 516 20172 518
rect 27650 570 27706 572
rect 27730 570 27786 572
rect 27810 570 27866 572
rect 27890 570 27946 572
rect 27650 518 27696 570
rect 27696 518 27706 570
rect 27730 518 27760 570
rect 27760 518 27772 570
rect 27772 518 27786 570
rect 27810 518 27824 570
rect 27824 518 27836 570
rect 27836 518 27866 570
rect 27890 518 27900 570
rect 27900 518 27946 570
rect 27650 516 27706 518
rect 27730 516 27786 518
rect 27810 516 27866 518
rect 27890 516 27946 518
<< metal3 >>
rect 11646 21932 11652 21996
rect 11716 21994 11722 21996
rect 11789 21994 11855 21997
rect 12249 21996 12315 21997
rect 23841 21996 23907 21997
rect 24945 21996 25011 21997
rect 25497 21996 25563 21997
rect 26049 21996 26115 21997
rect 11716 21992 11855 21994
rect 11716 21936 11794 21992
rect 11850 21936 11855 21992
rect 11716 21934 11855 21936
rect 11716 21932 11722 21934
rect 11789 21931 11855 21934
rect 12198 21932 12204 21996
rect 12268 21994 12315 21996
rect 23790 21994 23796 21996
rect 12268 21992 12360 21994
rect 12310 21936 12360 21992
rect 12268 21934 12360 21936
rect 23750 21934 23796 21994
rect 23860 21992 23907 21996
rect 24894 21994 24900 21996
rect 23902 21936 23907 21992
rect 12268 21932 12315 21934
rect 23790 21932 23796 21934
rect 23860 21932 23907 21936
rect 24854 21934 24900 21994
rect 24964 21992 25011 21996
rect 25446 21994 25452 21996
rect 25006 21936 25011 21992
rect 24894 21932 24900 21934
rect 24964 21932 25011 21936
rect 25406 21934 25452 21994
rect 25516 21992 25563 21996
rect 25998 21994 26004 21996
rect 25558 21936 25563 21992
rect 25446 21932 25452 21934
rect 25516 21932 25563 21936
rect 25958 21934 26004 21994
rect 26068 21992 26115 21996
rect 26110 21936 26115 21992
rect 25998 21932 26004 21934
rect 26068 21932 26115 21936
rect 27102 21932 27108 21996
rect 27172 21994 27178 21996
rect 27521 21994 27587 21997
rect 27172 21992 27587 21994
rect 27172 21936 27526 21992
rect 27582 21936 27587 21992
rect 27172 21934 27587 21936
rect 27172 21932 27178 21934
rect 12249 21931 12315 21932
rect 23841 21931 23907 21932
rect 24945 21931 25011 21932
rect 25497 21931 25563 21932
rect 26049 21931 26115 21932
rect 27521 21931 27587 21934
rect 27654 21932 27660 21996
rect 27724 21994 27730 21996
rect 28257 21994 28323 21997
rect 27724 21992 28323 21994
rect 27724 21936 28262 21992
rect 28318 21936 28323 21992
rect 27724 21934 28323 21936
rect 27724 21932 27730 21934
rect 28257 21931 28323 21934
rect 7782 21796 7788 21860
rect 7852 21858 7858 21860
rect 8661 21858 8727 21861
rect 21633 21860 21699 21861
rect 24393 21860 24459 21861
rect 21582 21858 21588 21860
rect 7852 21856 8727 21858
rect 7852 21800 8666 21856
rect 8722 21800 8727 21856
rect 7852 21798 8727 21800
rect 21542 21798 21588 21858
rect 21652 21856 21699 21860
rect 24342 21858 24348 21860
rect 21694 21800 21699 21856
rect 7852 21796 7858 21798
rect 8661 21795 8727 21798
rect 21582 21796 21588 21798
rect 21652 21796 21699 21800
rect 24302 21798 24348 21858
rect 24412 21856 24459 21860
rect 24454 21800 24459 21856
rect 24342 21796 24348 21798
rect 24412 21796 24459 21800
rect 21633 21795 21699 21796
rect 24393 21795 24459 21796
rect 26509 21860 26575 21861
rect 26509 21856 26556 21860
rect 26620 21858 26626 21860
rect 26509 21800 26514 21856
rect 26509 21796 26556 21800
rect 26620 21798 26666 21858
rect 26620 21796 26626 21798
rect 28206 21796 28212 21860
rect 28276 21858 28282 21860
rect 28993 21858 29059 21861
rect 28276 21856 29059 21858
rect 28276 21800 28998 21856
rect 29054 21800 29059 21856
rect 28276 21798 29059 21800
rect 28276 21796 28282 21798
rect 26509 21795 26575 21796
rect 28993 21795 29059 21798
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 11432 21792 11748 21793
rect 11432 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11748 21792
rect 11432 21727 11748 21728
rect 19206 21792 19522 21793
rect 19206 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19522 21792
rect 19206 21727 19522 21728
rect 26980 21792 27296 21793
rect 26980 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27296 21792
rect 26980 21727 27296 21728
rect 6126 21660 6132 21724
rect 6196 21722 6202 21724
rect 6453 21722 6519 21725
rect 7281 21724 7347 21725
rect 8385 21724 8451 21725
rect 6196 21720 6519 21722
rect 6196 21664 6458 21720
rect 6514 21664 6519 21720
rect 6196 21662 6519 21664
rect 6196 21660 6202 21662
rect 6453 21659 6519 21662
rect 7230 21660 7236 21724
rect 7300 21722 7347 21724
rect 7300 21720 7392 21722
rect 7342 21664 7392 21720
rect 7300 21662 7392 21664
rect 7300 21660 7347 21662
rect 8334 21660 8340 21724
rect 8404 21722 8451 21724
rect 9949 21724 10015 21725
rect 9949 21722 9996 21724
rect 8404 21720 8496 21722
rect 8446 21664 8496 21720
rect 8404 21662 8496 21664
rect 9904 21720 9996 21722
rect 9904 21664 9954 21720
rect 9904 21662 9996 21664
rect 8404 21660 8451 21662
rect 7281 21659 7347 21660
rect 8385 21659 8451 21660
rect 9949 21660 9996 21662
rect 10060 21660 10066 21724
rect 10317 21722 10383 21725
rect 12801 21724 12867 21725
rect 10542 21722 10548 21724
rect 10317 21720 10548 21722
rect 10317 21664 10322 21720
rect 10378 21664 10548 21720
rect 10317 21662 10548 21664
rect 9949 21659 10015 21660
rect 10317 21659 10383 21662
rect 10542 21660 10548 21662
rect 10612 21660 10618 21724
rect 12750 21660 12756 21724
rect 12820 21722 12867 21724
rect 12820 21720 12912 21722
rect 12862 21664 12912 21720
rect 12820 21662 12912 21664
rect 12820 21660 12867 21662
rect 12801 21659 12867 21660
rect 11094 21524 11100 21588
rect 11164 21586 11170 21588
rect 11697 21586 11763 21589
rect 11164 21584 11763 21586
rect 11164 21528 11702 21584
rect 11758 21528 11763 21584
rect 11164 21526 11763 21528
rect 11164 21524 11170 21526
rect 11697 21523 11763 21526
rect 16665 21586 16731 21589
rect 17718 21586 17724 21588
rect 16665 21584 17724 21586
rect 16665 21528 16670 21584
rect 16726 21528 17724 21584
rect 16665 21526 17724 21528
rect 16665 21523 16731 21526
rect 17718 21524 17724 21526
rect 17788 21524 17794 21588
rect 18822 21524 18828 21588
rect 18892 21586 18898 21588
rect 19425 21586 19491 21589
rect 18892 21584 19491 21586
rect 18892 21528 19430 21584
rect 19486 21528 19491 21584
rect 18892 21526 19491 21528
rect 18892 21524 18898 21526
rect 19425 21523 19491 21526
rect 18270 21388 18276 21452
rect 18340 21450 18346 21452
rect 19241 21450 19307 21453
rect 18340 21448 19307 21450
rect 18340 21392 19246 21448
rect 19302 21392 19307 21448
rect 18340 21390 19307 21392
rect 18340 21388 18346 21390
rect 19241 21387 19307 21390
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 12092 21248 12408 21249
rect 12092 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12408 21248
rect 12092 21183 12408 21184
rect 19866 21248 20182 21249
rect 19866 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20182 21248
rect 19866 21183 20182 21184
rect 27640 21248 27956 21249
rect 27640 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27956 21248
rect 27640 21183 27956 21184
rect 6269 21178 6335 21181
rect 6678 21178 6684 21180
rect 6269 21176 6684 21178
rect 6269 21120 6274 21176
rect 6330 21120 6684 21176
rect 6269 21118 6684 21120
rect 6269 21115 6335 21118
rect 6678 21116 6684 21118
rect 6748 21116 6754 21180
rect 8477 21178 8543 21181
rect 13813 21180 13879 21181
rect 9438 21178 9444 21180
rect 8477 21176 9444 21178
rect 8477 21120 8482 21176
rect 8538 21120 9444 21176
rect 8477 21118 9444 21120
rect 8477 21115 8543 21118
rect 9438 21116 9444 21118
rect 9508 21116 9514 21180
rect 13813 21178 13860 21180
rect 13768 21176 13860 21178
rect 13768 21120 13818 21176
rect 13768 21118 13860 21120
rect 13813 21116 13860 21118
rect 13924 21116 13930 21180
rect 13813 21115 13879 21116
rect 15469 21044 15535 21045
rect 15469 21042 15516 21044
rect 15424 21040 15516 21042
rect 15424 20984 15474 21040
rect 15424 20982 15516 20984
rect 15469 20980 15516 20982
rect 15580 20980 15586 21044
rect 15469 20979 15535 20980
rect 16757 20906 16823 20909
rect 18229 20906 18295 20909
rect 22921 20906 22987 20909
rect 16757 20904 22987 20906
rect 16757 20848 16762 20904
rect 16818 20848 18234 20904
rect 18290 20848 22926 20904
rect 22982 20848 22987 20904
rect 16757 20846 22987 20848
rect 16757 20843 16823 20846
rect 18229 20843 18295 20846
rect 22921 20843 22987 20846
rect 10174 20708 10180 20772
rect 10244 20770 10250 20772
rect 10501 20770 10567 20773
rect 10244 20768 10567 20770
rect 10244 20712 10506 20768
rect 10562 20712 10567 20768
rect 10244 20710 10567 20712
rect 10244 20708 10250 20710
rect 10501 20707 10567 20710
rect 16941 20770 17007 20773
rect 17166 20770 17172 20772
rect 16941 20768 17172 20770
rect 16941 20712 16946 20768
rect 17002 20712 17172 20768
rect 16941 20710 17172 20712
rect 16941 20707 17007 20710
rect 17166 20708 17172 20710
rect 17236 20770 17242 20772
rect 17677 20770 17743 20773
rect 17236 20768 17743 20770
rect 17236 20712 17682 20768
rect 17738 20712 17743 20768
rect 17236 20710 17743 20712
rect 17236 20708 17242 20710
rect 17677 20707 17743 20710
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 11432 20704 11748 20705
rect 11432 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11748 20704
rect 11432 20639 11748 20640
rect 19206 20704 19522 20705
rect 19206 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19522 20704
rect 19206 20639 19522 20640
rect 26980 20704 27296 20705
rect 26980 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27296 20704
rect 26980 20639 27296 20640
rect 8569 20634 8635 20637
rect 8886 20634 8892 20636
rect 8569 20632 8892 20634
rect 8569 20576 8574 20632
rect 8630 20576 8892 20632
rect 8569 20574 8892 20576
rect 8569 20571 8635 20574
rect 8886 20572 8892 20574
rect 8956 20572 8962 20636
rect 12893 20634 12959 20637
rect 13302 20634 13308 20636
rect 12893 20632 13308 20634
rect 12893 20576 12898 20632
rect 12954 20576 13308 20632
rect 12893 20574 13308 20576
rect 12893 20571 12959 20574
rect 13302 20572 13308 20574
rect 13372 20572 13378 20636
rect 13813 20634 13879 20637
rect 14406 20634 14412 20636
rect 13813 20632 14412 20634
rect 13813 20576 13818 20632
rect 13874 20576 14412 20632
rect 13813 20574 14412 20576
rect 13813 20571 13879 20574
rect 14406 20572 14412 20574
rect 14476 20572 14482 20636
rect 18045 20498 18111 20501
rect 19057 20498 19123 20501
rect 18045 20496 19123 20498
rect 18045 20440 18050 20496
rect 18106 20440 19062 20496
rect 19118 20440 19123 20496
rect 18045 20438 19123 20440
rect 18045 20435 18111 20438
rect 19057 20435 19123 20438
rect 18321 20362 18387 20365
rect 18873 20362 18939 20365
rect 18321 20360 18939 20362
rect 18321 20304 18326 20360
rect 18382 20304 18878 20360
rect 18934 20304 18939 20360
rect 18321 20302 18939 20304
rect 18321 20299 18387 20302
rect 18873 20299 18939 20302
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 12092 20160 12408 20161
rect 12092 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12408 20160
rect 12092 20095 12408 20096
rect 19866 20160 20182 20161
rect 19866 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20182 20160
rect 19866 20095 20182 20096
rect 27640 20160 27956 20161
rect 27640 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27956 20160
rect 27640 20095 27956 20096
rect 20345 20090 20411 20093
rect 23105 20090 23171 20093
rect 20345 20088 23171 20090
rect 20345 20032 20350 20088
rect 20406 20032 23110 20088
rect 23166 20032 23171 20088
rect 20345 20030 23171 20032
rect 20345 20027 20411 20030
rect 23105 20027 23171 20030
rect 16297 19954 16363 19957
rect 16614 19954 16620 19956
rect 16297 19952 16620 19954
rect 16297 19896 16302 19952
rect 16358 19896 16620 19952
rect 16297 19894 16620 19896
rect 16297 19891 16363 19894
rect 16614 19892 16620 19894
rect 16684 19892 16690 19956
rect 17585 19954 17651 19957
rect 26509 19954 26575 19957
rect 27521 19954 27587 19957
rect 17585 19952 27587 19954
rect 17585 19896 17590 19952
rect 17646 19896 26514 19952
rect 26570 19896 27526 19952
rect 27582 19896 27587 19952
rect 17585 19894 27587 19896
rect 17585 19891 17651 19894
rect 26509 19891 26575 19894
rect 27521 19891 27587 19894
rect 18505 19818 18571 19821
rect 19057 19818 19123 19821
rect 18505 19816 19123 19818
rect 18505 19760 18510 19816
rect 18566 19760 19062 19816
rect 19118 19760 19123 19816
rect 18505 19758 19123 19760
rect 18505 19755 18571 19758
rect 19057 19755 19123 19758
rect 22093 19818 22159 19821
rect 22737 19818 22803 19821
rect 22093 19816 22803 19818
rect 22093 19760 22098 19816
rect 22154 19760 22742 19816
rect 22798 19760 22803 19816
rect 22093 19758 22803 19760
rect 22093 19755 22159 19758
rect 22737 19755 22803 19758
rect 22277 19682 22343 19685
rect 22921 19682 22987 19685
rect 22277 19680 22987 19682
rect 22277 19624 22282 19680
rect 22338 19624 22926 19680
rect 22982 19624 22987 19680
rect 22277 19622 22987 19624
rect 22277 19619 22343 19622
rect 22921 19619 22987 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 3658 19551 3974 19552
rect 11432 19616 11748 19617
rect 11432 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11748 19616
rect 11432 19551 11748 19552
rect 19206 19616 19522 19617
rect 19206 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19522 19616
rect 19206 19551 19522 19552
rect 26980 19616 27296 19617
rect 26980 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27296 19616
rect 26980 19551 27296 19552
rect 6361 19274 6427 19277
rect 6637 19274 6703 19277
rect 6361 19272 6703 19274
rect 6361 19216 6366 19272
rect 6422 19216 6642 19272
rect 6698 19216 6703 19272
rect 6361 19214 6703 19216
rect 6361 19211 6427 19214
rect 6637 19211 6703 19214
rect 16798 19212 16804 19276
rect 16868 19274 16874 19276
rect 16941 19274 17007 19277
rect 16868 19272 17007 19274
rect 16868 19216 16946 19272
rect 17002 19216 17007 19272
rect 16868 19214 17007 19216
rect 16868 19212 16874 19214
rect 16941 19211 17007 19214
rect 17125 19274 17191 19277
rect 19149 19274 19215 19277
rect 17125 19272 19215 19274
rect 17125 19216 17130 19272
rect 17186 19216 19154 19272
rect 19210 19216 19215 19272
rect 17125 19214 19215 19216
rect 17125 19211 17191 19214
rect 19149 19211 19215 19214
rect 15653 19138 15719 19141
rect 16665 19138 16731 19141
rect 17033 19138 17099 19141
rect 15653 19136 17099 19138
rect 15653 19080 15658 19136
rect 15714 19080 16670 19136
rect 16726 19080 17038 19136
rect 17094 19080 17099 19136
rect 15653 19078 17099 19080
rect 15653 19075 15719 19078
rect 16665 19075 16731 19078
rect 17033 19075 17099 19078
rect 20253 19138 20319 19141
rect 23013 19138 23079 19141
rect 20253 19136 23079 19138
rect 20253 19080 20258 19136
rect 20314 19080 23018 19136
rect 23074 19080 23079 19136
rect 20253 19078 23079 19080
rect 20253 19075 20319 19078
rect 23013 19075 23079 19078
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 12092 19072 12408 19073
rect 12092 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12408 19072
rect 12092 19007 12408 19008
rect 19866 19072 20182 19073
rect 19866 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20182 19072
rect 19866 19007 20182 19008
rect 27640 19072 27956 19073
rect 27640 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27956 19072
rect 27640 19007 27956 19008
rect 17033 19002 17099 19005
rect 18505 19002 18571 19005
rect 17033 19000 18571 19002
rect 17033 18944 17038 19000
rect 17094 18944 18510 19000
rect 18566 18944 18571 19000
rect 17033 18942 18571 18944
rect 17033 18939 17099 18942
rect 18505 18939 18571 18942
rect 3969 18866 4035 18869
rect 4245 18866 4311 18869
rect 3969 18864 4311 18866
rect 3969 18808 3974 18864
rect 4030 18808 4250 18864
rect 4306 18808 4311 18864
rect 3969 18806 4311 18808
rect 3969 18803 4035 18806
rect 4245 18803 4311 18806
rect 16062 18804 16068 18868
rect 16132 18866 16138 18868
rect 16941 18866 17007 18869
rect 16132 18864 17007 18866
rect 16132 18808 16946 18864
rect 17002 18808 17007 18864
rect 16132 18806 17007 18808
rect 16132 18804 16138 18806
rect 16941 18803 17007 18806
rect 21449 18866 21515 18869
rect 27521 18866 27587 18869
rect 30189 18866 30255 18869
rect 21449 18864 30255 18866
rect 21449 18808 21454 18864
rect 21510 18808 27526 18864
rect 27582 18808 30194 18864
rect 30250 18808 30255 18864
rect 21449 18806 30255 18808
rect 21449 18803 21515 18806
rect 27521 18803 27587 18806
rect 30189 18803 30255 18806
rect 11881 18730 11947 18733
rect 24669 18730 24735 18733
rect 11881 18728 24735 18730
rect 11881 18672 11886 18728
rect 11942 18672 24674 18728
rect 24730 18672 24735 18728
rect 11881 18670 24735 18672
rect 11881 18667 11947 18670
rect 24669 18667 24735 18670
rect 16297 18594 16363 18597
rect 17493 18594 17559 18597
rect 20253 18596 20319 18597
rect 20253 18594 20300 18596
rect 16297 18592 17559 18594
rect 16297 18536 16302 18592
rect 16358 18536 17498 18592
rect 17554 18536 17559 18592
rect 16297 18534 17559 18536
rect 20208 18592 20300 18594
rect 20208 18536 20258 18592
rect 20208 18534 20300 18536
rect 16297 18531 16363 18534
rect 17493 18531 17559 18534
rect 20253 18532 20300 18534
rect 20364 18532 20370 18596
rect 20478 18532 20484 18596
rect 20548 18594 20554 18596
rect 20713 18594 20779 18597
rect 20548 18592 20779 18594
rect 20548 18536 20718 18592
rect 20774 18536 20779 18592
rect 20548 18534 20779 18536
rect 20548 18532 20554 18534
rect 20253 18531 20319 18532
rect 20713 18531 20779 18534
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 11432 18528 11748 18529
rect 11432 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11748 18528
rect 11432 18463 11748 18464
rect 19206 18528 19522 18529
rect 19206 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19522 18528
rect 19206 18463 19522 18464
rect 26980 18528 27296 18529
rect 26980 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27296 18528
rect 26980 18463 27296 18464
rect 14917 18460 14983 18461
rect 14917 18458 14964 18460
rect 14836 18456 14964 18458
rect 15028 18458 15034 18460
rect 15285 18458 15351 18461
rect 17217 18458 17283 18461
rect 17493 18458 17559 18461
rect 15028 18456 17559 18458
rect 14836 18400 14922 18456
rect 15028 18400 15290 18456
rect 15346 18400 17222 18456
rect 17278 18400 17498 18456
rect 17554 18400 17559 18456
rect 14836 18398 14964 18400
rect 14917 18396 14964 18398
rect 15028 18398 17559 18400
rect 15028 18396 15034 18398
rect 14917 18395 14983 18396
rect 15285 18395 15351 18398
rect 17217 18395 17283 18398
rect 17493 18395 17559 18398
rect 20069 18458 20135 18461
rect 22921 18458 22987 18461
rect 20069 18456 22987 18458
rect 20069 18400 20074 18456
rect 20130 18400 22926 18456
rect 22982 18400 22987 18456
rect 20069 18398 22987 18400
rect 20069 18395 20135 18398
rect 22921 18395 22987 18398
rect 10501 18322 10567 18325
rect 22461 18322 22527 18325
rect 10501 18320 22527 18322
rect 10501 18264 10506 18320
rect 10562 18264 22466 18320
rect 22522 18264 22527 18320
rect 10501 18262 22527 18264
rect 10501 18259 10567 18262
rect 22461 18259 22527 18262
rect 10041 18186 10107 18189
rect 21909 18186 21975 18189
rect 25313 18186 25379 18189
rect 10041 18184 25379 18186
rect 10041 18128 10046 18184
rect 10102 18128 21914 18184
rect 21970 18128 25318 18184
rect 25374 18128 25379 18184
rect 10041 18126 25379 18128
rect 10041 18123 10107 18126
rect 21909 18123 21975 18126
rect 25313 18123 25379 18126
rect 16297 18050 16363 18053
rect 18229 18050 18295 18053
rect 20437 18052 20503 18053
rect 20437 18050 20484 18052
rect 16297 18048 18295 18050
rect 16297 17992 16302 18048
rect 16358 17992 18234 18048
rect 18290 17992 18295 18048
rect 16297 17990 18295 17992
rect 20392 18048 20484 18050
rect 20392 17992 20442 18048
rect 20392 17990 20484 17992
rect 16297 17987 16363 17990
rect 18229 17987 18295 17990
rect 20437 17988 20484 17990
rect 20548 17988 20554 18052
rect 22461 18050 22527 18053
rect 25865 18050 25931 18053
rect 22461 18048 25931 18050
rect 22461 17992 22466 18048
rect 22522 17992 25870 18048
rect 25926 17992 25931 18048
rect 22461 17990 25931 17992
rect 20437 17987 20503 17988
rect 22461 17987 22527 17990
rect 25865 17987 25931 17990
rect 28073 18050 28139 18053
rect 28758 18050 28764 18052
rect 28073 18048 28764 18050
rect 28073 17992 28078 18048
rect 28134 17992 28764 18048
rect 28073 17990 28764 17992
rect 28073 17987 28139 17990
rect 28758 17988 28764 17990
rect 28828 17988 28834 18052
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 12092 17984 12408 17985
rect 12092 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12408 17984
rect 12092 17919 12408 17920
rect 19866 17984 20182 17985
rect 19866 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20182 17984
rect 19866 17919 20182 17920
rect 27640 17984 27956 17985
rect 27640 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27956 17984
rect 27640 17919 27956 17920
rect 13261 17914 13327 17917
rect 17033 17914 17099 17917
rect 13261 17912 17099 17914
rect 13261 17856 13266 17912
rect 13322 17856 17038 17912
rect 17094 17856 17099 17912
rect 13261 17854 17099 17856
rect 13261 17851 13327 17854
rect 17033 17851 17099 17854
rect 10133 17778 10199 17781
rect 11973 17778 12039 17781
rect 10133 17776 12039 17778
rect 10133 17720 10138 17776
rect 10194 17720 11978 17776
rect 12034 17720 12039 17776
rect 10133 17718 12039 17720
rect 10133 17715 10199 17718
rect 11973 17715 12039 17718
rect 13813 17778 13879 17781
rect 15561 17778 15627 17781
rect 17125 17778 17191 17781
rect 13813 17776 17191 17778
rect 13813 17720 13818 17776
rect 13874 17720 15566 17776
rect 15622 17720 17130 17776
rect 17186 17720 17191 17776
rect 13813 17718 17191 17720
rect 13813 17715 13879 17718
rect 15561 17715 15627 17718
rect 17125 17715 17191 17718
rect 11789 17642 11855 17645
rect 21265 17642 21331 17645
rect 11789 17640 21331 17642
rect 11789 17584 11794 17640
rect 11850 17584 21270 17640
rect 21326 17584 21331 17640
rect 11789 17582 21331 17584
rect 11789 17579 11855 17582
rect 21265 17579 21331 17582
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 11432 17440 11748 17441
rect 11432 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11748 17440
rect 11432 17375 11748 17376
rect 19206 17440 19522 17441
rect 19206 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19522 17440
rect 19206 17375 19522 17376
rect 26980 17440 27296 17441
rect 26980 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27296 17440
rect 26980 17375 27296 17376
rect 16665 17370 16731 17373
rect 16798 17370 16804 17372
rect 16665 17368 16804 17370
rect 16665 17312 16670 17368
rect 16726 17312 16804 17368
rect 16665 17310 16804 17312
rect 16665 17307 16731 17310
rect 16798 17308 16804 17310
rect 16868 17308 16874 17372
rect 3417 17098 3483 17101
rect 9397 17098 9463 17101
rect 3417 17096 9463 17098
rect 3417 17040 3422 17096
rect 3478 17040 9402 17096
rect 9458 17040 9463 17096
rect 3417 17038 9463 17040
rect 3417 17035 3483 17038
rect 9397 17035 9463 17038
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 12092 16896 12408 16897
rect 12092 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12408 16896
rect 12092 16831 12408 16832
rect 19866 16896 20182 16897
rect 19866 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20182 16896
rect 19866 16831 20182 16832
rect 27640 16896 27956 16897
rect 27640 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27956 16896
rect 27640 16831 27956 16832
rect 20437 16826 20503 16829
rect 20713 16826 20779 16829
rect 20437 16824 20779 16826
rect 20437 16768 20442 16824
rect 20498 16768 20718 16824
rect 20774 16768 20779 16824
rect 20437 16766 20779 16768
rect 20437 16763 20503 16766
rect 20713 16763 20779 16766
rect 22461 16826 22527 16829
rect 26141 16826 26207 16829
rect 26601 16826 26667 16829
rect 22461 16824 26667 16826
rect 22461 16768 22466 16824
rect 22522 16768 26146 16824
rect 26202 16768 26606 16824
rect 26662 16768 26667 16824
rect 22461 16766 26667 16768
rect 22461 16763 22527 16766
rect 26141 16763 26207 16766
rect 26601 16763 26667 16766
rect 17861 16690 17927 16693
rect 20161 16690 20227 16693
rect 17861 16688 20227 16690
rect 17861 16632 17866 16688
rect 17922 16632 20166 16688
rect 20222 16632 20227 16688
rect 17861 16630 20227 16632
rect 17861 16627 17927 16630
rect 20161 16627 20227 16630
rect 20437 16690 20503 16693
rect 20621 16690 20687 16693
rect 24393 16690 24459 16693
rect 20437 16688 24459 16690
rect 20437 16632 20442 16688
rect 20498 16632 20626 16688
rect 20682 16632 24398 16688
rect 24454 16632 24459 16688
rect 20437 16630 24459 16632
rect 20437 16627 20503 16630
rect 20621 16627 20687 16630
rect 24393 16627 24459 16630
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 11432 16352 11748 16353
rect 11432 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11748 16352
rect 11432 16287 11748 16288
rect 19206 16352 19522 16353
rect 19206 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19522 16352
rect 19206 16287 19522 16288
rect 26980 16352 27296 16353
rect 26980 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27296 16352
rect 26980 16287 27296 16288
rect 22093 16146 22159 16149
rect 22737 16146 22803 16149
rect 22093 16144 22803 16146
rect 22093 16088 22098 16144
rect 22154 16088 22742 16144
rect 22798 16088 22803 16144
rect 22093 16086 22803 16088
rect 22093 16083 22159 16086
rect 22737 16083 22803 16086
rect 9489 16010 9555 16013
rect 10777 16010 10843 16013
rect 9489 16008 10843 16010
rect 9489 15952 9494 16008
rect 9550 15952 10782 16008
rect 10838 15952 10843 16008
rect 9489 15950 10843 15952
rect 9489 15947 9555 15950
rect 10777 15947 10843 15950
rect 20805 16010 20871 16013
rect 22921 16010 22987 16013
rect 20805 16008 22987 16010
rect 20805 15952 20810 16008
rect 20866 15952 22926 16008
rect 22982 15952 22987 16008
rect 20805 15950 22987 15952
rect 20805 15947 20871 15950
rect 22921 15947 22987 15950
rect 20253 15874 20319 15877
rect 21633 15874 21699 15877
rect 20253 15872 21699 15874
rect 20253 15816 20258 15872
rect 20314 15816 21638 15872
rect 21694 15816 21699 15872
rect 20253 15814 21699 15816
rect 20253 15811 20319 15814
rect 21633 15811 21699 15814
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 12092 15808 12408 15809
rect 12092 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12408 15808
rect 12092 15743 12408 15744
rect 19866 15808 20182 15809
rect 19866 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20182 15808
rect 19866 15743 20182 15744
rect 27640 15808 27956 15809
rect 27640 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27956 15808
rect 27640 15743 27956 15744
rect 20805 15738 20871 15741
rect 24577 15738 24643 15741
rect 20805 15736 24643 15738
rect 20805 15680 20810 15736
rect 20866 15680 24582 15736
rect 24638 15680 24643 15736
rect 20805 15678 24643 15680
rect 20805 15675 20871 15678
rect 24577 15675 24643 15678
rect 14181 15602 14247 15605
rect 21817 15602 21883 15605
rect 14181 15600 21883 15602
rect 14181 15544 14186 15600
rect 14242 15544 21822 15600
rect 21878 15544 21883 15600
rect 14181 15542 21883 15544
rect 14181 15539 14247 15542
rect 21817 15539 21883 15542
rect 3693 15466 3759 15469
rect 5257 15466 5323 15469
rect 3693 15464 5323 15466
rect 3693 15408 3698 15464
rect 3754 15408 5262 15464
rect 5318 15408 5323 15464
rect 3693 15406 5323 15408
rect 3693 15403 3759 15406
rect 5257 15403 5323 15406
rect 10225 15466 10291 15469
rect 20478 15466 20484 15468
rect 10225 15464 20484 15466
rect 10225 15408 10230 15464
rect 10286 15408 20484 15464
rect 10225 15406 20484 15408
rect 10225 15403 10291 15406
rect 20478 15404 20484 15406
rect 20548 15466 20554 15468
rect 21081 15466 21147 15469
rect 20548 15464 21147 15466
rect 20548 15408 21086 15464
rect 21142 15408 21147 15464
rect 20548 15406 21147 15408
rect 20548 15404 20554 15406
rect 21081 15403 21147 15406
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 11432 15264 11748 15265
rect 11432 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11748 15264
rect 11432 15199 11748 15200
rect 19206 15264 19522 15265
rect 19206 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19522 15264
rect 19206 15199 19522 15200
rect 26980 15264 27296 15265
rect 26980 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27296 15264
rect 26980 15199 27296 15200
rect 1945 15058 2011 15061
rect 7373 15058 7439 15061
rect 1945 15056 7439 15058
rect 1945 15000 1950 15056
rect 2006 15000 7378 15056
rect 7434 15000 7439 15056
rect 1945 14998 7439 15000
rect 1945 14995 2011 14998
rect 7373 14995 7439 14998
rect 17585 15058 17651 15061
rect 20897 15058 20963 15061
rect 17585 15056 20963 15058
rect 17585 15000 17590 15056
rect 17646 15000 20902 15056
rect 20958 15000 20963 15056
rect 17585 14998 20963 15000
rect 17585 14995 17651 14998
rect 20897 14995 20963 14998
rect 11237 14922 11303 14925
rect 12617 14922 12683 14925
rect 21173 14922 21239 14925
rect 11237 14920 21239 14922
rect 11237 14864 11242 14920
rect 11298 14864 12622 14920
rect 12678 14864 21178 14920
rect 21234 14864 21239 14920
rect 11237 14862 21239 14864
rect 11237 14859 11303 14862
rect 12617 14859 12683 14862
rect 21173 14859 21239 14862
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 12092 14720 12408 14721
rect 12092 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12408 14720
rect 12092 14655 12408 14656
rect 19866 14720 20182 14721
rect 19866 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20182 14720
rect 19866 14655 20182 14656
rect 27640 14720 27956 14721
rect 27640 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27956 14720
rect 27640 14655 27956 14656
rect 13261 14650 13327 14653
rect 18045 14650 18111 14653
rect 13261 14648 18111 14650
rect 13261 14592 13266 14648
rect 13322 14592 18050 14648
rect 18106 14592 18111 14648
rect 13261 14590 18111 14592
rect 13261 14587 13327 14590
rect 18045 14587 18111 14590
rect 4889 14514 4955 14517
rect 16205 14514 16271 14517
rect 4889 14512 16271 14514
rect 4889 14456 4894 14512
rect 4950 14456 16210 14512
rect 16266 14456 16271 14512
rect 4889 14454 16271 14456
rect 4889 14451 4955 14454
rect 16205 14451 16271 14454
rect 22645 14514 22711 14517
rect 28257 14514 28323 14517
rect 22645 14512 28323 14514
rect 22645 14456 22650 14512
rect 22706 14456 28262 14512
rect 28318 14456 28323 14512
rect 22645 14454 28323 14456
rect 22645 14451 22711 14454
rect 28257 14451 28323 14454
rect 24393 14378 24459 14381
rect 26233 14378 26299 14381
rect 26969 14378 27035 14381
rect 28349 14378 28415 14381
rect 24393 14376 28415 14378
rect 24393 14320 24398 14376
rect 24454 14320 26238 14376
rect 26294 14320 26974 14376
rect 27030 14320 28354 14376
rect 28410 14320 28415 14376
rect 24393 14318 28415 14320
rect 24393 14315 24459 14318
rect 26233 14315 26299 14318
rect 26969 14315 27035 14318
rect 28349 14315 28415 14318
rect 19885 14242 19951 14245
rect 21725 14242 21791 14245
rect 22093 14242 22159 14245
rect 19885 14240 22159 14242
rect 19885 14184 19890 14240
rect 19946 14184 21730 14240
rect 21786 14184 22098 14240
rect 22154 14184 22159 14240
rect 19885 14182 22159 14184
rect 19885 14179 19951 14182
rect 21725 14179 21791 14182
rect 22093 14179 22159 14182
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 11432 14176 11748 14177
rect 11432 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11748 14176
rect 11432 14111 11748 14112
rect 19206 14176 19522 14177
rect 19206 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19522 14176
rect 19206 14111 19522 14112
rect 26980 14176 27296 14177
rect 26980 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27296 14176
rect 26980 14111 27296 14112
rect 22553 13970 22619 13973
rect 28257 13970 28323 13973
rect 30189 13970 30255 13973
rect 22553 13968 30255 13970
rect 22553 13912 22558 13968
rect 22614 13912 28262 13968
rect 28318 13912 30194 13968
rect 30250 13912 30255 13968
rect 22553 13910 30255 13912
rect 22553 13907 22619 13910
rect 28257 13907 28323 13910
rect 30189 13907 30255 13910
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 12092 13632 12408 13633
rect 12092 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12408 13632
rect 12092 13567 12408 13568
rect 19866 13632 20182 13633
rect 19866 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20182 13632
rect 19866 13567 20182 13568
rect 27640 13632 27956 13633
rect 27640 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27956 13632
rect 27640 13567 27956 13568
rect 19977 13426 20043 13429
rect 20294 13426 20300 13428
rect 19977 13424 20300 13426
rect 19977 13368 19982 13424
rect 20038 13368 20300 13424
rect 19977 13366 20300 13368
rect 19977 13363 20043 13366
rect 20294 13364 20300 13366
rect 20364 13364 20370 13428
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 11432 13088 11748 13089
rect 11432 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11748 13088
rect 11432 13023 11748 13024
rect 19206 13088 19522 13089
rect 19206 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19522 13088
rect 19206 13023 19522 13024
rect 26980 13088 27296 13089
rect 26980 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27296 13088
rect 26980 13023 27296 13024
rect 10593 12882 10659 12885
rect 15929 12882 15995 12885
rect 16297 12882 16363 12885
rect 16481 12882 16547 12885
rect 10593 12880 16547 12882
rect 10593 12824 10598 12880
rect 10654 12824 15934 12880
rect 15990 12824 16302 12880
rect 16358 12824 16486 12880
rect 16542 12824 16547 12880
rect 10593 12822 16547 12824
rect 10593 12819 10659 12822
rect 15929 12819 15995 12822
rect 16297 12819 16363 12822
rect 16481 12819 16547 12822
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 12092 12544 12408 12545
rect 12092 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12408 12544
rect 12092 12479 12408 12480
rect 19866 12544 20182 12545
rect 19866 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20182 12544
rect 19866 12479 20182 12480
rect 27640 12544 27956 12545
rect 27640 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27956 12544
rect 27640 12479 27956 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 11432 12000 11748 12001
rect 11432 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11748 12000
rect 11432 11935 11748 11936
rect 19206 12000 19522 12001
rect 19206 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19522 12000
rect 19206 11935 19522 11936
rect 26980 12000 27296 12001
rect 26980 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27296 12000
rect 26980 11935 27296 11936
rect 10041 11930 10107 11933
rect 10174 11930 10180 11932
rect 10041 11928 10180 11930
rect 10041 11872 10046 11928
rect 10102 11872 10180 11928
rect 10041 11870 10180 11872
rect 10041 11867 10107 11870
rect 10174 11868 10180 11870
rect 10244 11868 10250 11932
rect 3785 11794 3851 11797
rect 4429 11794 4495 11797
rect 3785 11792 4495 11794
rect 3785 11736 3790 11792
rect 3846 11736 4434 11792
rect 4490 11736 4495 11792
rect 3785 11734 4495 11736
rect 3785 11731 3851 11734
rect 4429 11731 4495 11734
rect 4061 11658 4127 11661
rect 8109 11658 8175 11661
rect 4061 11656 8175 11658
rect 4061 11600 4066 11656
rect 4122 11600 8114 11656
rect 8170 11600 8175 11656
rect 4061 11598 8175 11600
rect 4061 11595 4127 11598
rect 8109 11595 8175 11598
rect 11973 11658 12039 11661
rect 27061 11658 27127 11661
rect 11973 11656 27127 11658
rect 11973 11600 11978 11656
rect 12034 11600 27066 11656
rect 27122 11600 27127 11656
rect 11973 11598 27127 11600
rect 11973 11595 12039 11598
rect 27061 11595 27127 11598
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 12092 11456 12408 11457
rect 12092 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12408 11456
rect 12092 11391 12408 11392
rect 19866 11456 20182 11457
rect 19866 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20182 11456
rect 19866 11391 20182 11392
rect 27640 11456 27956 11457
rect 27640 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27956 11456
rect 27640 11391 27956 11392
rect 14089 11386 14155 11389
rect 17677 11386 17743 11389
rect 14089 11384 17743 11386
rect 14089 11328 14094 11384
rect 14150 11328 17682 11384
rect 17738 11328 17743 11384
rect 14089 11326 17743 11328
rect 14089 11323 14155 11326
rect 17677 11323 17743 11326
rect 5257 11250 5323 11253
rect 17769 11250 17835 11253
rect 5257 11248 17835 11250
rect 5257 11192 5262 11248
rect 5318 11192 17774 11248
rect 17830 11192 17835 11248
rect 5257 11190 17835 11192
rect 5257 11187 5323 11190
rect 17769 11187 17835 11190
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 11432 10912 11748 10913
rect 11432 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11748 10912
rect 11432 10847 11748 10848
rect 19206 10912 19522 10913
rect 19206 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19522 10912
rect 19206 10847 19522 10848
rect 26980 10912 27296 10913
rect 26980 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27296 10912
rect 26980 10847 27296 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 12092 10368 12408 10369
rect 12092 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12408 10368
rect 12092 10303 12408 10304
rect 19866 10368 20182 10369
rect 19866 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20182 10368
rect 19866 10303 20182 10304
rect 27640 10368 27956 10369
rect 27640 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27956 10368
rect 27640 10303 27956 10304
rect 6545 10162 6611 10165
rect 8569 10162 8635 10165
rect 6545 10160 8635 10162
rect 6545 10104 6550 10160
rect 6606 10104 8574 10160
rect 8630 10104 8635 10160
rect 6545 10102 8635 10104
rect 6545 10099 6611 10102
rect 8569 10099 8635 10102
rect 12065 10162 12131 10165
rect 16297 10162 16363 10165
rect 12065 10160 16363 10162
rect 12065 10104 12070 10160
rect 12126 10104 16302 10160
rect 16358 10104 16363 10160
rect 12065 10102 16363 10104
rect 12065 10099 12131 10102
rect 16297 10099 16363 10102
rect 3785 10026 3851 10029
rect 3558 10024 3851 10026
rect 3558 9992 3790 10024
rect 3512 9968 3790 9992
rect 3846 9968 3851 10024
rect 3512 9966 3851 9968
rect 3512 9932 3618 9966
rect 3785 9963 3851 9966
rect 4061 10026 4127 10029
rect 12341 10026 12407 10029
rect 16021 10026 16087 10029
rect 4061 10024 4170 10026
rect 4061 9968 4066 10024
rect 4122 9968 4170 10024
rect 4061 9963 4170 9968
rect 12341 10024 16087 10026
rect 12341 9968 12346 10024
rect 12402 9968 16026 10024
rect 16082 9968 16087 10024
rect 12341 9966 16087 9968
rect 12341 9963 12407 9966
rect 16021 9963 16087 9966
rect 3233 9890 3299 9893
rect 3512 9890 3572 9932
rect 3190 9888 3299 9890
rect 3190 9832 3238 9888
rect 3294 9832 3299 9888
rect 3190 9827 3299 9832
rect 3420 9830 3572 9890
rect 3190 9757 3250 9827
rect 3190 9752 3299 9757
rect 3190 9696 3238 9752
rect 3294 9696 3299 9752
rect 3190 9694 3299 9696
rect 3233 9691 3299 9694
rect 3420 9618 3480 9830
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 4110 9693 4170 9963
rect 11432 9824 11748 9825
rect 11432 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11748 9824
rect 11432 9759 11748 9760
rect 19206 9824 19522 9825
rect 19206 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19522 9824
rect 19206 9759 19522 9760
rect 26980 9824 27296 9825
rect 26980 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27296 9824
rect 26980 9759 27296 9760
rect 4061 9688 4170 9693
rect 4061 9632 4066 9688
rect 4122 9632 4170 9688
rect 4061 9630 4170 9632
rect 4061 9627 4127 9630
rect 3601 9618 3667 9621
rect 3420 9616 3667 9618
rect 3420 9560 3606 9616
rect 3662 9560 3667 9616
rect 3420 9558 3667 9560
rect 3601 9555 3667 9558
rect 3141 9482 3207 9485
rect 3969 9482 4035 9485
rect 3141 9480 4035 9482
rect 3141 9424 3146 9480
rect 3202 9424 3974 9480
rect 4030 9424 4035 9480
rect 3141 9422 4035 9424
rect 3141 9419 3207 9422
rect 3969 9419 4035 9422
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 12092 9280 12408 9281
rect 12092 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12408 9280
rect 12092 9215 12408 9216
rect 19866 9280 20182 9281
rect 19866 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20182 9280
rect 19866 9215 20182 9216
rect 27640 9280 27956 9281
rect 27640 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27956 9280
rect 27640 9215 27956 9216
rect 3693 9074 3759 9077
rect 7281 9074 7347 9077
rect 3693 9072 7347 9074
rect 3693 9016 3698 9072
rect 3754 9016 7286 9072
rect 7342 9016 7347 9072
rect 3693 9014 7347 9016
rect 3693 9011 3759 9014
rect 7281 9011 7347 9014
rect 11881 9074 11947 9077
rect 12801 9074 12867 9077
rect 15561 9074 15627 9077
rect 11881 9072 15627 9074
rect 11881 9016 11886 9072
rect 11942 9016 12806 9072
rect 12862 9016 15566 9072
rect 15622 9016 15627 9072
rect 11881 9014 15627 9016
rect 11881 9011 11947 9014
rect 12801 9011 12867 9014
rect 15561 9011 15627 9014
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 11432 8736 11748 8737
rect 11432 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11748 8736
rect 11432 8671 11748 8672
rect 19206 8736 19522 8737
rect 19206 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19522 8736
rect 19206 8671 19522 8672
rect 26980 8736 27296 8737
rect 26980 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27296 8736
rect 26980 8671 27296 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 12092 8192 12408 8193
rect 12092 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12408 8192
rect 12092 8127 12408 8128
rect 19866 8192 20182 8193
rect 19866 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20182 8192
rect 19866 8127 20182 8128
rect 27640 8192 27956 8193
rect 27640 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27956 8192
rect 27640 8127 27956 8128
rect 3049 7986 3115 7989
rect 7373 7986 7439 7989
rect 3049 7984 7439 7986
rect 3049 7928 3054 7984
rect 3110 7928 7378 7984
rect 7434 7928 7439 7984
rect 3049 7926 7439 7928
rect 3049 7923 3115 7926
rect 7373 7923 7439 7926
rect 9857 7986 9923 7989
rect 10133 7986 10199 7989
rect 10593 7986 10659 7989
rect 9857 7984 10659 7986
rect 9857 7928 9862 7984
rect 9918 7928 10138 7984
rect 10194 7928 10598 7984
rect 10654 7928 10659 7984
rect 9857 7926 10659 7928
rect 9857 7923 9923 7926
rect 10133 7923 10199 7926
rect 10593 7923 10659 7926
rect 10317 7850 10383 7853
rect 15561 7850 15627 7853
rect 10317 7848 15627 7850
rect 10317 7792 10322 7848
rect 10378 7792 15566 7848
rect 15622 7792 15627 7848
rect 10317 7790 15627 7792
rect 10317 7787 10383 7790
rect 15561 7787 15627 7790
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 11432 7648 11748 7649
rect 11432 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11748 7648
rect 11432 7583 11748 7584
rect 19206 7648 19522 7649
rect 19206 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19522 7648
rect 19206 7583 19522 7584
rect 26980 7648 27296 7649
rect 26980 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27296 7648
rect 26980 7583 27296 7584
rect 14917 7578 14983 7581
rect 16297 7578 16363 7581
rect 14917 7576 16363 7578
rect 14917 7520 14922 7576
rect 14978 7520 16302 7576
rect 16358 7520 16363 7576
rect 14917 7518 16363 7520
rect 14917 7515 14983 7518
rect 16297 7515 16363 7518
rect 4429 7442 4495 7445
rect 15009 7442 15075 7445
rect 4429 7440 15075 7442
rect 4429 7384 4434 7440
rect 4490 7384 15014 7440
rect 15070 7384 15075 7440
rect 4429 7382 15075 7384
rect 4429 7379 4495 7382
rect 15009 7379 15075 7382
rect 3877 7306 3943 7309
rect 8385 7306 8451 7309
rect 3877 7304 8451 7306
rect 3877 7248 3882 7304
rect 3938 7248 8390 7304
rect 8446 7248 8451 7304
rect 3877 7246 8451 7248
rect 3877 7243 3943 7246
rect 8385 7243 8451 7246
rect 11789 7306 11855 7309
rect 16573 7306 16639 7309
rect 20621 7306 20687 7309
rect 11789 7304 20687 7306
rect 11789 7248 11794 7304
rect 11850 7248 16578 7304
rect 16634 7248 20626 7304
rect 20682 7248 20687 7304
rect 11789 7246 20687 7248
rect 11789 7243 11855 7246
rect 16573 7243 16639 7246
rect 20621 7243 20687 7246
rect 13077 7170 13143 7173
rect 15653 7170 15719 7173
rect 13077 7168 15719 7170
rect 13077 7112 13082 7168
rect 13138 7112 15658 7168
rect 15714 7112 15719 7168
rect 13077 7110 15719 7112
rect 13077 7107 13143 7110
rect 15653 7107 15719 7110
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 12092 7104 12408 7105
rect 12092 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12408 7104
rect 12092 7039 12408 7040
rect 19866 7104 20182 7105
rect 19866 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20182 7104
rect 19866 7039 20182 7040
rect 27640 7104 27956 7105
rect 27640 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27956 7104
rect 27640 7039 27956 7040
rect 6085 6626 6151 6629
rect 7465 6626 7531 6629
rect 6085 6624 7531 6626
rect 6085 6568 6090 6624
rect 6146 6568 7470 6624
rect 7526 6568 7531 6624
rect 6085 6566 7531 6568
rect 6085 6563 6151 6566
rect 7465 6563 7531 6566
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 11432 6560 11748 6561
rect 11432 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11748 6560
rect 11432 6495 11748 6496
rect 19206 6560 19522 6561
rect 19206 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19522 6560
rect 19206 6495 19522 6496
rect 26980 6560 27296 6561
rect 26980 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27296 6560
rect 26980 6495 27296 6496
rect 2497 6490 2563 6493
rect 3509 6490 3575 6493
rect 2497 6488 3575 6490
rect 2497 6432 2502 6488
rect 2558 6432 3514 6488
rect 3570 6432 3575 6488
rect 2497 6430 3575 6432
rect 2497 6427 2563 6430
rect 3509 6427 3575 6430
rect 6269 6490 6335 6493
rect 6913 6490 6979 6493
rect 6269 6488 6979 6490
rect 6269 6432 6274 6488
rect 6330 6432 6918 6488
rect 6974 6432 6979 6488
rect 6269 6430 6979 6432
rect 6269 6427 6335 6430
rect 6913 6427 6979 6430
rect 2129 6354 2195 6357
rect 3233 6354 3299 6357
rect 2129 6352 3299 6354
rect 2129 6296 2134 6352
rect 2190 6296 3238 6352
rect 3294 6296 3299 6352
rect 2129 6294 3299 6296
rect 2129 6291 2195 6294
rect 3233 6291 3299 6294
rect 2589 6218 2655 6221
rect 3417 6218 3483 6221
rect 2589 6216 3483 6218
rect 2589 6160 2594 6216
rect 2650 6160 3422 6216
rect 3478 6160 3483 6216
rect 2589 6158 3483 6160
rect 2589 6155 2655 6158
rect 3417 6155 3483 6158
rect 6821 6218 6887 6221
rect 13077 6218 13143 6221
rect 6821 6216 13143 6218
rect 6821 6160 6826 6216
rect 6882 6160 13082 6216
rect 13138 6160 13143 6216
rect 6821 6158 13143 6160
rect 6821 6155 6887 6158
rect 13077 6155 13143 6158
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 12092 6016 12408 6017
rect 12092 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12408 6016
rect 12092 5951 12408 5952
rect 19866 6016 20182 6017
rect 19866 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20182 6016
rect 19866 5951 20182 5952
rect 27640 6016 27956 6017
rect 27640 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27956 6016
rect 27640 5951 27956 5952
rect 10961 5810 11027 5813
rect 12157 5810 12223 5813
rect 10961 5808 12223 5810
rect 10961 5752 10966 5808
rect 11022 5752 12162 5808
rect 12218 5752 12223 5808
rect 10961 5750 12223 5752
rect 10961 5747 11027 5750
rect 12157 5747 12223 5750
rect 13997 5810 14063 5813
rect 14181 5810 14247 5813
rect 15745 5810 15811 5813
rect 13997 5808 15811 5810
rect 13997 5752 14002 5808
rect 14058 5752 14186 5808
rect 14242 5752 15750 5808
rect 15806 5752 15811 5808
rect 13997 5750 15811 5752
rect 13997 5747 14063 5750
rect 14181 5747 14247 5750
rect 15745 5747 15811 5750
rect 12893 5674 12959 5677
rect 13537 5674 13603 5677
rect 14733 5674 14799 5677
rect 15193 5674 15259 5677
rect 12893 5672 15259 5674
rect 12893 5616 12898 5672
rect 12954 5616 13542 5672
rect 13598 5616 14738 5672
rect 14794 5616 15198 5672
rect 15254 5616 15259 5672
rect 12893 5614 15259 5616
rect 12893 5611 12959 5614
rect 13537 5611 13603 5614
rect 14733 5611 14799 5614
rect 15193 5611 15259 5614
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 11432 5472 11748 5473
rect 11432 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11748 5472
rect 11432 5407 11748 5408
rect 19206 5472 19522 5473
rect 19206 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19522 5472
rect 19206 5407 19522 5408
rect 26980 5472 27296 5473
rect 26980 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27296 5472
rect 26980 5407 27296 5408
rect 13813 5266 13879 5269
rect 16113 5266 16179 5269
rect 13813 5264 16179 5266
rect 13813 5208 13818 5264
rect 13874 5208 16118 5264
rect 16174 5208 16179 5264
rect 13813 5206 16179 5208
rect 13813 5203 13879 5206
rect 16113 5203 16179 5206
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 12092 4928 12408 4929
rect 12092 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12408 4928
rect 12092 4863 12408 4864
rect 19866 4928 20182 4929
rect 19866 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20182 4928
rect 19866 4863 20182 4864
rect 27640 4928 27956 4929
rect 27640 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27956 4928
rect 27640 4863 27956 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 11432 4384 11748 4385
rect 11432 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11748 4384
rect 11432 4319 11748 4320
rect 19206 4384 19522 4385
rect 19206 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19522 4384
rect 19206 4319 19522 4320
rect 26980 4384 27296 4385
rect 26980 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27296 4384
rect 26980 4319 27296 4320
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 12092 3840 12408 3841
rect 12092 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12408 3840
rect 12092 3775 12408 3776
rect 19866 3840 20182 3841
rect 19866 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20182 3840
rect 19866 3775 20182 3776
rect 27640 3840 27956 3841
rect 27640 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27956 3840
rect 27640 3775 27956 3776
rect 6177 3634 6243 3637
rect 8661 3634 8727 3637
rect 6177 3632 8727 3634
rect 6177 3576 6182 3632
rect 6238 3576 8666 3632
rect 8722 3576 8727 3632
rect 6177 3574 8727 3576
rect 6177 3571 6243 3574
rect 8661 3571 8727 3574
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 11432 3296 11748 3297
rect 11432 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11748 3296
rect 11432 3231 11748 3232
rect 19206 3296 19522 3297
rect 19206 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19522 3296
rect 19206 3231 19522 3232
rect 26980 3296 27296 3297
rect 26980 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27296 3296
rect 26980 3231 27296 3232
rect 26693 2954 26759 2957
rect 28809 2954 28875 2957
rect 26693 2952 28875 2954
rect 26693 2896 26698 2952
rect 26754 2896 28814 2952
rect 28870 2896 28875 2952
rect 26693 2894 28875 2896
rect 26693 2891 26759 2894
rect 28809 2891 28875 2894
rect 10685 2818 10751 2821
rect 11513 2818 11579 2821
rect 11881 2818 11947 2821
rect 10685 2816 11947 2818
rect 10685 2760 10690 2816
rect 10746 2760 11518 2816
rect 11574 2760 11886 2816
rect 11942 2760 11947 2816
rect 10685 2758 11947 2760
rect 10685 2755 10751 2758
rect 11513 2755 11579 2758
rect 11881 2755 11947 2758
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 12092 2752 12408 2753
rect 12092 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12408 2752
rect 12092 2687 12408 2688
rect 19866 2752 20182 2753
rect 19866 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20182 2752
rect 19866 2687 20182 2688
rect 27640 2752 27956 2753
rect 27640 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27956 2752
rect 27640 2687 27956 2688
rect 11697 2410 11763 2413
rect 15009 2410 15075 2413
rect 11697 2408 15075 2410
rect 11697 2352 11702 2408
rect 11758 2352 15014 2408
rect 15070 2352 15075 2408
rect 11697 2350 15075 2352
rect 11697 2347 11763 2350
rect 15009 2347 15075 2350
rect 21449 2410 21515 2413
rect 22093 2410 22159 2413
rect 21449 2408 22159 2410
rect 21449 2352 21454 2408
rect 21510 2352 22098 2408
rect 22154 2352 22159 2408
rect 21449 2350 22159 2352
rect 21449 2347 21515 2350
rect 22093 2347 22159 2350
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 11432 2208 11748 2209
rect 11432 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11748 2208
rect 11432 2143 11748 2144
rect 19206 2208 19522 2209
rect 19206 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19522 2208
rect 19206 2143 19522 2144
rect 26980 2208 27296 2209
rect 26980 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27296 2208
rect 26980 2143 27296 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 12092 1664 12408 1665
rect 12092 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12408 1664
rect 12092 1599 12408 1600
rect 19866 1664 20182 1665
rect 19866 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20182 1664
rect 19866 1599 20182 1600
rect 27640 1664 27956 1665
rect 27640 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27956 1664
rect 27640 1599 27956 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 11432 1120 11748 1121
rect 11432 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11748 1120
rect 11432 1055 11748 1056
rect 19206 1120 19522 1121
rect 19206 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19522 1120
rect 19206 1055 19522 1056
rect 26980 1120 27296 1121
rect 26980 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27296 1120
rect 26980 1055 27296 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 12092 576 12408 577
rect 12092 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12408 576
rect 12092 511 12408 512
rect 19866 576 20182 577
rect 19866 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20182 576
rect 19866 511 20182 512
rect 27640 576 27956 577
rect 27640 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27956 576
rect 27640 511 27956 512
<< via3 >>
rect 11652 21932 11716 21996
rect 12204 21992 12268 21996
rect 12204 21936 12254 21992
rect 12254 21936 12268 21992
rect 12204 21932 12268 21936
rect 23796 21992 23860 21996
rect 23796 21936 23846 21992
rect 23846 21936 23860 21992
rect 23796 21932 23860 21936
rect 24900 21992 24964 21996
rect 24900 21936 24950 21992
rect 24950 21936 24964 21992
rect 24900 21932 24964 21936
rect 25452 21992 25516 21996
rect 25452 21936 25502 21992
rect 25502 21936 25516 21992
rect 25452 21932 25516 21936
rect 26004 21992 26068 21996
rect 26004 21936 26054 21992
rect 26054 21936 26068 21992
rect 26004 21932 26068 21936
rect 27108 21932 27172 21996
rect 27660 21932 27724 21996
rect 7788 21796 7852 21860
rect 21588 21856 21652 21860
rect 21588 21800 21638 21856
rect 21638 21800 21652 21856
rect 21588 21796 21652 21800
rect 24348 21856 24412 21860
rect 24348 21800 24398 21856
rect 24398 21800 24412 21856
rect 24348 21796 24412 21800
rect 26556 21856 26620 21860
rect 26556 21800 26570 21856
rect 26570 21800 26620 21856
rect 26556 21796 26620 21800
rect 28212 21796 28276 21860
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 11438 21788 11502 21792
rect 11438 21732 11442 21788
rect 11442 21732 11498 21788
rect 11498 21732 11502 21788
rect 11438 21728 11502 21732
rect 11518 21788 11582 21792
rect 11518 21732 11522 21788
rect 11522 21732 11578 21788
rect 11578 21732 11582 21788
rect 11518 21728 11582 21732
rect 11598 21788 11662 21792
rect 11598 21732 11602 21788
rect 11602 21732 11658 21788
rect 11658 21732 11662 21788
rect 11598 21728 11662 21732
rect 11678 21788 11742 21792
rect 11678 21732 11682 21788
rect 11682 21732 11738 21788
rect 11738 21732 11742 21788
rect 11678 21728 11742 21732
rect 19212 21788 19276 21792
rect 19212 21732 19216 21788
rect 19216 21732 19272 21788
rect 19272 21732 19276 21788
rect 19212 21728 19276 21732
rect 19292 21788 19356 21792
rect 19292 21732 19296 21788
rect 19296 21732 19352 21788
rect 19352 21732 19356 21788
rect 19292 21728 19356 21732
rect 19372 21788 19436 21792
rect 19372 21732 19376 21788
rect 19376 21732 19432 21788
rect 19432 21732 19436 21788
rect 19372 21728 19436 21732
rect 19452 21788 19516 21792
rect 19452 21732 19456 21788
rect 19456 21732 19512 21788
rect 19512 21732 19516 21788
rect 19452 21728 19516 21732
rect 26986 21788 27050 21792
rect 26986 21732 26990 21788
rect 26990 21732 27046 21788
rect 27046 21732 27050 21788
rect 26986 21728 27050 21732
rect 27066 21788 27130 21792
rect 27066 21732 27070 21788
rect 27070 21732 27126 21788
rect 27126 21732 27130 21788
rect 27066 21728 27130 21732
rect 27146 21788 27210 21792
rect 27146 21732 27150 21788
rect 27150 21732 27206 21788
rect 27206 21732 27210 21788
rect 27146 21728 27210 21732
rect 27226 21788 27290 21792
rect 27226 21732 27230 21788
rect 27230 21732 27286 21788
rect 27286 21732 27290 21788
rect 27226 21728 27290 21732
rect 6132 21660 6196 21724
rect 7236 21720 7300 21724
rect 7236 21664 7286 21720
rect 7286 21664 7300 21720
rect 7236 21660 7300 21664
rect 8340 21720 8404 21724
rect 8340 21664 8390 21720
rect 8390 21664 8404 21720
rect 8340 21660 8404 21664
rect 9996 21720 10060 21724
rect 9996 21664 10010 21720
rect 10010 21664 10060 21720
rect 9996 21660 10060 21664
rect 10548 21660 10612 21724
rect 12756 21720 12820 21724
rect 12756 21664 12806 21720
rect 12806 21664 12820 21720
rect 12756 21660 12820 21664
rect 11100 21524 11164 21588
rect 17724 21524 17788 21588
rect 18828 21524 18892 21588
rect 18276 21388 18340 21452
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 12098 21244 12162 21248
rect 12098 21188 12102 21244
rect 12102 21188 12158 21244
rect 12158 21188 12162 21244
rect 12098 21184 12162 21188
rect 12178 21244 12242 21248
rect 12178 21188 12182 21244
rect 12182 21188 12238 21244
rect 12238 21188 12242 21244
rect 12178 21184 12242 21188
rect 12258 21244 12322 21248
rect 12258 21188 12262 21244
rect 12262 21188 12318 21244
rect 12318 21188 12322 21244
rect 12258 21184 12322 21188
rect 12338 21244 12402 21248
rect 12338 21188 12342 21244
rect 12342 21188 12398 21244
rect 12398 21188 12402 21244
rect 12338 21184 12402 21188
rect 19872 21244 19936 21248
rect 19872 21188 19876 21244
rect 19876 21188 19932 21244
rect 19932 21188 19936 21244
rect 19872 21184 19936 21188
rect 19952 21244 20016 21248
rect 19952 21188 19956 21244
rect 19956 21188 20012 21244
rect 20012 21188 20016 21244
rect 19952 21184 20016 21188
rect 20032 21244 20096 21248
rect 20032 21188 20036 21244
rect 20036 21188 20092 21244
rect 20092 21188 20096 21244
rect 20032 21184 20096 21188
rect 20112 21244 20176 21248
rect 20112 21188 20116 21244
rect 20116 21188 20172 21244
rect 20172 21188 20176 21244
rect 20112 21184 20176 21188
rect 27646 21244 27710 21248
rect 27646 21188 27650 21244
rect 27650 21188 27706 21244
rect 27706 21188 27710 21244
rect 27646 21184 27710 21188
rect 27726 21244 27790 21248
rect 27726 21188 27730 21244
rect 27730 21188 27786 21244
rect 27786 21188 27790 21244
rect 27726 21184 27790 21188
rect 27806 21244 27870 21248
rect 27806 21188 27810 21244
rect 27810 21188 27866 21244
rect 27866 21188 27870 21244
rect 27806 21184 27870 21188
rect 27886 21244 27950 21248
rect 27886 21188 27890 21244
rect 27890 21188 27946 21244
rect 27946 21188 27950 21244
rect 27886 21184 27950 21188
rect 6684 21116 6748 21180
rect 9444 21116 9508 21180
rect 13860 21176 13924 21180
rect 13860 21120 13874 21176
rect 13874 21120 13924 21176
rect 13860 21116 13924 21120
rect 15516 21040 15580 21044
rect 15516 20984 15530 21040
rect 15530 20984 15580 21040
rect 15516 20980 15580 20984
rect 10180 20708 10244 20772
rect 17172 20708 17236 20772
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 11438 20700 11502 20704
rect 11438 20644 11442 20700
rect 11442 20644 11498 20700
rect 11498 20644 11502 20700
rect 11438 20640 11502 20644
rect 11518 20700 11582 20704
rect 11518 20644 11522 20700
rect 11522 20644 11578 20700
rect 11578 20644 11582 20700
rect 11518 20640 11582 20644
rect 11598 20700 11662 20704
rect 11598 20644 11602 20700
rect 11602 20644 11658 20700
rect 11658 20644 11662 20700
rect 11598 20640 11662 20644
rect 11678 20700 11742 20704
rect 11678 20644 11682 20700
rect 11682 20644 11738 20700
rect 11738 20644 11742 20700
rect 11678 20640 11742 20644
rect 19212 20700 19276 20704
rect 19212 20644 19216 20700
rect 19216 20644 19272 20700
rect 19272 20644 19276 20700
rect 19212 20640 19276 20644
rect 19292 20700 19356 20704
rect 19292 20644 19296 20700
rect 19296 20644 19352 20700
rect 19352 20644 19356 20700
rect 19292 20640 19356 20644
rect 19372 20700 19436 20704
rect 19372 20644 19376 20700
rect 19376 20644 19432 20700
rect 19432 20644 19436 20700
rect 19372 20640 19436 20644
rect 19452 20700 19516 20704
rect 19452 20644 19456 20700
rect 19456 20644 19512 20700
rect 19512 20644 19516 20700
rect 19452 20640 19516 20644
rect 26986 20700 27050 20704
rect 26986 20644 26990 20700
rect 26990 20644 27046 20700
rect 27046 20644 27050 20700
rect 26986 20640 27050 20644
rect 27066 20700 27130 20704
rect 27066 20644 27070 20700
rect 27070 20644 27126 20700
rect 27126 20644 27130 20700
rect 27066 20640 27130 20644
rect 27146 20700 27210 20704
rect 27146 20644 27150 20700
rect 27150 20644 27206 20700
rect 27206 20644 27210 20700
rect 27146 20640 27210 20644
rect 27226 20700 27290 20704
rect 27226 20644 27230 20700
rect 27230 20644 27286 20700
rect 27286 20644 27290 20700
rect 27226 20640 27290 20644
rect 8892 20572 8956 20636
rect 13308 20572 13372 20636
rect 14412 20572 14476 20636
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 12098 20156 12162 20160
rect 12098 20100 12102 20156
rect 12102 20100 12158 20156
rect 12158 20100 12162 20156
rect 12098 20096 12162 20100
rect 12178 20156 12242 20160
rect 12178 20100 12182 20156
rect 12182 20100 12238 20156
rect 12238 20100 12242 20156
rect 12178 20096 12242 20100
rect 12258 20156 12322 20160
rect 12258 20100 12262 20156
rect 12262 20100 12318 20156
rect 12318 20100 12322 20156
rect 12258 20096 12322 20100
rect 12338 20156 12402 20160
rect 12338 20100 12342 20156
rect 12342 20100 12398 20156
rect 12398 20100 12402 20156
rect 12338 20096 12402 20100
rect 19872 20156 19936 20160
rect 19872 20100 19876 20156
rect 19876 20100 19932 20156
rect 19932 20100 19936 20156
rect 19872 20096 19936 20100
rect 19952 20156 20016 20160
rect 19952 20100 19956 20156
rect 19956 20100 20012 20156
rect 20012 20100 20016 20156
rect 19952 20096 20016 20100
rect 20032 20156 20096 20160
rect 20032 20100 20036 20156
rect 20036 20100 20092 20156
rect 20092 20100 20096 20156
rect 20032 20096 20096 20100
rect 20112 20156 20176 20160
rect 20112 20100 20116 20156
rect 20116 20100 20172 20156
rect 20172 20100 20176 20156
rect 20112 20096 20176 20100
rect 27646 20156 27710 20160
rect 27646 20100 27650 20156
rect 27650 20100 27706 20156
rect 27706 20100 27710 20156
rect 27646 20096 27710 20100
rect 27726 20156 27790 20160
rect 27726 20100 27730 20156
rect 27730 20100 27786 20156
rect 27786 20100 27790 20156
rect 27726 20096 27790 20100
rect 27806 20156 27870 20160
rect 27806 20100 27810 20156
rect 27810 20100 27866 20156
rect 27866 20100 27870 20156
rect 27806 20096 27870 20100
rect 27886 20156 27950 20160
rect 27886 20100 27890 20156
rect 27890 20100 27946 20156
rect 27946 20100 27950 20156
rect 27886 20096 27950 20100
rect 16620 19892 16684 19956
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 11438 19612 11502 19616
rect 11438 19556 11442 19612
rect 11442 19556 11498 19612
rect 11498 19556 11502 19612
rect 11438 19552 11502 19556
rect 11518 19612 11582 19616
rect 11518 19556 11522 19612
rect 11522 19556 11578 19612
rect 11578 19556 11582 19612
rect 11518 19552 11582 19556
rect 11598 19612 11662 19616
rect 11598 19556 11602 19612
rect 11602 19556 11658 19612
rect 11658 19556 11662 19612
rect 11598 19552 11662 19556
rect 11678 19612 11742 19616
rect 11678 19556 11682 19612
rect 11682 19556 11738 19612
rect 11738 19556 11742 19612
rect 11678 19552 11742 19556
rect 19212 19612 19276 19616
rect 19212 19556 19216 19612
rect 19216 19556 19272 19612
rect 19272 19556 19276 19612
rect 19212 19552 19276 19556
rect 19292 19612 19356 19616
rect 19292 19556 19296 19612
rect 19296 19556 19352 19612
rect 19352 19556 19356 19612
rect 19292 19552 19356 19556
rect 19372 19612 19436 19616
rect 19372 19556 19376 19612
rect 19376 19556 19432 19612
rect 19432 19556 19436 19612
rect 19372 19552 19436 19556
rect 19452 19612 19516 19616
rect 19452 19556 19456 19612
rect 19456 19556 19512 19612
rect 19512 19556 19516 19612
rect 19452 19552 19516 19556
rect 26986 19612 27050 19616
rect 26986 19556 26990 19612
rect 26990 19556 27046 19612
rect 27046 19556 27050 19612
rect 26986 19552 27050 19556
rect 27066 19612 27130 19616
rect 27066 19556 27070 19612
rect 27070 19556 27126 19612
rect 27126 19556 27130 19612
rect 27066 19552 27130 19556
rect 27146 19612 27210 19616
rect 27146 19556 27150 19612
rect 27150 19556 27206 19612
rect 27206 19556 27210 19612
rect 27146 19552 27210 19556
rect 27226 19612 27290 19616
rect 27226 19556 27230 19612
rect 27230 19556 27286 19612
rect 27286 19556 27290 19612
rect 27226 19552 27290 19556
rect 16804 19212 16868 19276
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 12098 19068 12162 19072
rect 12098 19012 12102 19068
rect 12102 19012 12158 19068
rect 12158 19012 12162 19068
rect 12098 19008 12162 19012
rect 12178 19068 12242 19072
rect 12178 19012 12182 19068
rect 12182 19012 12238 19068
rect 12238 19012 12242 19068
rect 12178 19008 12242 19012
rect 12258 19068 12322 19072
rect 12258 19012 12262 19068
rect 12262 19012 12318 19068
rect 12318 19012 12322 19068
rect 12258 19008 12322 19012
rect 12338 19068 12402 19072
rect 12338 19012 12342 19068
rect 12342 19012 12398 19068
rect 12398 19012 12402 19068
rect 12338 19008 12402 19012
rect 19872 19068 19936 19072
rect 19872 19012 19876 19068
rect 19876 19012 19932 19068
rect 19932 19012 19936 19068
rect 19872 19008 19936 19012
rect 19952 19068 20016 19072
rect 19952 19012 19956 19068
rect 19956 19012 20012 19068
rect 20012 19012 20016 19068
rect 19952 19008 20016 19012
rect 20032 19068 20096 19072
rect 20032 19012 20036 19068
rect 20036 19012 20092 19068
rect 20092 19012 20096 19068
rect 20032 19008 20096 19012
rect 20112 19068 20176 19072
rect 20112 19012 20116 19068
rect 20116 19012 20172 19068
rect 20172 19012 20176 19068
rect 20112 19008 20176 19012
rect 27646 19068 27710 19072
rect 27646 19012 27650 19068
rect 27650 19012 27706 19068
rect 27706 19012 27710 19068
rect 27646 19008 27710 19012
rect 27726 19068 27790 19072
rect 27726 19012 27730 19068
rect 27730 19012 27786 19068
rect 27786 19012 27790 19068
rect 27726 19008 27790 19012
rect 27806 19068 27870 19072
rect 27806 19012 27810 19068
rect 27810 19012 27866 19068
rect 27866 19012 27870 19068
rect 27806 19008 27870 19012
rect 27886 19068 27950 19072
rect 27886 19012 27890 19068
rect 27890 19012 27946 19068
rect 27946 19012 27950 19068
rect 27886 19008 27950 19012
rect 16068 18804 16132 18868
rect 20300 18592 20364 18596
rect 20300 18536 20314 18592
rect 20314 18536 20364 18592
rect 20300 18532 20364 18536
rect 20484 18532 20548 18596
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 11438 18524 11502 18528
rect 11438 18468 11442 18524
rect 11442 18468 11498 18524
rect 11498 18468 11502 18524
rect 11438 18464 11502 18468
rect 11518 18524 11582 18528
rect 11518 18468 11522 18524
rect 11522 18468 11578 18524
rect 11578 18468 11582 18524
rect 11518 18464 11582 18468
rect 11598 18524 11662 18528
rect 11598 18468 11602 18524
rect 11602 18468 11658 18524
rect 11658 18468 11662 18524
rect 11598 18464 11662 18468
rect 11678 18524 11742 18528
rect 11678 18468 11682 18524
rect 11682 18468 11738 18524
rect 11738 18468 11742 18524
rect 11678 18464 11742 18468
rect 19212 18524 19276 18528
rect 19212 18468 19216 18524
rect 19216 18468 19272 18524
rect 19272 18468 19276 18524
rect 19212 18464 19276 18468
rect 19292 18524 19356 18528
rect 19292 18468 19296 18524
rect 19296 18468 19352 18524
rect 19352 18468 19356 18524
rect 19292 18464 19356 18468
rect 19372 18524 19436 18528
rect 19372 18468 19376 18524
rect 19376 18468 19432 18524
rect 19432 18468 19436 18524
rect 19372 18464 19436 18468
rect 19452 18524 19516 18528
rect 19452 18468 19456 18524
rect 19456 18468 19512 18524
rect 19512 18468 19516 18524
rect 19452 18464 19516 18468
rect 26986 18524 27050 18528
rect 26986 18468 26990 18524
rect 26990 18468 27046 18524
rect 27046 18468 27050 18524
rect 26986 18464 27050 18468
rect 27066 18524 27130 18528
rect 27066 18468 27070 18524
rect 27070 18468 27126 18524
rect 27126 18468 27130 18524
rect 27066 18464 27130 18468
rect 27146 18524 27210 18528
rect 27146 18468 27150 18524
rect 27150 18468 27206 18524
rect 27206 18468 27210 18524
rect 27146 18464 27210 18468
rect 27226 18524 27290 18528
rect 27226 18468 27230 18524
rect 27230 18468 27286 18524
rect 27286 18468 27290 18524
rect 27226 18464 27290 18468
rect 14964 18456 15028 18460
rect 14964 18400 14978 18456
rect 14978 18400 15028 18456
rect 14964 18396 15028 18400
rect 20484 18048 20548 18052
rect 20484 17992 20498 18048
rect 20498 17992 20548 18048
rect 20484 17988 20548 17992
rect 28764 17988 28828 18052
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 12098 17980 12162 17984
rect 12098 17924 12102 17980
rect 12102 17924 12158 17980
rect 12158 17924 12162 17980
rect 12098 17920 12162 17924
rect 12178 17980 12242 17984
rect 12178 17924 12182 17980
rect 12182 17924 12238 17980
rect 12238 17924 12242 17980
rect 12178 17920 12242 17924
rect 12258 17980 12322 17984
rect 12258 17924 12262 17980
rect 12262 17924 12318 17980
rect 12318 17924 12322 17980
rect 12258 17920 12322 17924
rect 12338 17980 12402 17984
rect 12338 17924 12342 17980
rect 12342 17924 12398 17980
rect 12398 17924 12402 17980
rect 12338 17920 12402 17924
rect 19872 17980 19936 17984
rect 19872 17924 19876 17980
rect 19876 17924 19932 17980
rect 19932 17924 19936 17980
rect 19872 17920 19936 17924
rect 19952 17980 20016 17984
rect 19952 17924 19956 17980
rect 19956 17924 20012 17980
rect 20012 17924 20016 17980
rect 19952 17920 20016 17924
rect 20032 17980 20096 17984
rect 20032 17924 20036 17980
rect 20036 17924 20092 17980
rect 20092 17924 20096 17980
rect 20032 17920 20096 17924
rect 20112 17980 20176 17984
rect 20112 17924 20116 17980
rect 20116 17924 20172 17980
rect 20172 17924 20176 17980
rect 20112 17920 20176 17924
rect 27646 17980 27710 17984
rect 27646 17924 27650 17980
rect 27650 17924 27706 17980
rect 27706 17924 27710 17980
rect 27646 17920 27710 17924
rect 27726 17980 27790 17984
rect 27726 17924 27730 17980
rect 27730 17924 27786 17980
rect 27786 17924 27790 17980
rect 27726 17920 27790 17924
rect 27806 17980 27870 17984
rect 27806 17924 27810 17980
rect 27810 17924 27866 17980
rect 27866 17924 27870 17980
rect 27806 17920 27870 17924
rect 27886 17980 27950 17984
rect 27886 17924 27890 17980
rect 27890 17924 27946 17980
rect 27946 17924 27950 17980
rect 27886 17920 27950 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 11438 17436 11502 17440
rect 11438 17380 11442 17436
rect 11442 17380 11498 17436
rect 11498 17380 11502 17436
rect 11438 17376 11502 17380
rect 11518 17436 11582 17440
rect 11518 17380 11522 17436
rect 11522 17380 11578 17436
rect 11578 17380 11582 17436
rect 11518 17376 11582 17380
rect 11598 17436 11662 17440
rect 11598 17380 11602 17436
rect 11602 17380 11658 17436
rect 11658 17380 11662 17436
rect 11598 17376 11662 17380
rect 11678 17436 11742 17440
rect 11678 17380 11682 17436
rect 11682 17380 11738 17436
rect 11738 17380 11742 17436
rect 11678 17376 11742 17380
rect 19212 17436 19276 17440
rect 19212 17380 19216 17436
rect 19216 17380 19272 17436
rect 19272 17380 19276 17436
rect 19212 17376 19276 17380
rect 19292 17436 19356 17440
rect 19292 17380 19296 17436
rect 19296 17380 19352 17436
rect 19352 17380 19356 17436
rect 19292 17376 19356 17380
rect 19372 17436 19436 17440
rect 19372 17380 19376 17436
rect 19376 17380 19432 17436
rect 19432 17380 19436 17436
rect 19372 17376 19436 17380
rect 19452 17436 19516 17440
rect 19452 17380 19456 17436
rect 19456 17380 19512 17436
rect 19512 17380 19516 17436
rect 19452 17376 19516 17380
rect 26986 17436 27050 17440
rect 26986 17380 26990 17436
rect 26990 17380 27046 17436
rect 27046 17380 27050 17436
rect 26986 17376 27050 17380
rect 27066 17436 27130 17440
rect 27066 17380 27070 17436
rect 27070 17380 27126 17436
rect 27126 17380 27130 17436
rect 27066 17376 27130 17380
rect 27146 17436 27210 17440
rect 27146 17380 27150 17436
rect 27150 17380 27206 17436
rect 27206 17380 27210 17436
rect 27146 17376 27210 17380
rect 27226 17436 27290 17440
rect 27226 17380 27230 17436
rect 27230 17380 27286 17436
rect 27286 17380 27290 17436
rect 27226 17376 27290 17380
rect 16804 17308 16868 17372
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 12098 16892 12162 16896
rect 12098 16836 12102 16892
rect 12102 16836 12158 16892
rect 12158 16836 12162 16892
rect 12098 16832 12162 16836
rect 12178 16892 12242 16896
rect 12178 16836 12182 16892
rect 12182 16836 12238 16892
rect 12238 16836 12242 16892
rect 12178 16832 12242 16836
rect 12258 16892 12322 16896
rect 12258 16836 12262 16892
rect 12262 16836 12318 16892
rect 12318 16836 12322 16892
rect 12258 16832 12322 16836
rect 12338 16892 12402 16896
rect 12338 16836 12342 16892
rect 12342 16836 12398 16892
rect 12398 16836 12402 16892
rect 12338 16832 12402 16836
rect 19872 16892 19936 16896
rect 19872 16836 19876 16892
rect 19876 16836 19932 16892
rect 19932 16836 19936 16892
rect 19872 16832 19936 16836
rect 19952 16892 20016 16896
rect 19952 16836 19956 16892
rect 19956 16836 20012 16892
rect 20012 16836 20016 16892
rect 19952 16832 20016 16836
rect 20032 16892 20096 16896
rect 20032 16836 20036 16892
rect 20036 16836 20092 16892
rect 20092 16836 20096 16892
rect 20032 16832 20096 16836
rect 20112 16892 20176 16896
rect 20112 16836 20116 16892
rect 20116 16836 20172 16892
rect 20172 16836 20176 16892
rect 20112 16832 20176 16836
rect 27646 16892 27710 16896
rect 27646 16836 27650 16892
rect 27650 16836 27706 16892
rect 27706 16836 27710 16892
rect 27646 16832 27710 16836
rect 27726 16892 27790 16896
rect 27726 16836 27730 16892
rect 27730 16836 27786 16892
rect 27786 16836 27790 16892
rect 27726 16832 27790 16836
rect 27806 16892 27870 16896
rect 27806 16836 27810 16892
rect 27810 16836 27866 16892
rect 27866 16836 27870 16892
rect 27806 16832 27870 16836
rect 27886 16892 27950 16896
rect 27886 16836 27890 16892
rect 27890 16836 27946 16892
rect 27946 16836 27950 16892
rect 27886 16832 27950 16836
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 11438 16348 11502 16352
rect 11438 16292 11442 16348
rect 11442 16292 11498 16348
rect 11498 16292 11502 16348
rect 11438 16288 11502 16292
rect 11518 16348 11582 16352
rect 11518 16292 11522 16348
rect 11522 16292 11578 16348
rect 11578 16292 11582 16348
rect 11518 16288 11582 16292
rect 11598 16348 11662 16352
rect 11598 16292 11602 16348
rect 11602 16292 11658 16348
rect 11658 16292 11662 16348
rect 11598 16288 11662 16292
rect 11678 16348 11742 16352
rect 11678 16292 11682 16348
rect 11682 16292 11738 16348
rect 11738 16292 11742 16348
rect 11678 16288 11742 16292
rect 19212 16348 19276 16352
rect 19212 16292 19216 16348
rect 19216 16292 19272 16348
rect 19272 16292 19276 16348
rect 19212 16288 19276 16292
rect 19292 16348 19356 16352
rect 19292 16292 19296 16348
rect 19296 16292 19352 16348
rect 19352 16292 19356 16348
rect 19292 16288 19356 16292
rect 19372 16348 19436 16352
rect 19372 16292 19376 16348
rect 19376 16292 19432 16348
rect 19432 16292 19436 16348
rect 19372 16288 19436 16292
rect 19452 16348 19516 16352
rect 19452 16292 19456 16348
rect 19456 16292 19512 16348
rect 19512 16292 19516 16348
rect 19452 16288 19516 16292
rect 26986 16348 27050 16352
rect 26986 16292 26990 16348
rect 26990 16292 27046 16348
rect 27046 16292 27050 16348
rect 26986 16288 27050 16292
rect 27066 16348 27130 16352
rect 27066 16292 27070 16348
rect 27070 16292 27126 16348
rect 27126 16292 27130 16348
rect 27066 16288 27130 16292
rect 27146 16348 27210 16352
rect 27146 16292 27150 16348
rect 27150 16292 27206 16348
rect 27206 16292 27210 16348
rect 27146 16288 27210 16292
rect 27226 16348 27290 16352
rect 27226 16292 27230 16348
rect 27230 16292 27286 16348
rect 27286 16292 27290 16348
rect 27226 16288 27290 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 12098 15804 12162 15808
rect 12098 15748 12102 15804
rect 12102 15748 12158 15804
rect 12158 15748 12162 15804
rect 12098 15744 12162 15748
rect 12178 15804 12242 15808
rect 12178 15748 12182 15804
rect 12182 15748 12238 15804
rect 12238 15748 12242 15804
rect 12178 15744 12242 15748
rect 12258 15804 12322 15808
rect 12258 15748 12262 15804
rect 12262 15748 12318 15804
rect 12318 15748 12322 15804
rect 12258 15744 12322 15748
rect 12338 15804 12402 15808
rect 12338 15748 12342 15804
rect 12342 15748 12398 15804
rect 12398 15748 12402 15804
rect 12338 15744 12402 15748
rect 19872 15804 19936 15808
rect 19872 15748 19876 15804
rect 19876 15748 19932 15804
rect 19932 15748 19936 15804
rect 19872 15744 19936 15748
rect 19952 15804 20016 15808
rect 19952 15748 19956 15804
rect 19956 15748 20012 15804
rect 20012 15748 20016 15804
rect 19952 15744 20016 15748
rect 20032 15804 20096 15808
rect 20032 15748 20036 15804
rect 20036 15748 20092 15804
rect 20092 15748 20096 15804
rect 20032 15744 20096 15748
rect 20112 15804 20176 15808
rect 20112 15748 20116 15804
rect 20116 15748 20172 15804
rect 20172 15748 20176 15804
rect 20112 15744 20176 15748
rect 27646 15804 27710 15808
rect 27646 15748 27650 15804
rect 27650 15748 27706 15804
rect 27706 15748 27710 15804
rect 27646 15744 27710 15748
rect 27726 15804 27790 15808
rect 27726 15748 27730 15804
rect 27730 15748 27786 15804
rect 27786 15748 27790 15804
rect 27726 15744 27790 15748
rect 27806 15804 27870 15808
rect 27806 15748 27810 15804
rect 27810 15748 27866 15804
rect 27866 15748 27870 15804
rect 27806 15744 27870 15748
rect 27886 15804 27950 15808
rect 27886 15748 27890 15804
rect 27890 15748 27946 15804
rect 27946 15748 27950 15804
rect 27886 15744 27950 15748
rect 20484 15404 20548 15468
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 11438 15260 11502 15264
rect 11438 15204 11442 15260
rect 11442 15204 11498 15260
rect 11498 15204 11502 15260
rect 11438 15200 11502 15204
rect 11518 15260 11582 15264
rect 11518 15204 11522 15260
rect 11522 15204 11578 15260
rect 11578 15204 11582 15260
rect 11518 15200 11582 15204
rect 11598 15260 11662 15264
rect 11598 15204 11602 15260
rect 11602 15204 11658 15260
rect 11658 15204 11662 15260
rect 11598 15200 11662 15204
rect 11678 15260 11742 15264
rect 11678 15204 11682 15260
rect 11682 15204 11738 15260
rect 11738 15204 11742 15260
rect 11678 15200 11742 15204
rect 19212 15260 19276 15264
rect 19212 15204 19216 15260
rect 19216 15204 19272 15260
rect 19272 15204 19276 15260
rect 19212 15200 19276 15204
rect 19292 15260 19356 15264
rect 19292 15204 19296 15260
rect 19296 15204 19352 15260
rect 19352 15204 19356 15260
rect 19292 15200 19356 15204
rect 19372 15260 19436 15264
rect 19372 15204 19376 15260
rect 19376 15204 19432 15260
rect 19432 15204 19436 15260
rect 19372 15200 19436 15204
rect 19452 15260 19516 15264
rect 19452 15204 19456 15260
rect 19456 15204 19512 15260
rect 19512 15204 19516 15260
rect 19452 15200 19516 15204
rect 26986 15260 27050 15264
rect 26986 15204 26990 15260
rect 26990 15204 27046 15260
rect 27046 15204 27050 15260
rect 26986 15200 27050 15204
rect 27066 15260 27130 15264
rect 27066 15204 27070 15260
rect 27070 15204 27126 15260
rect 27126 15204 27130 15260
rect 27066 15200 27130 15204
rect 27146 15260 27210 15264
rect 27146 15204 27150 15260
rect 27150 15204 27206 15260
rect 27206 15204 27210 15260
rect 27146 15200 27210 15204
rect 27226 15260 27290 15264
rect 27226 15204 27230 15260
rect 27230 15204 27286 15260
rect 27286 15204 27290 15260
rect 27226 15200 27290 15204
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 12098 14716 12162 14720
rect 12098 14660 12102 14716
rect 12102 14660 12158 14716
rect 12158 14660 12162 14716
rect 12098 14656 12162 14660
rect 12178 14716 12242 14720
rect 12178 14660 12182 14716
rect 12182 14660 12238 14716
rect 12238 14660 12242 14716
rect 12178 14656 12242 14660
rect 12258 14716 12322 14720
rect 12258 14660 12262 14716
rect 12262 14660 12318 14716
rect 12318 14660 12322 14716
rect 12258 14656 12322 14660
rect 12338 14716 12402 14720
rect 12338 14660 12342 14716
rect 12342 14660 12398 14716
rect 12398 14660 12402 14716
rect 12338 14656 12402 14660
rect 19872 14716 19936 14720
rect 19872 14660 19876 14716
rect 19876 14660 19932 14716
rect 19932 14660 19936 14716
rect 19872 14656 19936 14660
rect 19952 14716 20016 14720
rect 19952 14660 19956 14716
rect 19956 14660 20012 14716
rect 20012 14660 20016 14716
rect 19952 14656 20016 14660
rect 20032 14716 20096 14720
rect 20032 14660 20036 14716
rect 20036 14660 20092 14716
rect 20092 14660 20096 14716
rect 20032 14656 20096 14660
rect 20112 14716 20176 14720
rect 20112 14660 20116 14716
rect 20116 14660 20172 14716
rect 20172 14660 20176 14716
rect 20112 14656 20176 14660
rect 27646 14716 27710 14720
rect 27646 14660 27650 14716
rect 27650 14660 27706 14716
rect 27706 14660 27710 14716
rect 27646 14656 27710 14660
rect 27726 14716 27790 14720
rect 27726 14660 27730 14716
rect 27730 14660 27786 14716
rect 27786 14660 27790 14716
rect 27726 14656 27790 14660
rect 27806 14716 27870 14720
rect 27806 14660 27810 14716
rect 27810 14660 27866 14716
rect 27866 14660 27870 14716
rect 27806 14656 27870 14660
rect 27886 14716 27950 14720
rect 27886 14660 27890 14716
rect 27890 14660 27946 14716
rect 27946 14660 27950 14716
rect 27886 14656 27950 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 11438 14172 11502 14176
rect 11438 14116 11442 14172
rect 11442 14116 11498 14172
rect 11498 14116 11502 14172
rect 11438 14112 11502 14116
rect 11518 14172 11582 14176
rect 11518 14116 11522 14172
rect 11522 14116 11578 14172
rect 11578 14116 11582 14172
rect 11518 14112 11582 14116
rect 11598 14172 11662 14176
rect 11598 14116 11602 14172
rect 11602 14116 11658 14172
rect 11658 14116 11662 14172
rect 11598 14112 11662 14116
rect 11678 14172 11742 14176
rect 11678 14116 11682 14172
rect 11682 14116 11738 14172
rect 11738 14116 11742 14172
rect 11678 14112 11742 14116
rect 19212 14172 19276 14176
rect 19212 14116 19216 14172
rect 19216 14116 19272 14172
rect 19272 14116 19276 14172
rect 19212 14112 19276 14116
rect 19292 14172 19356 14176
rect 19292 14116 19296 14172
rect 19296 14116 19352 14172
rect 19352 14116 19356 14172
rect 19292 14112 19356 14116
rect 19372 14172 19436 14176
rect 19372 14116 19376 14172
rect 19376 14116 19432 14172
rect 19432 14116 19436 14172
rect 19372 14112 19436 14116
rect 19452 14172 19516 14176
rect 19452 14116 19456 14172
rect 19456 14116 19512 14172
rect 19512 14116 19516 14172
rect 19452 14112 19516 14116
rect 26986 14172 27050 14176
rect 26986 14116 26990 14172
rect 26990 14116 27046 14172
rect 27046 14116 27050 14172
rect 26986 14112 27050 14116
rect 27066 14172 27130 14176
rect 27066 14116 27070 14172
rect 27070 14116 27126 14172
rect 27126 14116 27130 14172
rect 27066 14112 27130 14116
rect 27146 14172 27210 14176
rect 27146 14116 27150 14172
rect 27150 14116 27206 14172
rect 27206 14116 27210 14172
rect 27146 14112 27210 14116
rect 27226 14172 27290 14176
rect 27226 14116 27230 14172
rect 27230 14116 27286 14172
rect 27286 14116 27290 14172
rect 27226 14112 27290 14116
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 12098 13628 12162 13632
rect 12098 13572 12102 13628
rect 12102 13572 12158 13628
rect 12158 13572 12162 13628
rect 12098 13568 12162 13572
rect 12178 13628 12242 13632
rect 12178 13572 12182 13628
rect 12182 13572 12238 13628
rect 12238 13572 12242 13628
rect 12178 13568 12242 13572
rect 12258 13628 12322 13632
rect 12258 13572 12262 13628
rect 12262 13572 12318 13628
rect 12318 13572 12322 13628
rect 12258 13568 12322 13572
rect 12338 13628 12402 13632
rect 12338 13572 12342 13628
rect 12342 13572 12398 13628
rect 12398 13572 12402 13628
rect 12338 13568 12402 13572
rect 19872 13628 19936 13632
rect 19872 13572 19876 13628
rect 19876 13572 19932 13628
rect 19932 13572 19936 13628
rect 19872 13568 19936 13572
rect 19952 13628 20016 13632
rect 19952 13572 19956 13628
rect 19956 13572 20012 13628
rect 20012 13572 20016 13628
rect 19952 13568 20016 13572
rect 20032 13628 20096 13632
rect 20032 13572 20036 13628
rect 20036 13572 20092 13628
rect 20092 13572 20096 13628
rect 20032 13568 20096 13572
rect 20112 13628 20176 13632
rect 20112 13572 20116 13628
rect 20116 13572 20172 13628
rect 20172 13572 20176 13628
rect 20112 13568 20176 13572
rect 27646 13628 27710 13632
rect 27646 13572 27650 13628
rect 27650 13572 27706 13628
rect 27706 13572 27710 13628
rect 27646 13568 27710 13572
rect 27726 13628 27790 13632
rect 27726 13572 27730 13628
rect 27730 13572 27786 13628
rect 27786 13572 27790 13628
rect 27726 13568 27790 13572
rect 27806 13628 27870 13632
rect 27806 13572 27810 13628
rect 27810 13572 27866 13628
rect 27866 13572 27870 13628
rect 27806 13568 27870 13572
rect 27886 13628 27950 13632
rect 27886 13572 27890 13628
rect 27890 13572 27946 13628
rect 27946 13572 27950 13628
rect 27886 13568 27950 13572
rect 20300 13364 20364 13428
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 11438 13084 11502 13088
rect 11438 13028 11442 13084
rect 11442 13028 11498 13084
rect 11498 13028 11502 13084
rect 11438 13024 11502 13028
rect 11518 13084 11582 13088
rect 11518 13028 11522 13084
rect 11522 13028 11578 13084
rect 11578 13028 11582 13084
rect 11518 13024 11582 13028
rect 11598 13084 11662 13088
rect 11598 13028 11602 13084
rect 11602 13028 11658 13084
rect 11658 13028 11662 13084
rect 11598 13024 11662 13028
rect 11678 13084 11742 13088
rect 11678 13028 11682 13084
rect 11682 13028 11738 13084
rect 11738 13028 11742 13084
rect 11678 13024 11742 13028
rect 19212 13084 19276 13088
rect 19212 13028 19216 13084
rect 19216 13028 19272 13084
rect 19272 13028 19276 13084
rect 19212 13024 19276 13028
rect 19292 13084 19356 13088
rect 19292 13028 19296 13084
rect 19296 13028 19352 13084
rect 19352 13028 19356 13084
rect 19292 13024 19356 13028
rect 19372 13084 19436 13088
rect 19372 13028 19376 13084
rect 19376 13028 19432 13084
rect 19432 13028 19436 13084
rect 19372 13024 19436 13028
rect 19452 13084 19516 13088
rect 19452 13028 19456 13084
rect 19456 13028 19512 13084
rect 19512 13028 19516 13084
rect 19452 13024 19516 13028
rect 26986 13084 27050 13088
rect 26986 13028 26990 13084
rect 26990 13028 27046 13084
rect 27046 13028 27050 13084
rect 26986 13024 27050 13028
rect 27066 13084 27130 13088
rect 27066 13028 27070 13084
rect 27070 13028 27126 13084
rect 27126 13028 27130 13084
rect 27066 13024 27130 13028
rect 27146 13084 27210 13088
rect 27146 13028 27150 13084
rect 27150 13028 27206 13084
rect 27206 13028 27210 13084
rect 27146 13024 27210 13028
rect 27226 13084 27290 13088
rect 27226 13028 27230 13084
rect 27230 13028 27286 13084
rect 27286 13028 27290 13084
rect 27226 13024 27290 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 12098 12540 12162 12544
rect 12098 12484 12102 12540
rect 12102 12484 12158 12540
rect 12158 12484 12162 12540
rect 12098 12480 12162 12484
rect 12178 12540 12242 12544
rect 12178 12484 12182 12540
rect 12182 12484 12238 12540
rect 12238 12484 12242 12540
rect 12178 12480 12242 12484
rect 12258 12540 12322 12544
rect 12258 12484 12262 12540
rect 12262 12484 12318 12540
rect 12318 12484 12322 12540
rect 12258 12480 12322 12484
rect 12338 12540 12402 12544
rect 12338 12484 12342 12540
rect 12342 12484 12398 12540
rect 12398 12484 12402 12540
rect 12338 12480 12402 12484
rect 19872 12540 19936 12544
rect 19872 12484 19876 12540
rect 19876 12484 19932 12540
rect 19932 12484 19936 12540
rect 19872 12480 19936 12484
rect 19952 12540 20016 12544
rect 19952 12484 19956 12540
rect 19956 12484 20012 12540
rect 20012 12484 20016 12540
rect 19952 12480 20016 12484
rect 20032 12540 20096 12544
rect 20032 12484 20036 12540
rect 20036 12484 20092 12540
rect 20092 12484 20096 12540
rect 20032 12480 20096 12484
rect 20112 12540 20176 12544
rect 20112 12484 20116 12540
rect 20116 12484 20172 12540
rect 20172 12484 20176 12540
rect 20112 12480 20176 12484
rect 27646 12540 27710 12544
rect 27646 12484 27650 12540
rect 27650 12484 27706 12540
rect 27706 12484 27710 12540
rect 27646 12480 27710 12484
rect 27726 12540 27790 12544
rect 27726 12484 27730 12540
rect 27730 12484 27786 12540
rect 27786 12484 27790 12540
rect 27726 12480 27790 12484
rect 27806 12540 27870 12544
rect 27806 12484 27810 12540
rect 27810 12484 27866 12540
rect 27866 12484 27870 12540
rect 27806 12480 27870 12484
rect 27886 12540 27950 12544
rect 27886 12484 27890 12540
rect 27890 12484 27946 12540
rect 27946 12484 27950 12540
rect 27886 12480 27950 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 11438 11996 11502 12000
rect 11438 11940 11442 11996
rect 11442 11940 11498 11996
rect 11498 11940 11502 11996
rect 11438 11936 11502 11940
rect 11518 11996 11582 12000
rect 11518 11940 11522 11996
rect 11522 11940 11578 11996
rect 11578 11940 11582 11996
rect 11518 11936 11582 11940
rect 11598 11996 11662 12000
rect 11598 11940 11602 11996
rect 11602 11940 11658 11996
rect 11658 11940 11662 11996
rect 11598 11936 11662 11940
rect 11678 11996 11742 12000
rect 11678 11940 11682 11996
rect 11682 11940 11738 11996
rect 11738 11940 11742 11996
rect 11678 11936 11742 11940
rect 19212 11996 19276 12000
rect 19212 11940 19216 11996
rect 19216 11940 19272 11996
rect 19272 11940 19276 11996
rect 19212 11936 19276 11940
rect 19292 11996 19356 12000
rect 19292 11940 19296 11996
rect 19296 11940 19352 11996
rect 19352 11940 19356 11996
rect 19292 11936 19356 11940
rect 19372 11996 19436 12000
rect 19372 11940 19376 11996
rect 19376 11940 19432 11996
rect 19432 11940 19436 11996
rect 19372 11936 19436 11940
rect 19452 11996 19516 12000
rect 19452 11940 19456 11996
rect 19456 11940 19512 11996
rect 19512 11940 19516 11996
rect 19452 11936 19516 11940
rect 26986 11996 27050 12000
rect 26986 11940 26990 11996
rect 26990 11940 27046 11996
rect 27046 11940 27050 11996
rect 26986 11936 27050 11940
rect 27066 11996 27130 12000
rect 27066 11940 27070 11996
rect 27070 11940 27126 11996
rect 27126 11940 27130 11996
rect 27066 11936 27130 11940
rect 27146 11996 27210 12000
rect 27146 11940 27150 11996
rect 27150 11940 27206 11996
rect 27206 11940 27210 11996
rect 27146 11936 27210 11940
rect 27226 11996 27290 12000
rect 27226 11940 27230 11996
rect 27230 11940 27286 11996
rect 27286 11940 27290 11996
rect 27226 11936 27290 11940
rect 10180 11868 10244 11932
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 12098 11452 12162 11456
rect 12098 11396 12102 11452
rect 12102 11396 12158 11452
rect 12158 11396 12162 11452
rect 12098 11392 12162 11396
rect 12178 11452 12242 11456
rect 12178 11396 12182 11452
rect 12182 11396 12238 11452
rect 12238 11396 12242 11452
rect 12178 11392 12242 11396
rect 12258 11452 12322 11456
rect 12258 11396 12262 11452
rect 12262 11396 12318 11452
rect 12318 11396 12322 11452
rect 12258 11392 12322 11396
rect 12338 11452 12402 11456
rect 12338 11396 12342 11452
rect 12342 11396 12398 11452
rect 12398 11396 12402 11452
rect 12338 11392 12402 11396
rect 19872 11452 19936 11456
rect 19872 11396 19876 11452
rect 19876 11396 19932 11452
rect 19932 11396 19936 11452
rect 19872 11392 19936 11396
rect 19952 11452 20016 11456
rect 19952 11396 19956 11452
rect 19956 11396 20012 11452
rect 20012 11396 20016 11452
rect 19952 11392 20016 11396
rect 20032 11452 20096 11456
rect 20032 11396 20036 11452
rect 20036 11396 20092 11452
rect 20092 11396 20096 11452
rect 20032 11392 20096 11396
rect 20112 11452 20176 11456
rect 20112 11396 20116 11452
rect 20116 11396 20172 11452
rect 20172 11396 20176 11452
rect 20112 11392 20176 11396
rect 27646 11452 27710 11456
rect 27646 11396 27650 11452
rect 27650 11396 27706 11452
rect 27706 11396 27710 11452
rect 27646 11392 27710 11396
rect 27726 11452 27790 11456
rect 27726 11396 27730 11452
rect 27730 11396 27786 11452
rect 27786 11396 27790 11452
rect 27726 11392 27790 11396
rect 27806 11452 27870 11456
rect 27806 11396 27810 11452
rect 27810 11396 27866 11452
rect 27866 11396 27870 11452
rect 27806 11392 27870 11396
rect 27886 11452 27950 11456
rect 27886 11396 27890 11452
rect 27890 11396 27946 11452
rect 27946 11396 27950 11452
rect 27886 11392 27950 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 11438 10908 11502 10912
rect 11438 10852 11442 10908
rect 11442 10852 11498 10908
rect 11498 10852 11502 10908
rect 11438 10848 11502 10852
rect 11518 10908 11582 10912
rect 11518 10852 11522 10908
rect 11522 10852 11578 10908
rect 11578 10852 11582 10908
rect 11518 10848 11582 10852
rect 11598 10908 11662 10912
rect 11598 10852 11602 10908
rect 11602 10852 11658 10908
rect 11658 10852 11662 10908
rect 11598 10848 11662 10852
rect 11678 10908 11742 10912
rect 11678 10852 11682 10908
rect 11682 10852 11738 10908
rect 11738 10852 11742 10908
rect 11678 10848 11742 10852
rect 19212 10908 19276 10912
rect 19212 10852 19216 10908
rect 19216 10852 19272 10908
rect 19272 10852 19276 10908
rect 19212 10848 19276 10852
rect 19292 10908 19356 10912
rect 19292 10852 19296 10908
rect 19296 10852 19352 10908
rect 19352 10852 19356 10908
rect 19292 10848 19356 10852
rect 19372 10908 19436 10912
rect 19372 10852 19376 10908
rect 19376 10852 19432 10908
rect 19432 10852 19436 10908
rect 19372 10848 19436 10852
rect 19452 10908 19516 10912
rect 19452 10852 19456 10908
rect 19456 10852 19512 10908
rect 19512 10852 19516 10908
rect 19452 10848 19516 10852
rect 26986 10908 27050 10912
rect 26986 10852 26990 10908
rect 26990 10852 27046 10908
rect 27046 10852 27050 10908
rect 26986 10848 27050 10852
rect 27066 10908 27130 10912
rect 27066 10852 27070 10908
rect 27070 10852 27126 10908
rect 27126 10852 27130 10908
rect 27066 10848 27130 10852
rect 27146 10908 27210 10912
rect 27146 10852 27150 10908
rect 27150 10852 27206 10908
rect 27206 10852 27210 10908
rect 27146 10848 27210 10852
rect 27226 10908 27290 10912
rect 27226 10852 27230 10908
rect 27230 10852 27286 10908
rect 27286 10852 27290 10908
rect 27226 10848 27290 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 12098 10364 12162 10368
rect 12098 10308 12102 10364
rect 12102 10308 12158 10364
rect 12158 10308 12162 10364
rect 12098 10304 12162 10308
rect 12178 10364 12242 10368
rect 12178 10308 12182 10364
rect 12182 10308 12238 10364
rect 12238 10308 12242 10364
rect 12178 10304 12242 10308
rect 12258 10364 12322 10368
rect 12258 10308 12262 10364
rect 12262 10308 12318 10364
rect 12318 10308 12322 10364
rect 12258 10304 12322 10308
rect 12338 10364 12402 10368
rect 12338 10308 12342 10364
rect 12342 10308 12398 10364
rect 12398 10308 12402 10364
rect 12338 10304 12402 10308
rect 19872 10364 19936 10368
rect 19872 10308 19876 10364
rect 19876 10308 19932 10364
rect 19932 10308 19936 10364
rect 19872 10304 19936 10308
rect 19952 10364 20016 10368
rect 19952 10308 19956 10364
rect 19956 10308 20012 10364
rect 20012 10308 20016 10364
rect 19952 10304 20016 10308
rect 20032 10364 20096 10368
rect 20032 10308 20036 10364
rect 20036 10308 20092 10364
rect 20092 10308 20096 10364
rect 20032 10304 20096 10308
rect 20112 10364 20176 10368
rect 20112 10308 20116 10364
rect 20116 10308 20172 10364
rect 20172 10308 20176 10364
rect 20112 10304 20176 10308
rect 27646 10364 27710 10368
rect 27646 10308 27650 10364
rect 27650 10308 27706 10364
rect 27706 10308 27710 10364
rect 27646 10304 27710 10308
rect 27726 10364 27790 10368
rect 27726 10308 27730 10364
rect 27730 10308 27786 10364
rect 27786 10308 27790 10364
rect 27726 10304 27790 10308
rect 27806 10364 27870 10368
rect 27806 10308 27810 10364
rect 27810 10308 27866 10364
rect 27866 10308 27870 10364
rect 27806 10304 27870 10308
rect 27886 10364 27950 10368
rect 27886 10308 27890 10364
rect 27890 10308 27946 10364
rect 27946 10308 27950 10364
rect 27886 10304 27950 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 11438 9820 11502 9824
rect 11438 9764 11442 9820
rect 11442 9764 11498 9820
rect 11498 9764 11502 9820
rect 11438 9760 11502 9764
rect 11518 9820 11582 9824
rect 11518 9764 11522 9820
rect 11522 9764 11578 9820
rect 11578 9764 11582 9820
rect 11518 9760 11582 9764
rect 11598 9820 11662 9824
rect 11598 9764 11602 9820
rect 11602 9764 11658 9820
rect 11658 9764 11662 9820
rect 11598 9760 11662 9764
rect 11678 9820 11742 9824
rect 11678 9764 11682 9820
rect 11682 9764 11738 9820
rect 11738 9764 11742 9820
rect 11678 9760 11742 9764
rect 19212 9820 19276 9824
rect 19212 9764 19216 9820
rect 19216 9764 19272 9820
rect 19272 9764 19276 9820
rect 19212 9760 19276 9764
rect 19292 9820 19356 9824
rect 19292 9764 19296 9820
rect 19296 9764 19352 9820
rect 19352 9764 19356 9820
rect 19292 9760 19356 9764
rect 19372 9820 19436 9824
rect 19372 9764 19376 9820
rect 19376 9764 19432 9820
rect 19432 9764 19436 9820
rect 19372 9760 19436 9764
rect 19452 9820 19516 9824
rect 19452 9764 19456 9820
rect 19456 9764 19512 9820
rect 19512 9764 19516 9820
rect 19452 9760 19516 9764
rect 26986 9820 27050 9824
rect 26986 9764 26990 9820
rect 26990 9764 27046 9820
rect 27046 9764 27050 9820
rect 26986 9760 27050 9764
rect 27066 9820 27130 9824
rect 27066 9764 27070 9820
rect 27070 9764 27126 9820
rect 27126 9764 27130 9820
rect 27066 9760 27130 9764
rect 27146 9820 27210 9824
rect 27146 9764 27150 9820
rect 27150 9764 27206 9820
rect 27206 9764 27210 9820
rect 27146 9760 27210 9764
rect 27226 9820 27290 9824
rect 27226 9764 27230 9820
rect 27230 9764 27286 9820
rect 27286 9764 27290 9820
rect 27226 9760 27290 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 12098 9276 12162 9280
rect 12098 9220 12102 9276
rect 12102 9220 12158 9276
rect 12158 9220 12162 9276
rect 12098 9216 12162 9220
rect 12178 9276 12242 9280
rect 12178 9220 12182 9276
rect 12182 9220 12238 9276
rect 12238 9220 12242 9276
rect 12178 9216 12242 9220
rect 12258 9276 12322 9280
rect 12258 9220 12262 9276
rect 12262 9220 12318 9276
rect 12318 9220 12322 9276
rect 12258 9216 12322 9220
rect 12338 9276 12402 9280
rect 12338 9220 12342 9276
rect 12342 9220 12398 9276
rect 12398 9220 12402 9276
rect 12338 9216 12402 9220
rect 19872 9276 19936 9280
rect 19872 9220 19876 9276
rect 19876 9220 19932 9276
rect 19932 9220 19936 9276
rect 19872 9216 19936 9220
rect 19952 9276 20016 9280
rect 19952 9220 19956 9276
rect 19956 9220 20012 9276
rect 20012 9220 20016 9276
rect 19952 9216 20016 9220
rect 20032 9276 20096 9280
rect 20032 9220 20036 9276
rect 20036 9220 20092 9276
rect 20092 9220 20096 9276
rect 20032 9216 20096 9220
rect 20112 9276 20176 9280
rect 20112 9220 20116 9276
rect 20116 9220 20172 9276
rect 20172 9220 20176 9276
rect 20112 9216 20176 9220
rect 27646 9276 27710 9280
rect 27646 9220 27650 9276
rect 27650 9220 27706 9276
rect 27706 9220 27710 9276
rect 27646 9216 27710 9220
rect 27726 9276 27790 9280
rect 27726 9220 27730 9276
rect 27730 9220 27786 9276
rect 27786 9220 27790 9276
rect 27726 9216 27790 9220
rect 27806 9276 27870 9280
rect 27806 9220 27810 9276
rect 27810 9220 27866 9276
rect 27866 9220 27870 9276
rect 27806 9216 27870 9220
rect 27886 9276 27950 9280
rect 27886 9220 27890 9276
rect 27890 9220 27946 9276
rect 27946 9220 27950 9276
rect 27886 9216 27950 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 11438 8732 11502 8736
rect 11438 8676 11442 8732
rect 11442 8676 11498 8732
rect 11498 8676 11502 8732
rect 11438 8672 11502 8676
rect 11518 8732 11582 8736
rect 11518 8676 11522 8732
rect 11522 8676 11578 8732
rect 11578 8676 11582 8732
rect 11518 8672 11582 8676
rect 11598 8732 11662 8736
rect 11598 8676 11602 8732
rect 11602 8676 11658 8732
rect 11658 8676 11662 8732
rect 11598 8672 11662 8676
rect 11678 8732 11742 8736
rect 11678 8676 11682 8732
rect 11682 8676 11738 8732
rect 11738 8676 11742 8732
rect 11678 8672 11742 8676
rect 19212 8732 19276 8736
rect 19212 8676 19216 8732
rect 19216 8676 19272 8732
rect 19272 8676 19276 8732
rect 19212 8672 19276 8676
rect 19292 8732 19356 8736
rect 19292 8676 19296 8732
rect 19296 8676 19352 8732
rect 19352 8676 19356 8732
rect 19292 8672 19356 8676
rect 19372 8732 19436 8736
rect 19372 8676 19376 8732
rect 19376 8676 19432 8732
rect 19432 8676 19436 8732
rect 19372 8672 19436 8676
rect 19452 8732 19516 8736
rect 19452 8676 19456 8732
rect 19456 8676 19512 8732
rect 19512 8676 19516 8732
rect 19452 8672 19516 8676
rect 26986 8732 27050 8736
rect 26986 8676 26990 8732
rect 26990 8676 27046 8732
rect 27046 8676 27050 8732
rect 26986 8672 27050 8676
rect 27066 8732 27130 8736
rect 27066 8676 27070 8732
rect 27070 8676 27126 8732
rect 27126 8676 27130 8732
rect 27066 8672 27130 8676
rect 27146 8732 27210 8736
rect 27146 8676 27150 8732
rect 27150 8676 27206 8732
rect 27206 8676 27210 8732
rect 27146 8672 27210 8676
rect 27226 8732 27290 8736
rect 27226 8676 27230 8732
rect 27230 8676 27286 8732
rect 27286 8676 27290 8732
rect 27226 8672 27290 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 12098 8188 12162 8192
rect 12098 8132 12102 8188
rect 12102 8132 12158 8188
rect 12158 8132 12162 8188
rect 12098 8128 12162 8132
rect 12178 8188 12242 8192
rect 12178 8132 12182 8188
rect 12182 8132 12238 8188
rect 12238 8132 12242 8188
rect 12178 8128 12242 8132
rect 12258 8188 12322 8192
rect 12258 8132 12262 8188
rect 12262 8132 12318 8188
rect 12318 8132 12322 8188
rect 12258 8128 12322 8132
rect 12338 8188 12402 8192
rect 12338 8132 12342 8188
rect 12342 8132 12398 8188
rect 12398 8132 12402 8188
rect 12338 8128 12402 8132
rect 19872 8188 19936 8192
rect 19872 8132 19876 8188
rect 19876 8132 19932 8188
rect 19932 8132 19936 8188
rect 19872 8128 19936 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 27646 8188 27710 8192
rect 27646 8132 27650 8188
rect 27650 8132 27706 8188
rect 27706 8132 27710 8188
rect 27646 8128 27710 8132
rect 27726 8188 27790 8192
rect 27726 8132 27730 8188
rect 27730 8132 27786 8188
rect 27786 8132 27790 8188
rect 27726 8128 27790 8132
rect 27806 8188 27870 8192
rect 27806 8132 27810 8188
rect 27810 8132 27866 8188
rect 27866 8132 27870 8188
rect 27806 8128 27870 8132
rect 27886 8188 27950 8192
rect 27886 8132 27890 8188
rect 27890 8132 27946 8188
rect 27946 8132 27950 8188
rect 27886 8128 27950 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 11438 7644 11502 7648
rect 11438 7588 11442 7644
rect 11442 7588 11498 7644
rect 11498 7588 11502 7644
rect 11438 7584 11502 7588
rect 11518 7644 11582 7648
rect 11518 7588 11522 7644
rect 11522 7588 11578 7644
rect 11578 7588 11582 7644
rect 11518 7584 11582 7588
rect 11598 7644 11662 7648
rect 11598 7588 11602 7644
rect 11602 7588 11658 7644
rect 11658 7588 11662 7644
rect 11598 7584 11662 7588
rect 11678 7644 11742 7648
rect 11678 7588 11682 7644
rect 11682 7588 11738 7644
rect 11738 7588 11742 7644
rect 11678 7584 11742 7588
rect 19212 7644 19276 7648
rect 19212 7588 19216 7644
rect 19216 7588 19272 7644
rect 19272 7588 19276 7644
rect 19212 7584 19276 7588
rect 19292 7644 19356 7648
rect 19292 7588 19296 7644
rect 19296 7588 19352 7644
rect 19352 7588 19356 7644
rect 19292 7584 19356 7588
rect 19372 7644 19436 7648
rect 19372 7588 19376 7644
rect 19376 7588 19432 7644
rect 19432 7588 19436 7644
rect 19372 7584 19436 7588
rect 19452 7644 19516 7648
rect 19452 7588 19456 7644
rect 19456 7588 19512 7644
rect 19512 7588 19516 7644
rect 19452 7584 19516 7588
rect 26986 7644 27050 7648
rect 26986 7588 26990 7644
rect 26990 7588 27046 7644
rect 27046 7588 27050 7644
rect 26986 7584 27050 7588
rect 27066 7644 27130 7648
rect 27066 7588 27070 7644
rect 27070 7588 27126 7644
rect 27126 7588 27130 7644
rect 27066 7584 27130 7588
rect 27146 7644 27210 7648
rect 27146 7588 27150 7644
rect 27150 7588 27206 7644
rect 27206 7588 27210 7644
rect 27146 7584 27210 7588
rect 27226 7644 27290 7648
rect 27226 7588 27230 7644
rect 27230 7588 27286 7644
rect 27286 7588 27290 7644
rect 27226 7584 27290 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 12098 7100 12162 7104
rect 12098 7044 12102 7100
rect 12102 7044 12158 7100
rect 12158 7044 12162 7100
rect 12098 7040 12162 7044
rect 12178 7100 12242 7104
rect 12178 7044 12182 7100
rect 12182 7044 12238 7100
rect 12238 7044 12242 7100
rect 12178 7040 12242 7044
rect 12258 7100 12322 7104
rect 12258 7044 12262 7100
rect 12262 7044 12318 7100
rect 12318 7044 12322 7100
rect 12258 7040 12322 7044
rect 12338 7100 12402 7104
rect 12338 7044 12342 7100
rect 12342 7044 12398 7100
rect 12398 7044 12402 7100
rect 12338 7040 12402 7044
rect 19872 7100 19936 7104
rect 19872 7044 19876 7100
rect 19876 7044 19932 7100
rect 19932 7044 19936 7100
rect 19872 7040 19936 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 27646 7100 27710 7104
rect 27646 7044 27650 7100
rect 27650 7044 27706 7100
rect 27706 7044 27710 7100
rect 27646 7040 27710 7044
rect 27726 7100 27790 7104
rect 27726 7044 27730 7100
rect 27730 7044 27786 7100
rect 27786 7044 27790 7100
rect 27726 7040 27790 7044
rect 27806 7100 27870 7104
rect 27806 7044 27810 7100
rect 27810 7044 27866 7100
rect 27866 7044 27870 7100
rect 27806 7040 27870 7044
rect 27886 7100 27950 7104
rect 27886 7044 27890 7100
rect 27890 7044 27946 7100
rect 27946 7044 27950 7100
rect 27886 7040 27950 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 11438 6556 11502 6560
rect 11438 6500 11442 6556
rect 11442 6500 11498 6556
rect 11498 6500 11502 6556
rect 11438 6496 11502 6500
rect 11518 6556 11582 6560
rect 11518 6500 11522 6556
rect 11522 6500 11578 6556
rect 11578 6500 11582 6556
rect 11518 6496 11582 6500
rect 11598 6556 11662 6560
rect 11598 6500 11602 6556
rect 11602 6500 11658 6556
rect 11658 6500 11662 6556
rect 11598 6496 11662 6500
rect 11678 6556 11742 6560
rect 11678 6500 11682 6556
rect 11682 6500 11738 6556
rect 11738 6500 11742 6556
rect 11678 6496 11742 6500
rect 19212 6556 19276 6560
rect 19212 6500 19216 6556
rect 19216 6500 19272 6556
rect 19272 6500 19276 6556
rect 19212 6496 19276 6500
rect 19292 6556 19356 6560
rect 19292 6500 19296 6556
rect 19296 6500 19352 6556
rect 19352 6500 19356 6556
rect 19292 6496 19356 6500
rect 19372 6556 19436 6560
rect 19372 6500 19376 6556
rect 19376 6500 19432 6556
rect 19432 6500 19436 6556
rect 19372 6496 19436 6500
rect 19452 6556 19516 6560
rect 19452 6500 19456 6556
rect 19456 6500 19512 6556
rect 19512 6500 19516 6556
rect 19452 6496 19516 6500
rect 26986 6556 27050 6560
rect 26986 6500 26990 6556
rect 26990 6500 27046 6556
rect 27046 6500 27050 6556
rect 26986 6496 27050 6500
rect 27066 6556 27130 6560
rect 27066 6500 27070 6556
rect 27070 6500 27126 6556
rect 27126 6500 27130 6556
rect 27066 6496 27130 6500
rect 27146 6556 27210 6560
rect 27146 6500 27150 6556
rect 27150 6500 27206 6556
rect 27206 6500 27210 6556
rect 27146 6496 27210 6500
rect 27226 6556 27290 6560
rect 27226 6500 27230 6556
rect 27230 6500 27286 6556
rect 27286 6500 27290 6556
rect 27226 6496 27290 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 12098 6012 12162 6016
rect 12098 5956 12102 6012
rect 12102 5956 12158 6012
rect 12158 5956 12162 6012
rect 12098 5952 12162 5956
rect 12178 6012 12242 6016
rect 12178 5956 12182 6012
rect 12182 5956 12238 6012
rect 12238 5956 12242 6012
rect 12178 5952 12242 5956
rect 12258 6012 12322 6016
rect 12258 5956 12262 6012
rect 12262 5956 12318 6012
rect 12318 5956 12322 6012
rect 12258 5952 12322 5956
rect 12338 6012 12402 6016
rect 12338 5956 12342 6012
rect 12342 5956 12398 6012
rect 12398 5956 12402 6012
rect 12338 5952 12402 5956
rect 19872 6012 19936 6016
rect 19872 5956 19876 6012
rect 19876 5956 19932 6012
rect 19932 5956 19936 6012
rect 19872 5952 19936 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 27646 6012 27710 6016
rect 27646 5956 27650 6012
rect 27650 5956 27706 6012
rect 27706 5956 27710 6012
rect 27646 5952 27710 5956
rect 27726 6012 27790 6016
rect 27726 5956 27730 6012
rect 27730 5956 27786 6012
rect 27786 5956 27790 6012
rect 27726 5952 27790 5956
rect 27806 6012 27870 6016
rect 27806 5956 27810 6012
rect 27810 5956 27866 6012
rect 27866 5956 27870 6012
rect 27806 5952 27870 5956
rect 27886 6012 27950 6016
rect 27886 5956 27890 6012
rect 27890 5956 27946 6012
rect 27946 5956 27950 6012
rect 27886 5952 27950 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 11438 5468 11502 5472
rect 11438 5412 11442 5468
rect 11442 5412 11498 5468
rect 11498 5412 11502 5468
rect 11438 5408 11502 5412
rect 11518 5468 11582 5472
rect 11518 5412 11522 5468
rect 11522 5412 11578 5468
rect 11578 5412 11582 5468
rect 11518 5408 11582 5412
rect 11598 5468 11662 5472
rect 11598 5412 11602 5468
rect 11602 5412 11658 5468
rect 11658 5412 11662 5468
rect 11598 5408 11662 5412
rect 11678 5468 11742 5472
rect 11678 5412 11682 5468
rect 11682 5412 11738 5468
rect 11738 5412 11742 5468
rect 11678 5408 11742 5412
rect 19212 5468 19276 5472
rect 19212 5412 19216 5468
rect 19216 5412 19272 5468
rect 19272 5412 19276 5468
rect 19212 5408 19276 5412
rect 19292 5468 19356 5472
rect 19292 5412 19296 5468
rect 19296 5412 19352 5468
rect 19352 5412 19356 5468
rect 19292 5408 19356 5412
rect 19372 5468 19436 5472
rect 19372 5412 19376 5468
rect 19376 5412 19432 5468
rect 19432 5412 19436 5468
rect 19372 5408 19436 5412
rect 19452 5468 19516 5472
rect 19452 5412 19456 5468
rect 19456 5412 19512 5468
rect 19512 5412 19516 5468
rect 19452 5408 19516 5412
rect 26986 5468 27050 5472
rect 26986 5412 26990 5468
rect 26990 5412 27046 5468
rect 27046 5412 27050 5468
rect 26986 5408 27050 5412
rect 27066 5468 27130 5472
rect 27066 5412 27070 5468
rect 27070 5412 27126 5468
rect 27126 5412 27130 5468
rect 27066 5408 27130 5412
rect 27146 5468 27210 5472
rect 27146 5412 27150 5468
rect 27150 5412 27206 5468
rect 27206 5412 27210 5468
rect 27146 5408 27210 5412
rect 27226 5468 27290 5472
rect 27226 5412 27230 5468
rect 27230 5412 27286 5468
rect 27286 5412 27290 5468
rect 27226 5408 27290 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 12098 4924 12162 4928
rect 12098 4868 12102 4924
rect 12102 4868 12158 4924
rect 12158 4868 12162 4924
rect 12098 4864 12162 4868
rect 12178 4924 12242 4928
rect 12178 4868 12182 4924
rect 12182 4868 12238 4924
rect 12238 4868 12242 4924
rect 12178 4864 12242 4868
rect 12258 4924 12322 4928
rect 12258 4868 12262 4924
rect 12262 4868 12318 4924
rect 12318 4868 12322 4924
rect 12258 4864 12322 4868
rect 12338 4924 12402 4928
rect 12338 4868 12342 4924
rect 12342 4868 12398 4924
rect 12398 4868 12402 4924
rect 12338 4864 12402 4868
rect 19872 4924 19936 4928
rect 19872 4868 19876 4924
rect 19876 4868 19932 4924
rect 19932 4868 19936 4924
rect 19872 4864 19936 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 27646 4924 27710 4928
rect 27646 4868 27650 4924
rect 27650 4868 27706 4924
rect 27706 4868 27710 4924
rect 27646 4864 27710 4868
rect 27726 4924 27790 4928
rect 27726 4868 27730 4924
rect 27730 4868 27786 4924
rect 27786 4868 27790 4924
rect 27726 4864 27790 4868
rect 27806 4924 27870 4928
rect 27806 4868 27810 4924
rect 27810 4868 27866 4924
rect 27866 4868 27870 4924
rect 27806 4864 27870 4868
rect 27886 4924 27950 4928
rect 27886 4868 27890 4924
rect 27890 4868 27946 4924
rect 27946 4868 27950 4924
rect 27886 4864 27950 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 11438 4380 11502 4384
rect 11438 4324 11442 4380
rect 11442 4324 11498 4380
rect 11498 4324 11502 4380
rect 11438 4320 11502 4324
rect 11518 4380 11582 4384
rect 11518 4324 11522 4380
rect 11522 4324 11578 4380
rect 11578 4324 11582 4380
rect 11518 4320 11582 4324
rect 11598 4380 11662 4384
rect 11598 4324 11602 4380
rect 11602 4324 11658 4380
rect 11658 4324 11662 4380
rect 11598 4320 11662 4324
rect 11678 4380 11742 4384
rect 11678 4324 11682 4380
rect 11682 4324 11738 4380
rect 11738 4324 11742 4380
rect 11678 4320 11742 4324
rect 19212 4380 19276 4384
rect 19212 4324 19216 4380
rect 19216 4324 19272 4380
rect 19272 4324 19276 4380
rect 19212 4320 19276 4324
rect 19292 4380 19356 4384
rect 19292 4324 19296 4380
rect 19296 4324 19352 4380
rect 19352 4324 19356 4380
rect 19292 4320 19356 4324
rect 19372 4380 19436 4384
rect 19372 4324 19376 4380
rect 19376 4324 19432 4380
rect 19432 4324 19436 4380
rect 19372 4320 19436 4324
rect 19452 4380 19516 4384
rect 19452 4324 19456 4380
rect 19456 4324 19512 4380
rect 19512 4324 19516 4380
rect 19452 4320 19516 4324
rect 26986 4380 27050 4384
rect 26986 4324 26990 4380
rect 26990 4324 27046 4380
rect 27046 4324 27050 4380
rect 26986 4320 27050 4324
rect 27066 4380 27130 4384
rect 27066 4324 27070 4380
rect 27070 4324 27126 4380
rect 27126 4324 27130 4380
rect 27066 4320 27130 4324
rect 27146 4380 27210 4384
rect 27146 4324 27150 4380
rect 27150 4324 27206 4380
rect 27206 4324 27210 4380
rect 27146 4320 27210 4324
rect 27226 4380 27290 4384
rect 27226 4324 27230 4380
rect 27230 4324 27286 4380
rect 27286 4324 27290 4380
rect 27226 4320 27290 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 12098 3836 12162 3840
rect 12098 3780 12102 3836
rect 12102 3780 12158 3836
rect 12158 3780 12162 3836
rect 12098 3776 12162 3780
rect 12178 3836 12242 3840
rect 12178 3780 12182 3836
rect 12182 3780 12238 3836
rect 12238 3780 12242 3836
rect 12178 3776 12242 3780
rect 12258 3836 12322 3840
rect 12258 3780 12262 3836
rect 12262 3780 12318 3836
rect 12318 3780 12322 3836
rect 12258 3776 12322 3780
rect 12338 3836 12402 3840
rect 12338 3780 12342 3836
rect 12342 3780 12398 3836
rect 12398 3780 12402 3836
rect 12338 3776 12402 3780
rect 19872 3836 19936 3840
rect 19872 3780 19876 3836
rect 19876 3780 19932 3836
rect 19932 3780 19936 3836
rect 19872 3776 19936 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 27646 3836 27710 3840
rect 27646 3780 27650 3836
rect 27650 3780 27706 3836
rect 27706 3780 27710 3836
rect 27646 3776 27710 3780
rect 27726 3836 27790 3840
rect 27726 3780 27730 3836
rect 27730 3780 27786 3836
rect 27786 3780 27790 3836
rect 27726 3776 27790 3780
rect 27806 3836 27870 3840
rect 27806 3780 27810 3836
rect 27810 3780 27866 3836
rect 27866 3780 27870 3836
rect 27806 3776 27870 3780
rect 27886 3836 27950 3840
rect 27886 3780 27890 3836
rect 27890 3780 27946 3836
rect 27946 3780 27950 3836
rect 27886 3776 27950 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 11438 3292 11502 3296
rect 11438 3236 11442 3292
rect 11442 3236 11498 3292
rect 11498 3236 11502 3292
rect 11438 3232 11502 3236
rect 11518 3292 11582 3296
rect 11518 3236 11522 3292
rect 11522 3236 11578 3292
rect 11578 3236 11582 3292
rect 11518 3232 11582 3236
rect 11598 3292 11662 3296
rect 11598 3236 11602 3292
rect 11602 3236 11658 3292
rect 11658 3236 11662 3292
rect 11598 3232 11662 3236
rect 11678 3292 11742 3296
rect 11678 3236 11682 3292
rect 11682 3236 11738 3292
rect 11738 3236 11742 3292
rect 11678 3232 11742 3236
rect 19212 3292 19276 3296
rect 19212 3236 19216 3292
rect 19216 3236 19272 3292
rect 19272 3236 19276 3292
rect 19212 3232 19276 3236
rect 19292 3292 19356 3296
rect 19292 3236 19296 3292
rect 19296 3236 19352 3292
rect 19352 3236 19356 3292
rect 19292 3232 19356 3236
rect 19372 3292 19436 3296
rect 19372 3236 19376 3292
rect 19376 3236 19432 3292
rect 19432 3236 19436 3292
rect 19372 3232 19436 3236
rect 19452 3292 19516 3296
rect 19452 3236 19456 3292
rect 19456 3236 19512 3292
rect 19512 3236 19516 3292
rect 19452 3232 19516 3236
rect 26986 3292 27050 3296
rect 26986 3236 26990 3292
rect 26990 3236 27046 3292
rect 27046 3236 27050 3292
rect 26986 3232 27050 3236
rect 27066 3292 27130 3296
rect 27066 3236 27070 3292
rect 27070 3236 27126 3292
rect 27126 3236 27130 3292
rect 27066 3232 27130 3236
rect 27146 3292 27210 3296
rect 27146 3236 27150 3292
rect 27150 3236 27206 3292
rect 27206 3236 27210 3292
rect 27146 3232 27210 3236
rect 27226 3292 27290 3296
rect 27226 3236 27230 3292
rect 27230 3236 27286 3292
rect 27286 3236 27290 3292
rect 27226 3232 27290 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 12098 2748 12162 2752
rect 12098 2692 12102 2748
rect 12102 2692 12158 2748
rect 12158 2692 12162 2748
rect 12098 2688 12162 2692
rect 12178 2748 12242 2752
rect 12178 2692 12182 2748
rect 12182 2692 12238 2748
rect 12238 2692 12242 2748
rect 12178 2688 12242 2692
rect 12258 2748 12322 2752
rect 12258 2692 12262 2748
rect 12262 2692 12318 2748
rect 12318 2692 12322 2748
rect 12258 2688 12322 2692
rect 12338 2748 12402 2752
rect 12338 2692 12342 2748
rect 12342 2692 12398 2748
rect 12398 2692 12402 2748
rect 12338 2688 12402 2692
rect 19872 2748 19936 2752
rect 19872 2692 19876 2748
rect 19876 2692 19932 2748
rect 19932 2692 19936 2748
rect 19872 2688 19936 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 27646 2748 27710 2752
rect 27646 2692 27650 2748
rect 27650 2692 27706 2748
rect 27706 2692 27710 2748
rect 27646 2688 27710 2692
rect 27726 2748 27790 2752
rect 27726 2692 27730 2748
rect 27730 2692 27786 2748
rect 27786 2692 27790 2748
rect 27726 2688 27790 2692
rect 27806 2748 27870 2752
rect 27806 2692 27810 2748
rect 27810 2692 27866 2748
rect 27866 2692 27870 2748
rect 27806 2688 27870 2692
rect 27886 2748 27950 2752
rect 27886 2692 27890 2748
rect 27890 2692 27946 2748
rect 27946 2692 27950 2748
rect 27886 2688 27950 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 11438 2204 11502 2208
rect 11438 2148 11442 2204
rect 11442 2148 11498 2204
rect 11498 2148 11502 2204
rect 11438 2144 11502 2148
rect 11518 2204 11582 2208
rect 11518 2148 11522 2204
rect 11522 2148 11578 2204
rect 11578 2148 11582 2204
rect 11518 2144 11582 2148
rect 11598 2204 11662 2208
rect 11598 2148 11602 2204
rect 11602 2148 11658 2204
rect 11658 2148 11662 2204
rect 11598 2144 11662 2148
rect 11678 2204 11742 2208
rect 11678 2148 11682 2204
rect 11682 2148 11738 2204
rect 11738 2148 11742 2204
rect 11678 2144 11742 2148
rect 19212 2204 19276 2208
rect 19212 2148 19216 2204
rect 19216 2148 19272 2204
rect 19272 2148 19276 2204
rect 19212 2144 19276 2148
rect 19292 2204 19356 2208
rect 19292 2148 19296 2204
rect 19296 2148 19352 2204
rect 19352 2148 19356 2204
rect 19292 2144 19356 2148
rect 19372 2204 19436 2208
rect 19372 2148 19376 2204
rect 19376 2148 19432 2204
rect 19432 2148 19436 2204
rect 19372 2144 19436 2148
rect 19452 2204 19516 2208
rect 19452 2148 19456 2204
rect 19456 2148 19512 2204
rect 19512 2148 19516 2204
rect 19452 2144 19516 2148
rect 26986 2204 27050 2208
rect 26986 2148 26990 2204
rect 26990 2148 27046 2204
rect 27046 2148 27050 2204
rect 26986 2144 27050 2148
rect 27066 2204 27130 2208
rect 27066 2148 27070 2204
rect 27070 2148 27126 2204
rect 27126 2148 27130 2204
rect 27066 2144 27130 2148
rect 27146 2204 27210 2208
rect 27146 2148 27150 2204
rect 27150 2148 27206 2204
rect 27206 2148 27210 2204
rect 27146 2144 27210 2148
rect 27226 2204 27290 2208
rect 27226 2148 27230 2204
rect 27230 2148 27286 2204
rect 27286 2148 27290 2204
rect 27226 2144 27290 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 12098 1660 12162 1664
rect 12098 1604 12102 1660
rect 12102 1604 12158 1660
rect 12158 1604 12162 1660
rect 12098 1600 12162 1604
rect 12178 1660 12242 1664
rect 12178 1604 12182 1660
rect 12182 1604 12238 1660
rect 12238 1604 12242 1660
rect 12178 1600 12242 1604
rect 12258 1660 12322 1664
rect 12258 1604 12262 1660
rect 12262 1604 12318 1660
rect 12318 1604 12322 1660
rect 12258 1600 12322 1604
rect 12338 1660 12402 1664
rect 12338 1604 12342 1660
rect 12342 1604 12398 1660
rect 12398 1604 12402 1660
rect 12338 1600 12402 1604
rect 19872 1660 19936 1664
rect 19872 1604 19876 1660
rect 19876 1604 19932 1660
rect 19932 1604 19936 1660
rect 19872 1600 19936 1604
rect 19952 1660 20016 1664
rect 19952 1604 19956 1660
rect 19956 1604 20012 1660
rect 20012 1604 20016 1660
rect 19952 1600 20016 1604
rect 20032 1660 20096 1664
rect 20032 1604 20036 1660
rect 20036 1604 20092 1660
rect 20092 1604 20096 1660
rect 20032 1600 20096 1604
rect 20112 1660 20176 1664
rect 20112 1604 20116 1660
rect 20116 1604 20172 1660
rect 20172 1604 20176 1660
rect 20112 1600 20176 1604
rect 27646 1660 27710 1664
rect 27646 1604 27650 1660
rect 27650 1604 27706 1660
rect 27706 1604 27710 1660
rect 27646 1600 27710 1604
rect 27726 1660 27790 1664
rect 27726 1604 27730 1660
rect 27730 1604 27786 1660
rect 27786 1604 27790 1660
rect 27726 1600 27790 1604
rect 27806 1660 27870 1664
rect 27806 1604 27810 1660
rect 27810 1604 27866 1660
rect 27866 1604 27870 1660
rect 27806 1600 27870 1604
rect 27886 1660 27950 1664
rect 27886 1604 27890 1660
rect 27890 1604 27946 1660
rect 27946 1604 27950 1660
rect 27886 1600 27950 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 11438 1116 11502 1120
rect 11438 1060 11442 1116
rect 11442 1060 11498 1116
rect 11498 1060 11502 1116
rect 11438 1056 11502 1060
rect 11518 1116 11582 1120
rect 11518 1060 11522 1116
rect 11522 1060 11578 1116
rect 11578 1060 11582 1116
rect 11518 1056 11582 1060
rect 11598 1116 11662 1120
rect 11598 1060 11602 1116
rect 11602 1060 11658 1116
rect 11658 1060 11662 1116
rect 11598 1056 11662 1060
rect 11678 1116 11742 1120
rect 11678 1060 11682 1116
rect 11682 1060 11738 1116
rect 11738 1060 11742 1116
rect 11678 1056 11742 1060
rect 19212 1116 19276 1120
rect 19212 1060 19216 1116
rect 19216 1060 19272 1116
rect 19272 1060 19276 1116
rect 19212 1056 19276 1060
rect 19292 1116 19356 1120
rect 19292 1060 19296 1116
rect 19296 1060 19352 1116
rect 19352 1060 19356 1116
rect 19292 1056 19356 1060
rect 19372 1116 19436 1120
rect 19372 1060 19376 1116
rect 19376 1060 19432 1116
rect 19432 1060 19436 1116
rect 19372 1056 19436 1060
rect 19452 1116 19516 1120
rect 19452 1060 19456 1116
rect 19456 1060 19512 1116
rect 19512 1060 19516 1116
rect 19452 1056 19516 1060
rect 26986 1116 27050 1120
rect 26986 1060 26990 1116
rect 26990 1060 27046 1116
rect 27046 1060 27050 1116
rect 26986 1056 27050 1060
rect 27066 1116 27130 1120
rect 27066 1060 27070 1116
rect 27070 1060 27126 1116
rect 27126 1060 27130 1116
rect 27066 1056 27130 1060
rect 27146 1116 27210 1120
rect 27146 1060 27150 1116
rect 27150 1060 27206 1116
rect 27206 1060 27210 1116
rect 27146 1056 27210 1060
rect 27226 1116 27290 1120
rect 27226 1060 27230 1116
rect 27230 1060 27286 1116
rect 27286 1060 27290 1116
rect 27226 1056 27290 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 12098 572 12162 576
rect 12098 516 12102 572
rect 12102 516 12158 572
rect 12158 516 12162 572
rect 12098 512 12162 516
rect 12178 572 12242 576
rect 12178 516 12182 572
rect 12182 516 12238 572
rect 12238 516 12242 572
rect 12178 512 12242 516
rect 12258 572 12322 576
rect 12258 516 12262 572
rect 12262 516 12318 572
rect 12318 516 12322 572
rect 12258 512 12322 516
rect 12338 572 12402 576
rect 12338 516 12342 572
rect 12342 516 12398 572
rect 12398 516 12402 572
rect 12338 512 12402 516
rect 19872 572 19936 576
rect 19872 516 19876 572
rect 19876 516 19932 572
rect 19932 516 19936 572
rect 19872 512 19936 516
rect 19952 572 20016 576
rect 19952 516 19956 572
rect 19956 516 20012 572
rect 20012 516 20016 572
rect 19952 512 20016 516
rect 20032 572 20096 576
rect 20032 516 20036 572
rect 20036 516 20092 572
rect 20092 516 20096 572
rect 20032 512 20096 516
rect 20112 572 20176 576
rect 20112 516 20116 572
rect 20116 516 20172 572
rect 20172 516 20176 572
rect 20112 512 20176 516
rect 27646 572 27710 576
rect 27646 516 27650 572
rect 27650 516 27706 572
rect 27706 516 27710 572
rect 27646 512 27710 516
rect 27726 572 27790 576
rect 27726 516 27730 572
rect 27730 516 27786 572
rect 27786 516 27790 572
rect 27726 512 27790 516
rect 27806 572 27870 576
rect 27806 516 27810 572
rect 27810 516 27866 572
rect 27866 516 27870 572
rect 27806 512 27870 516
rect 27886 572 27950 576
rect 27886 516 27890 572
rect 27890 516 27946 572
rect 27946 516 27950 572
rect 27886 512 27950 516
<< metal4 >>
rect 3656 21792 3976 21808
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 21248 4636 21808
rect 6134 21725 6194 22304
rect 6131 21724 6197 21725
rect 6131 21660 6132 21724
rect 6196 21660 6197 21724
rect 6131 21659 6197 21660
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 6686 21181 6746 22304
rect 7238 21725 7298 22304
rect 7790 21861 7850 22304
rect 7787 21860 7853 21861
rect 7787 21796 7788 21860
rect 7852 21796 7853 21860
rect 7787 21795 7853 21796
rect 8342 21725 8402 22304
rect 7235 21724 7301 21725
rect 7235 21660 7236 21724
rect 7300 21660 7301 21724
rect 7235 21659 7301 21660
rect 8339 21724 8405 21725
rect 8339 21660 8340 21724
rect 8404 21660 8405 21724
rect 8339 21659 8405 21660
rect 6683 21180 6749 21181
rect 6683 21116 6684 21180
rect 6748 21116 6749 21180
rect 6683 21115 6749 21116
rect 8894 20637 8954 22304
rect 9446 21181 9506 22304
rect 9998 21725 10058 22304
rect 10550 21725 10610 22304
rect 9995 21724 10061 21725
rect 9995 21660 9996 21724
rect 10060 21660 10061 21724
rect 9995 21659 10061 21660
rect 10547 21724 10613 21725
rect 10547 21660 10548 21724
rect 10612 21660 10613 21724
rect 10547 21659 10613 21660
rect 11102 21589 11162 22304
rect 11654 21997 11714 22304
rect 12206 21997 12266 22304
rect 11651 21996 11717 21997
rect 11651 21932 11652 21996
rect 11716 21932 11717 21996
rect 11651 21931 11717 21932
rect 12203 21996 12269 21997
rect 12203 21932 12204 21996
rect 12268 21932 12269 21996
rect 12203 21931 12269 21932
rect 11430 21792 11750 21808
rect 11430 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11750 21792
rect 11099 21588 11165 21589
rect 11099 21524 11100 21588
rect 11164 21524 11165 21588
rect 11099 21523 11165 21524
rect 9443 21180 9509 21181
rect 9443 21116 9444 21180
rect 9508 21116 9509 21180
rect 9443 21115 9509 21116
rect 10179 20772 10245 20773
rect 10179 20708 10180 20772
rect 10244 20708 10245 20772
rect 10179 20707 10245 20708
rect 8891 20636 8957 20637
rect 8891 20572 8892 20636
rect 8956 20572 8957 20636
rect 8891 20571 8957 20572
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 10182 11933 10242 20707
rect 11430 20704 11750 21728
rect 11430 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11750 20704
rect 11430 19616 11750 20640
rect 11430 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11750 19616
rect 11430 18528 11750 19552
rect 11430 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11750 18528
rect 11430 17440 11750 18464
rect 11430 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11750 17440
rect 11430 16352 11750 17376
rect 11430 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11750 16352
rect 11430 15264 11750 16288
rect 11430 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11750 15264
rect 11430 14176 11750 15200
rect 11430 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11750 14176
rect 11430 13088 11750 14112
rect 11430 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11750 13088
rect 11430 12000 11750 13024
rect 11430 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11750 12000
rect 10179 11932 10245 11933
rect 10179 11868 10180 11932
rect 10244 11868 10245 11932
rect 10179 11867 10245 11868
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 11430 10912 11750 11936
rect 11430 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11750 10912
rect 11430 9824 11750 10848
rect 11430 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11750 9824
rect 11430 8736 11750 9760
rect 11430 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11750 8736
rect 11430 7648 11750 8672
rect 11430 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11750 7648
rect 11430 6560 11750 7584
rect 11430 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11750 6560
rect 11430 5472 11750 6496
rect 11430 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11750 5472
rect 11430 4384 11750 5408
rect 11430 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11750 4384
rect 11430 3296 11750 4320
rect 11430 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11750 3296
rect 11430 2208 11750 3232
rect 11430 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11750 2208
rect 11430 1120 11750 2144
rect 11430 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11750 1120
rect 11430 496 11750 1056
rect 12090 21248 12410 21808
rect 12758 21725 12818 22304
rect 12755 21724 12821 21725
rect 12755 21660 12756 21724
rect 12820 21660 12821 21724
rect 12755 21659 12821 21660
rect 12090 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12410 21248
rect 12090 20160 12410 21184
rect 13310 20637 13370 22304
rect 13862 21181 13922 22304
rect 13859 21180 13925 21181
rect 13859 21116 13860 21180
rect 13924 21116 13925 21180
rect 13859 21115 13925 21116
rect 14414 20637 14474 22304
rect 13307 20636 13373 20637
rect 13307 20572 13308 20636
rect 13372 20572 13373 20636
rect 13307 20571 13373 20572
rect 14411 20636 14477 20637
rect 14411 20572 14412 20636
rect 14476 20572 14477 20636
rect 14411 20571 14477 20572
rect 12090 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12410 20160
rect 12090 19072 12410 20096
rect 12090 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12410 19072
rect 12090 17984 12410 19008
rect 14966 18461 15026 22304
rect 15518 21045 15578 22304
rect 15515 21044 15581 21045
rect 15515 20980 15516 21044
rect 15580 20980 15581 21044
rect 15515 20979 15581 20980
rect 16070 18869 16130 22304
rect 16622 19957 16682 22304
rect 17174 20773 17234 22304
rect 17726 21589 17786 22304
rect 17723 21588 17789 21589
rect 17723 21524 17724 21588
rect 17788 21524 17789 21588
rect 17723 21523 17789 21524
rect 18278 21453 18338 22304
rect 18830 21589 18890 22304
rect 19382 22104 19442 22304
rect 19934 22104 19994 22304
rect 20486 22104 20546 22304
rect 21038 22104 21098 22304
rect 21590 21861 21650 22304
rect 22142 22104 22202 22304
rect 22694 22104 22754 22304
rect 23246 22104 23306 22304
rect 23798 21997 23858 22304
rect 23795 21996 23861 21997
rect 23795 21932 23796 21996
rect 23860 21932 23861 21996
rect 23795 21931 23861 21932
rect 24350 21861 24410 22304
rect 24902 21997 24962 22304
rect 25454 21997 25514 22304
rect 26006 21997 26066 22304
rect 24899 21996 24965 21997
rect 24899 21932 24900 21996
rect 24964 21932 24965 21996
rect 24899 21931 24965 21932
rect 25451 21996 25517 21997
rect 25451 21932 25452 21996
rect 25516 21932 25517 21996
rect 25451 21931 25517 21932
rect 26003 21996 26069 21997
rect 26003 21932 26004 21996
rect 26068 21932 26069 21996
rect 26003 21931 26069 21932
rect 26558 21861 26618 22304
rect 27110 21997 27170 22304
rect 27662 21997 27722 22304
rect 27107 21996 27173 21997
rect 27107 21932 27108 21996
rect 27172 21932 27173 21996
rect 27107 21931 27173 21932
rect 27659 21996 27725 21997
rect 27659 21932 27660 21996
rect 27724 21932 27725 21996
rect 27659 21931 27725 21932
rect 28214 21861 28274 22304
rect 21587 21860 21653 21861
rect 19204 21792 19524 21808
rect 19204 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19524 21792
rect 18827 21588 18893 21589
rect 18827 21524 18828 21588
rect 18892 21524 18893 21588
rect 18827 21523 18893 21524
rect 18275 21452 18341 21453
rect 18275 21388 18276 21452
rect 18340 21388 18341 21452
rect 18275 21387 18341 21388
rect 17171 20772 17237 20773
rect 17171 20708 17172 20772
rect 17236 20708 17237 20772
rect 17171 20707 17237 20708
rect 19204 20704 19524 21728
rect 19204 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19524 20704
rect 16619 19956 16685 19957
rect 16619 19892 16620 19956
rect 16684 19892 16685 19956
rect 16619 19891 16685 19892
rect 19204 19616 19524 20640
rect 19204 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19524 19616
rect 16803 19276 16869 19277
rect 16803 19212 16804 19276
rect 16868 19212 16869 19276
rect 16803 19211 16869 19212
rect 16067 18868 16133 18869
rect 16067 18804 16068 18868
rect 16132 18804 16133 18868
rect 16067 18803 16133 18804
rect 14963 18460 15029 18461
rect 14963 18396 14964 18460
rect 15028 18396 15029 18460
rect 14963 18395 15029 18396
rect 12090 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12410 17984
rect 12090 16896 12410 17920
rect 16806 17373 16866 19211
rect 19204 18528 19524 19552
rect 19204 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19524 18528
rect 19204 17440 19524 18464
rect 19204 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19524 17440
rect 16803 17372 16869 17373
rect 16803 17308 16804 17372
rect 16868 17308 16869 17372
rect 16803 17307 16869 17308
rect 12090 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12410 16896
rect 12090 15808 12410 16832
rect 12090 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12410 15808
rect 12090 14720 12410 15744
rect 12090 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12410 14720
rect 12090 13632 12410 14656
rect 12090 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12410 13632
rect 12090 12544 12410 13568
rect 12090 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12410 12544
rect 12090 11456 12410 12480
rect 12090 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12410 11456
rect 12090 10368 12410 11392
rect 12090 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12410 10368
rect 12090 9280 12410 10304
rect 12090 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12410 9280
rect 12090 8192 12410 9216
rect 12090 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12410 8192
rect 12090 7104 12410 8128
rect 12090 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12410 7104
rect 12090 6016 12410 7040
rect 12090 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12410 6016
rect 12090 4928 12410 5952
rect 12090 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12410 4928
rect 12090 3840 12410 4864
rect 12090 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12410 3840
rect 12090 2752 12410 3776
rect 12090 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12410 2752
rect 12090 1664 12410 2688
rect 12090 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12410 1664
rect 12090 576 12410 1600
rect 12090 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12410 576
rect 12090 496 12410 512
rect 19204 16352 19524 17376
rect 19204 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19524 16352
rect 19204 15264 19524 16288
rect 19204 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19524 15264
rect 19204 14176 19524 15200
rect 19204 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19524 14176
rect 19204 13088 19524 14112
rect 19204 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19524 13088
rect 19204 12000 19524 13024
rect 19204 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19524 12000
rect 19204 10912 19524 11936
rect 19204 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19524 10912
rect 19204 9824 19524 10848
rect 19204 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19524 9824
rect 19204 8736 19524 9760
rect 19204 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19524 8736
rect 19204 7648 19524 8672
rect 19204 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19524 7648
rect 19204 6560 19524 7584
rect 19204 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19524 6560
rect 19204 5472 19524 6496
rect 19204 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19524 5472
rect 19204 4384 19524 5408
rect 19204 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19524 4384
rect 19204 3296 19524 4320
rect 19204 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19524 3296
rect 19204 2208 19524 3232
rect 19204 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19524 2208
rect 19204 1120 19524 2144
rect 19204 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19524 1120
rect 19204 496 19524 1056
rect 19864 21248 20184 21808
rect 21587 21796 21588 21860
rect 21652 21796 21653 21860
rect 21587 21795 21653 21796
rect 24347 21860 24413 21861
rect 24347 21796 24348 21860
rect 24412 21796 24413 21860
rect 24347 21795 24413 21796
rect 26555 21860 26621 21861
rect 26555 21796 26556 21860
rect 26620 21796 26621 21860
rect 28211 21860 28277 21861
rect 26555 21795 26621 21796
rect 19864 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20184 21248
rect 19864 20160 20184 21184
rect 19864 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20184 20160
rect 19864 19072 20184 20096
rect 19864 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20184 19072
rect 19864 17984 20184 19008
rect 26978 21792 27298 21808
rect 26978 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27298 21792
rect 26978 20704 27298 21728
rect 26978 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27298 20704
rect 26978 19616 27298 20640
rect 26978 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27298 19616
rect 20299 18596 20365 18597
rect 20299 18532 20300 18596
rect 20364 18532 20365 18596
rect 20299 18531 20365 18532
rect 20483 18596 20549 18597
rect 20483 18532 20484 18596
rect 20548 18532 20549 18596
rect 20483 18531 20549 18532
rect 19864 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20184 17984
rect 19864 16896 20184 17920
rect 19864 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20184 16896
rect 19864 15808 20184 16832
rect 19864 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20184 15808
rect 19864 14720 20184 15744
rect 19864 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20184 14720
rect 19864 13632 20184 14656
rect 19864 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20184 13632
rect 19864 12544 20184 13568
rect 20302 13429 20362 18531
rect 20486 18053 20546 18531
rect 26978 18528 27298 19552
rect 26978 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27298 18528
rect 20483 18052 20549 18053
rect 20483 17988 20484 18052
rect 20548 17988 20549 18052
rect 20483 17987 20549 17988
rect 20486 15469 20546 17987
rect 26978 17440 27298 18464
rect 26978 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27298 17440
rect 26978 16352 27298 17376
rect 26978 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27298 16352
rect 20483 15468 20549 15469
rect 20483 15404 20484 15468
rect 20548 15404 20549 15468
rect 20483 15403 20549 15404
rect 26978 15264 27298 16288
rect 26978 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27298 15264
rect 26978 14176 27298 15200
rect 26978 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27298 14176
rect 20299 13428 20365 13429
rect 20299 13364 20300 13428
rect 20364 13364 20365 13428
rect 20299 13363 20365 13364
rect 19864 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20184 12544
rect 19864 11456 20184 12480
rect 19864 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20184 11456
rect 19864 10368 20184 11392
rect 19864 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20184 10368
rect 19864 9280 20184 10304
rect 19864 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20184 9280
rect 19864 8192 20184 9216
rect 19864 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20184 8192
rect 19864 7104 20184 8128
rect 19864 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20184 7104
rect 19864 6016 20184 7040
rect 19864 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20184 6016
rect 19864 4928 20184 5952
rect 19864 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20184 4928
rect 19864 3840 20184 4864
rect 19864 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20184 3840
rect 19864 2752 20184 3776
rect 19864 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20184 2752
rect 19864 1664 20184 2688
rect 19864 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20184 1664
rect 19864 576 20184 1600
rect 19864 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20184 576
rect 19864 496 20184 512
rect 26978 13088 27298 14112
rect 26978 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27298 13088
rect 26978 12000 27298 13024
rect 26978 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27298 12000
rect 26978 10912 27298 11936
rect 26978 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27298 10912
rect 26978 9824 27298 10848
rect 26978 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27298 9824
rect 26978 8736 27298 9760
rect 26978 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27298 8736
rect 26978 7648 27298 8672
rect 26978 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27298 7648
rect 26978 6560 27298 7584
rect 26978 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27298 6560
rect 26978 5472 27298 6496
rect 26978 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27298 5472
rect 26978 4384 27298 5408
rect 26978 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27298 4384
rect 26978 3296 27298 4320
rect 26978 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27298 3296
rect 26978 2208 27298 3232
rect 26978 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27298 2208
rect 26978 1120 27298 2144
rect 26978 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27298 1120
rect 26978 496 27298 1056
rect 27638 21248 27958 21808
rect 28211 21796 28212 21860
rect 28276 21796 28277 21860
rect 28211 21795 28277 21796
rect 27638 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27958 21248
rect 27638 20160 27958 21184
rect 27638 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27958 20160
rect 27638 19072 27958 20096
rect 27638 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27958 19072
rect 27638 17984 27958 19008
rect 28766 18053 28826 22304
rect 29318 22104 29378 22304
rect 28763 18052 28829 18053
rect 28763 17988 28764 18052
rect 28828 17988 28829 18052
rect 28763 17987 28829 17988
rect 27638 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27958 17984
rect 27638 16896 27958 17920
rect 27638 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27958 16896
rect 27638 15808 27958 16832
rect 27638 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27958 15808
rect 27638 14720 27958 15744
rect 27638 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27958 14720
rect 27638 13632 27958 14656
rect 27638 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27958 13632
rect 27638 12544 27958 13568
rect 27638 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27958 12544
rect 27638 11456 27958 12480
rect 27638 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27958 11456
rect 27638 10368 27958 11392
rect 27638 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27958 10368
rect 27638 9280 27958 10304
rect 27638 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27958 9280
rect 27638 8192 27958 9216
rect 27638 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27958 8192
rect 27638 7104 27958 8128
rect 27638 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27958 7104
rect 27638 6016 27958 7040
rect 27638 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27958 6016
rect 27638 4928 27958 5952
rect 27638 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27958 4928
rect 27638 3840 27958 4864
rect 27638 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27958 3840
rect 27638 2752 27958 3776
rect 27638 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27958 2752
rect 27638 1664 27958 2688
rect 27638 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27958 1664
rect 27638 576 27958 1600
rect 27638 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27958 576
rect 27638 496 27958 512
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1
transform 1 0 6256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1
transform 1 0 6716 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1
transform -1 0 7084 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1
transform 1 0 7820 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1
transform -1 0 11224 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1
transform -1 0 10396 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1
transform -1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1
transform -1 0 14352 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1
transform -1 0 23000 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1
transform 1 0 9384 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1
transform -1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1
transform -1 0 29164 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1
transform -1 0 27048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1
transform -1 0 26680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1
transform -1 0 27048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1
transform 1 0 11132 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1
transform -1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1
transform -1 0 18032 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1
transform -1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1
transform -1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1
transform -1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1
transform -1 0 9384 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1
transform -1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1
transform 1 0 7636 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1
transform 1 0 7544 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1
transform 1 0 5152 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753__1
timestamp 1
transform -1 0 12328 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753__2
timestamp 1
transform -1 0 11316 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0754_
timestamp 1
transform 1 0 5796 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _0755_
timestamp 1
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _0756_
timestamp 1
transform -1 0 7820 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__mux4_1  _0757_
timestamp 1
transform -1 0 26312 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0758_
timestamp 1
transform -1 0 25852 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0759_
timestamp 1
transform 1 0 20976 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _0760_
timestamp 1
transform -1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _0761_
timestamp 1
transform -1 0 27324 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0762_
timestamp 1
transform -1 0 28060 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1
transform 1 0 25300 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _0764_
timestamp 1
transform 1 0 20516 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0765_
timestamp 1
transform -1 0 9936 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0766_
timestamp 1
transform 1 0 6164 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0767_
timestamp 1
transform -1 0 10396 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0768_
timestamp 1
transform -1 0 9016 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0769_
timestamp 1
transform -1 0 9568 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0770_
timestamp 1
transform -1 0 9844 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1
transform 1 0 7728 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 1
transform 1 0 7452 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0773_
timestamp 1
transform 1 0 6256 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0774_
timestamp 1
transform 1 0 8556 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0775_
timestamp 1
transform 1 0 7176 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0776_
timestamp 1
transform -1 0 10856 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0777_
timestamp 1
transform -1 0 9936 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0778_
timestamp 1
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0779_
timestamp 1
transform 1 0 4232 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0780_
timestamp 1
transform 1 0 5888 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0781_
timestamp 1
transform 1 0 4508 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0782_
timestamp 1
transform 1 0 7268 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_1  _0783_
timestamp 1
transform 1 0 6440 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0784_
timestamp 1
transform -1 0 9384 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_1  _0785_
timestamp 1
transform 1 0 9476 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0786_
timestamp 1
transform 1 0 8832 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0787_
timestamp 1
transform 1 0 8372 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0788_
timestamp 1
transform 1 0 7728 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0789_
timestamp 1
transform 1 0 7452 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0790_
timestamp 1
transform -1 0 9108 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _0791_
timestamp 1
transform 1 0 13800 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0792_
timestamp 1
transform 1 0 6808 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0793_
timestamp 1
transform 1 0 3496 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0794_
timestamp 1
transform 1 0 1196 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0795_
timestamp 1
transform -1 0 3956 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0796_
timestamp 1
transform -1 0 4416 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0797_
timestamp 1
transform 1 0 3404 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0798_
timestamp 1
transform -1 0 2760 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0799_
timestamp 1
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1
transform 1 0 12972 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0801_
timestamp 1
transform 1 0 11408 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0803_
timestamp 1
transform 1 0 6992 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0804_
timestamp 1
transform 1 0 2392 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0805_
timestamp 1
transform -1 0 2484 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0806_
timestamp 1
transform 1 0 3220 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0807_
timestamp 1
transform -1 0 2392 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0808_
timestamp 1
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0809_
timestamp 1
transform -1 0 3220 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0810_
timestamp 1
transform 1 0 3220 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0811_
timestamp 1
transform -1 0 2576 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_4  _0812_
timestamp 1
transform -1 0 7912 0 1 12512
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_2  _0813_
timestamp 1
transform 1 0 7360 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0814_
timestamp 1
transform 1 0 3404 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1
transform 1 0 1472 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0816_
timestamp 1
transform 1 0 4968 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1
transform 1 0 5060 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0818_
timestamp 1
transform 1 0 3956 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0819_
timestamp 1
transform -1 0 2852 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0820_
timestamp 1
transform 1 0 8372 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0821_
timestamp 1
transform 1 0 6348 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1
transform -1 0 6348 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0823_
timestamp 1
transform 1 0 3220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0824_
timestamp 1
transform -1 0 2944 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0825_
timestamp 1
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1
transform -1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0827_
timestamp 1
transform -1 0 9108 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0828_
timestamp 1
transform 1 0 9476 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0830_
timestamp 1
transform 1 0 11868 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0831_
timestamp 1
transform 1 0 12696 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0832_
timestamp 1
transform 1 0 14812 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0833_
timestamp 1
transform -1 0 16836 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0834_
timestamp 1
transform 1 0 10948 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0835_
timestamp 1
transform 1 0 13064 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0836_
timestamp 1
transform -1 0 14352 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0837_
timestamp 1
transform 1 0 14076 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0838_
timestamp 1
transform 1 0 16468 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0839_
timestamp 1
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0840_
timestamp 1
transform 1 0 14904 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0841_
timestamp 1
transform -1 0 16008 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1
transform 1 0 15364 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0843_
timestamp 1
transform 1 0 15640 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0844_
timestamp 1
transform -1 0 18216 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0845_
timestamp 1
transform 1 0 16284 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0846_
timestamp 1
transform 1 0 17112 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0847_
timestamp 1
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0848_
timestamp 1
transform -1 0 14996 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_1  _0849_
timestamp 1
transform 1 0 14996 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0850_
timestamp 1
transform -1 0 15088 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0851_
timestamp 1
transform 1 0 14352 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0852_
timestamp 1
transform -1 0 13064 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0853_
timestamp 1
transform 1 0 12328 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _0854_
timestamp 1
transform -1 0 6624 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _0855_
timestamp 1
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0856_
timestamp 1
transform -1 0 19872 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1
transform -1 0 21712 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0858_
timestamp 1
transform 1 0 20424 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0859_
timestamp 1
transform -1 0 21712 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0860_
timestamp 1
transform -1 0 20148 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0861_
timestamp 1
transform 1 0 19780 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0862_
timestamp 1
transform -1 0 19780 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0863_
timestamp 1
transform -1 0 21160 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _0864_
timestamp 1
transform 1 0 20516 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0865_
timestamp 1
transform -1 0 21712 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1
transform 1 0 17940 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0867_
timestamp 1
transform 1 0 18952 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0868_
timestamp 1
transform 1 0 18768 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_2  _0869_
timestamp 1
transform 1 0 8464 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0870_
timestamp 1
transform 1 0 10948 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0871_
timestamp 1
transform 1 0 15272 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0872_
timestamp 1
transform 1 0 11316 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0873_
timestamp 1
transform -1 0 11408 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0874_
timestamp 1
transform 1 0 15916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1
transform -1 0 15456 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0876_
timestamp 1
transform 1 0 14536 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1
transform 1 0 13984 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0878_
timestamp 1
transform 1 0 12328 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0879_
timestamp 1
transform 1 0 12696 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1
transform 1 0 13524 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0881_
timestamp 1
transform 1 0 13340 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0882_
timestamp 1
transform 1 0 13064 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0883_
timestamp 1
transform 1 0 15640 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1
transform 1 0 15548 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0885_
timestamp 1
transform 1 0 11132 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0886_
timestamp 1
transform 1 0 9936 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0887_
timestamp 1
transform 1 0 7820 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0888_
timestamp 1
transform -1 0 10212 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0889_
timestamp 1
transform 1 0 18124 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0890_
timestamp 1
transform -1 0 19412 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1
transform 1 0 19412 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0892_
timestamp 1
transform 1 0 17756 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0893_
timestamp 1
transform 1 0 16652 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0894_
timestamp 1
transform 1 0 18676 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1
transform -1 0 18584 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0896_
timestamp 1
transform -1 0 12604 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0897_
timestamp 1
transform 1 0 18400 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1
transform 1 0 18124 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0899_
timestamp 1
transform 1 0 21620 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1
transform 1 0 18676 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0901_
timestamp 1
transform 1 0 18676 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0902_
timestamp 1
transform 1 0 18032 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0903_
timestamp 1
transform 1 0 15824 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0904_
timestamp 1
transform -1 0 15916 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0905_
timestamp 1
transform -1 0 13340 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _0906_
timestamp 1
transform -1 0 21436 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0908_
timestamp 1
transform 1 0 21252 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1
transform 1 0 20792 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0910_
timestamp 1
transform 1 0 22724 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1
transform 1 0 22448 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0912_
timestamp 1
transform -1 0 22724 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1
transform 1 0 22908 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0914_
timestamp 1
transform -1 0 22264 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0915_
timestamp 1
transform 1 0 21712 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _0916_
timestamp 1
transform 1 0 21160 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0917_
timestamp 1
transform 1 0 9936 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0918_
timestamp 1
transform -1 0 11868 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0919_
timestamp 1
transform -1 0 11408 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1
transform -1 0 9936 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0921_
timestamp 1
transform -1 0 11224 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1
transform 1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1
transform -1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0924_
timestamp 1
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0925_
timestamp 1
transform -1 0 7728 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1
transform 1 0 6164 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1
transform -1 0 4968 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0928_
timestamp 1
transform -1 0 4416 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1
transform -1 0 3680 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1
transform -1 0 13248 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0931_
timestamp 1
transform -1 0 3588 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0932_
timestamp 1
transform -1 0 3128 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1
transform 1 0 4600 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0934_
timestamp 1
transform -1 0 3956 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0935_
timestamp 1
transform 1 0 3956 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0936_
timestamp 1
transform 1 0 5796 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 1
transform 1 0 8004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0938_
timestamp 1
transform -1 0 9016 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0939_
timestamp 1
transform 1 0 7268 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0940_
timestamp 1
transform -1 0 10856 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 1
transform 1 0 17112 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0942_
timestamp 1
transform 1 0 14812 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0943_
timestamp 1
transform 1 0 11776 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1
transform -1 0 10856 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1
transform 1 0 9936 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0946_
timestamp 1
transform -1 0 12052 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0947_
timestamp 1
transform 1 0 10856 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1
transform 1 0 10948 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0949_
timestamp 1
transform 1 0 11132 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0950_
timestamp 1
transform 1 0 10120 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 1
transform 1 0 10488 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0952_
timestamp 1
transform 1 0 12052 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0953_
timestamp 1
transform 1 0 12512 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0954_
timestamp 1
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0955_
timestamp 1
transform 1 0 12696 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0956_
timestamp 1
transform -1 0 16192 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0957_
timestamp 1
transform 1 0 16192 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0958_
timestamp 1
transform -1 0 16008 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0959_
timestamp 1
transform 1 0 15364 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1
transform 1 0 16652 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0961_
timestamp 1
transform -1 0 18216 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0962_
timestamp 1
transform -1 0 18676 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0963_
timestamp 1
transform 1 0 17388 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0964_
timestamp 1
transform 1 0 25484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0965_
timestamp 1
transform -1 0 28060 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1
transform -1 0 29440 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0967_
timestamp 1
transform -1 0 28336 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1
transform 1 0 28428 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0969_
timestamp 1
transform -1 0 27324 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0970_
timestamp 1
transform 1 0 25668 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1
transform -1 0 25668 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0972_
timestamp 1
transform -1 0 22264 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1
transform -1 0 21804 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0974_
timestamp 1
transform -1 0 20976 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0975_
timestamp 1
transform 1 0 20240 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0976_
timestamp 1
transform 1 0 21252 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0977_
timestamp 1
transform -1 0 20608 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0978_
timestamp 1
transform 1 0 22264 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0979_
timestamp 1
transform -1 0 19964 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0980_
timestamp 1
transform -1 0 22632 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 1
transform -1 0 21068 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0982_
timestamp 1
transform 1 0 25208 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0983_
timestamp 1
transform -1 0 24472 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0984_
timestamp 1
transform 1 0 26128 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0985_
timestamp 1
transform -1 0 23736 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0986_
timestamp 1
transform -1 0 26864 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1
transform -1 0 25668 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0988_
timestamp 1
transform -1 0 26864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1
transform -1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0990_
timestamp 1
transform -1 0 27692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0991_
timestamp 1
transform 1 0 28980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0992_
timestamp 1
transform -1 0 29348 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0993_
timestamp 1
transform -1 0 28612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0994_
timestamp 1
transform 1 0 29164 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0995_
timestamp 1
transform 1 0 28612 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0996_
timestamp 1
transform -1 0 30360 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0997_
timestamp 1
transform 1 0 30636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0998_
timestamp 1
transform 1 0 27692 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0999_
timestamp 1
transform -1 0 26220 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1000_
timestamp 1
transform 1 0 28336 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1001_
timestamp 1
transform 1 0 25852 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1002_
timestamp 1
transform 1 0 28520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1003_
timestamp 1
transform 1 0 28888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1004_
timestamp 1
transform 1 0 28060 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1005_
timestamp 1
transform 1 0 16376 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1
transform 1 0 20792 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1007_
timestamp 1
transform -1 0 23092 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1
transform -1 0 23276 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1009_
timestamp 1
transform -1 0 22172 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1010_
timestamp 1
transform 1 0 9568 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1011_
timestamp 1
transform -1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1
transform 1 0 10396 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1013_
timestamp 1
transform 1 0 9476 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1014_
timestamp 1
transform -1 0 11592 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1015_
timestamp 1
transform 1 0 10120 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1
transform -1 0 14904 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1
transform -1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1
transform 1 0 16008 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1019_
timestamp 1
transform -1 0 16928 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1
transform -1 0 15272 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1021_
timestamp 1
transform -1 0 14536 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1
transform 1 0 18124 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _1023_
timestamp 1
transform 1 0 13524 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1
transform 1 0 20424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1025_
timestamp 1
transform -1 0 21160 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1
transform 1 0 9844 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1027_
timestamp 1
transform -1 0 10672 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1028_
timestamp 1
transform 1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1029_
timestamp 1
transform -1 0 16284 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1
transform 1 0 17388 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1
transform 1 0 16652 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 1
transform -1 0 20240 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1033_
timestamp 1
transform 1 0 20332 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1034_
timestamp 1
transform -1 0 23736 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1035_
timestamp 1
transform -1 0 23552 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1
transform -1 0 22540 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1037_
timestamp 1
transform -1 0 21712 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1038_
timestamp 1
transform 1 0 21252 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1
transform 1 0 21252 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1040_
timestamp 1
transform -1 0 24288 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1041_
timestamp 1
transform -1 0 23460 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1
transform 1 0 22448 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1
transform 1 0 22448 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1
transform 1 0 25024 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1
transform -1 0 23736 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1
transform -1 0 24288 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1047_
timestamp 1
transform -1 0 23000 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1
transform -1 0 21712 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1049_
timestamp 1
transform -1 0 20608 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1050_
timestamp 1
transform -1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1051_
timestamp 1
transform -1 0 3772 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1052_
timestamp 1
transform 1 0 4140 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1053_
timestamp 1
transform 1 0 3956 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1
transform 1 0 1840 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1055_
timestamp 1
transform 1 0 3404 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1
transform 1 0 2484 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1057_
timestamp 1
transform 1 0 2208 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1058_
timestamp 1
transform -1 0 4416 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1059_
timestamp 1
transform 1 0 3128 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1060_
timestamp 1
transform 1 0 1932 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1061_
timestamp 1
transform 1 0 1656 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1062_
timestamp 1
transform -1 0 3680 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1063_
timestamp 1
transform 1 0 2392 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1064_
timestamp 1
transform -1 0 1932 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1
transform -1 0 3128 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1
transform 1 0 1932 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1
transform 1 0 2392 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1
transform -1 0 7176 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1069_
timestamp 1
transform 1 0 16008 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1
transform -1 0 17940 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1071_
timestamp 1
transform 1 0 18308 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1072_
timestamp 1
transform 1 0 15732 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1073_
timestamp 1
transform 1 0 12788 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1074_
timestamp 1
transform 1 0 16928 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1075_
timestamp 1
transform 1 0 13524 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1076_
timestamp 1
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1077_
timestamp 1
transform -1 0 19596 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1078_
timestamp 1
transform -1 0 18584 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _1079_
timestamp 1
transform -1 0 17940 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _1080_
timestamp 1
transform 1 0 18400 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1081_
timestamp 1
transform 1 0 17572 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1082_
timestamp 1
transform 1 0 18124 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1083_
timestamp 1
transform 1 0 17020 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1084_
timestamp 1
transform 1 0 16284 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1085_
timestamp 1
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1
transform 1 0 16192 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1087_
timestamp 1
transform 1 0 15548 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1088_
timestamp 1
transform 1 0 15640 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1089_
timestamp 1
transform 1 0 14628 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1090_
timestamp 1
transform -1 0 17480 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1091_
timestamp 1
transform -1 0 15732 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1
transform 1 0 15364 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1093_
timestamp 1
transform 1 0 16100 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1094_
timestamp 1
transform -1 0 15364 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1095_
timestamp 1
transform 1 0 17204 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1096_
timestamp 1
transform 1 0 17204 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1097_
timestamp 1
transform -1 0 16008 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1098_
timestamp 1
transform 1 0 16100 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1
transform 1 0 14720 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1100_
timestamp 1
transform -1 0 16928 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1101_
timestamp 1
transform -1 0 16008 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1102_
timestamp 1
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1103_
timestamp 1
transform 1 0 15180 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1104_
timestamp 1
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1105_
timestamp 1
transform 1 0 25668 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1106_
timestamp 1
transform 1 0 28428 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1
transform 1 0 28888 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1108_
timestamp 1
transform -1 0 30912 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1109_
timestamp 1
transform -1 0 28336 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1110_
timestamp 1
transform -1 0 31280 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 1
transform -1 0 29808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1112_
timestamp 1
transform -1 0 30452 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1113_
timestamp 1
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1
transform 1 0 30084 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1115_
timestamp 1
transform -1 0 28428 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1116_
timestamp 1
transform -1 0 29992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1117_
timestamp 1
transform 1 0 26588 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1118_
timestamp 1
transform 1 0 26312 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1119_
timestamp 1
transform -1 0 26312 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1120_
timestamp 1
transform 1 0 17572 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1121_
timestamp 1
transform 1 0 9016 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1122_
timestamp 1
transform 1 0 10304 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1
transform -1 0 10764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_4  _1124_
timestamp 1
transform 1 0 9384 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1
transform -1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1
transform -1 0 8280 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1127_
timestamp 1
transform 1 0 6256 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1128_
timestamp 1
transform 1 0 5428 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1129_
timestamp 1
transform 1 0 7452 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1130_
timestamp 1
transform 1 0 6624 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 1
transform -1 0 7912 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1132_
timestamp 1
transform 1 0 7636 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1133_
timestamp 1
transform 1 0 7912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1134_
timestamp 1
transform 1 0 7084 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _1135_
timestamp 1
transform 1 0 6624 0 1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1136_
timestamp 1
transform -1 0 8188 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1
transform -1 0 7636 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1138_
timestamp 1
transform 1 0 9016 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1139_
timestamp 1
transform -1 0 6256 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1140_
timestamp 1
transform -1 0 4692 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1141_
timestamp 1
transform 1 0 3220 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 1
transform 1 0 2576 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1
transform 1 0 4324 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1144_
timestamp 1
transform -1 0 4324 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 1
transform -1 0 5520 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1146_
timestamp 1
transform -1 0 5244 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1147_
timestamp 1
transform 1 0 3588 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1148_
timestamp 1
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1149_
timestamp 1
transform -1 0 4416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1150_
timestamp 1
transform 1 0 6440 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1151_
timestamp 1
transform -1 0 10396 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1152_
timestamp 1
transform 1 0 11592 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1153_
timestamp 1
transform 1 0 25300 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1154_
timestamp 1
transform 1 0 24196 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1155_
timestamp 1
transform -1 0 25024 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1156_
timestamp 1
transform 1 0 23184 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1157_
timestamp 1
transform 1 0 24656 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1158_
timestamp 1
transform -1 0 25668 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1159_
timestamp 1
transform 1 0 25116 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1160_
timestamp 1
transform -1 0 26312 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1161_
timestamp 1
transform -1 0 26588 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1162_
timestamp 1
transform 1 0 25300 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1163_
timestamp 1
transform -1 0 26036 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1164_
timestamp 1
transform 1 0 25760 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1165_
timestamp 1
transform -1 0 27508 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1166_
timestamp 1
transform -1 0 28888 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1167_
timestamp 1
transform -1 0 27140 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 1
transform 1 0 11868 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1169_
timestamp 1
transform 1 0 12512 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1170_
timestamp 1
transform -1 0 12604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1171_
timestamp 1
transform 1 0 11684 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1172_
timestamp 1
transform -1 0 11684 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1173_
timestamp 1
transform -1 0 11500 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1174_
timestamp 1
transform 1 0 10396 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1
transform 1 0 6532 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1176_
timestamp 1
transform 1 0 9476 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1177_
timestamp 1
transform 1 0 7452 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1178_
timestamp 1
transform -1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1179_
timestamp 1
transform -1 0 10304 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1180_
timestamp 1
transform -1 0 12972 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1181_
timestamp 1
transform -1 0 13064 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1182_
timestamp 1
transform -1 0 12512 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1183_
timestamp 1
transform -1 0 11776 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1184_
timestamp 1
transform 1 0 9844 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1185_
timestamp 1
transform -1 0 10856 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1186_
timestamp 1
transform -1 0 10212 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1187_
timestamp 1
transform 1 0 9108 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1188_
timestamp 1
transform 1 0 4508 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1189_
timestamp 1
transform -1 0 6440 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 1
transform -1 0 7452 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1191_
timestamp 1
transform -1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1192_
timestamp 1
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1193_
timestamp 1
transform -1 0 10580 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1194_
timestamp 1
transform -1 0 10856 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1195_
timestamp 1
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1196_
timestamp 1
transform 1 0 9936 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1197_
timestamp 1
transform -1 0 4600 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1198_
timestamp 1
transform 1 0 3036 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__nand3_1  _1199_
timestamp 1
transform 1 0 6164 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1200_
timestamp 1
transform -1 0 4692 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1201_
timestamp 1
transform 1 0 6532 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1202_
timestamp 1
transform 1 0 4968 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1203_
timestamp 1
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1204_
timestamp 1
transform -1 0 7636 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1205_
timestamp 1
transform 1 0 8648 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1206_
timestamp 1
transform 1 0 21896 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1207_
timestamp 1
transform 1 0 20056 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1208_
timestamp 1
transform -1 0 22908 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1209_
timestamp 1
transform -1 0 24196 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1210_
timestamp 1
transform 1 0 22264 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1211_
timestamp 1
transform -1 0 23184 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1212_
timestamp 1
transform 1 0 22908 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1213_
timestamp 1
transform -1 0 21436 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1
transform 1 0 20240 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1215_
timestamp 1
transform 1 0 19228 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1216_
timestamp 1
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1217_
timestamp 1
transform -1 0 20792 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1218_
timestamp 1
transform -1 0 22908 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1219_
timestamp 1
transform -1 0 23460 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1
transform 1 0 24012 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1221_
timestamp 1
transform 1 0 23920 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1222_
timestamp 1
transform 1 0 24012 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1223_
timestamp 1
transform 1 0 23736 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1224_
timestamp 1
transform 1 0 23276 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1225_
timestamp 1
transform 1 0 26404 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1226_
timestamp 1
transform 1 0 26404 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1227_
timestamp 1
transform 1 0 25116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1228_
timestamp 1
transform -1 0 25576 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1229_
timestamp 1
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1230_
timestamp 1
transform 1 0 27600 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1231_
timestamp 1
transform 1 0 27876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1232_
timestamp 1
transform 1 0 27140 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1233_
timestamp 1
transform 1 0 26956 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1234_
timestamp 1
transform -1 0 27876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1
transform 1 0 28980 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1236_
timestamp 1
transform -1 0 31188 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp 1
transform 1 0 28888 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1238_
timestamp 1
transform 1 0 28980 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1
transform -1 0 28888 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1
transform 1 0 29900 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1241_
timestamp 1
transform 1 0 28796 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1
transform 1 0 29072 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1243_
timestamp 1
transform -1 0 28796 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1244_
timestamp 1
transform -1 0 31188 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1
transform -1 0 30176 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1246_
timestamp 1
transform -1 0 29716 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1247_
timestamp 1
transform -1 0 30452 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1248_
timestamp 1
transform -1 0 31096 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1249_
timestamp 1
transform -1 0 28152 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1250_
timestamp 1
transform 1 0 27692 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1251_
timestamp 1
transform -1 0 28888 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1252_
timestamp 1
transform 1 0 28888 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1253_
timestamp 1
transform -1 0 28152 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1254_
timestamp 1
transform -1 0 28888 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1255_
timestamp 1
transform 1 0 28980 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1256_
timestamp 1
transform -1 0 28888 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1257_
timestamp 1
transform -1 0 30268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1258_
timestamp 1
transform 1 0 29900 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1
transform -1 0 29808 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1260_
timestamp 1
transform 1 0 27692 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1261_
timestamp 1
transform -1 0 29072 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1262_
timestamp 1
transform -1 0 29900 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1263_
timestamp 1
transform 1 0 29808 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1264_
timestamp 1
transform -1 0 29532 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1265_
timestamp 1
transform 1 0 25852 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1266_
timestamp 1
transform -1 0 27048 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1267_
timestamp 1
transform -1 0 27232 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1268_
timestamp 1
transform 1 0 27232 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1269_
timestamp 1
transform -1 0 27416 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1270_
timestamp 1
transform 1 0 23276 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1271_
timestamp 1
transform -1 0 25300 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1272_
timestamp 1
transform 1 0 24748 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1273_
timestamp 1
transform 1 0 24104 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1
transform -1 0 24564 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1
transform 1 0 24748 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1
transform -1 0 26772 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1277_
timestamp 1
transform -1 0 26036 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1278_
timestamp 1
transform -1 0 26312 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1279_
timestamp 1
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1280_
timestamp 1
transform 1 0 23184 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1281_
timestamp 1
transform 1 0 23000 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1282_
timestamp 1
transform 1 0 23828 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1283_
timestamp 1
transform -1 0 23736 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1284_
timestamp 1
transform -1 0 24564 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1285_
timestamp 1
transform -1 0 21252 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1286_
timestamp 1
transform -1 0 22080 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1287_
timestamp 1
transform -1 0 22724 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1288_
timestamp 1
transform -1 0 23460 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1
transform 1 0 14720 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1290_
timestamp 1
transform 1 0 13892 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _1291_
timestamp 1
transform -1 0 20148 0 1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _1292_
timestamp 1
transform -1 0 17204 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1293_
timestamp 1
transform 1 0 16836 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1294_
timestamp 1
transform -1 0 16560 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1295_
timestamp 1
transform -1 0 16008 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1296_
timestamp 1
transform -1 0 16928 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1297_
timestamp 1
transform 1 0 17112 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1298_
timestamp 1
transform 1 0 18400 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1299_
timestamp 1
transform 1 0 19412 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1300_
timestamp 1
transform 1 0 18676 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1301_
timestamp 1
transform -1 0 19228 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1302_
timestamp 1
transform 1 0 20424 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1303_
timestamp 1
transform 1 0 17848 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1304_
timestamp 1
transform -1 0 26588 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1305_
timestamp 1
transform -1 0 23184 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1306_
timestamp 1
transform -1 0 11684 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1307_
timestamp 1
transform 1 0 11040 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1308_
timestamp 1
transform 1 0 11316 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1309__3
timestamp 1
transform 1 0 18124 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1310__4
timestamp 1
transform -1 0 19872 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1311__5
timestamp 1
transform 1 0 16928 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1312__6
timestamp 1
transform -1 0 15732 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1313__7
timestamp 1
transform -1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1314__8
timestamp 1
transform -1 0 23736 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1315__9
timestamp 1
transform -1 0 24564 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1316__10
timestamp 1
transform 1 0 24840 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1317__11
timestamp 1
transform 1 0 24380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1318__12
timestamp 1
transform -1 0 27784 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1319__13
timestamp 1
transform 1 0 28980 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1320__14
timestamp 1
transform 1 0 29256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1321__15
timestamp 1
transform 1 0 30452 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1322__16
timestamp 1
transform -1 0 29256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1323__17
timestamp 1
transform 1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1324__18
timestamp 1
transform 1 0 31004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1325__19
timestamp 1
transform 1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1326__20
timestamp 1
transform -1 0 26220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1327__21
timestamp 1
transform 1 0 24748 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1328__22
timestamp 1
transform 1 0 18676 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1329__23
timestamp 1
transform 1 0 8004 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1330__24
timestamp 1
transform -1 0 11776 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1331__25
timestamp 1
transform 1 0 8372 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1332__26
timestamp 1
transform -1 0 9936 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1333__27
timestamp 1
transform 1 0 13156 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1334__28
timestamp 1
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1335__29
timestamp 1
transform -1 0 12696 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1336__30
timestamp 1
transform -1 0 5612 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1337__31
timestamp 1
transform -1 0 2852 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1338__32
timestamp 1
transform -1 0 3128 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339__33
timestamp 1
transform -1 0 6256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1340__34
timestamp 1
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1341__35
timestamp 1
transform -1 0 4692 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1342__36
timestamp 1
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1343__37
timestamp 1
transform -1 0 19044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1344__38
timestamp 1
transform 1 0 25484 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1345__39
timestamp 1
transform -1 0 27784 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1346__40
timestamp 1
transform -1 0 29256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1347__41
timestamp 1
transform -1 0 31096 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1348__42
timestamp 1
transform 1 0 29808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1349__43
timestamp 1
transform -1 0 29532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1350__44
timestamp 1
transform 1 0 27140 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1351__45
timestamp 1
transform -1 0 13892 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1352__46
timestamp 1
transform -1 0 15824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1353__47
timestamp 1
transform 1 0 13156 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1354__48
timestamp 1
transform 1 0 13616 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1355__49
timestamp 1
transform 1 0 6072 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1356__50
timestamp 1
transform -1 0 1472 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1357__51
timestamp 1
transform 1 0 4140 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1358__52
timestamp 1
transform -1 0 2300 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1359__53
timestamp 1
transform -1 0 4048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1360__54
timestamp 1
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1361__55
timestamp 1
transform -1 0 2024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1362__56
timestamp 1
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1363__57
timestamp 1
transform 1 0 1564 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1364__58
timestamp 1
transform -1 0 20976 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1365__59
timestamp 1
transform -1 0 22264 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1366__60
timestamp 1
transform -1 0 25760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1367__61
timestamp 1
transform 1 0 22172 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1368__62
timestamp 1
transform -1 0 23828 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1369__63
timestamp 1
transform 1 0 20424 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1370__64
timestamp 1
transform -1 0 22080 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1371__65
timestamp 1
transform -1 0 24196 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1372__66
timestamp 1
transform -1 0 17204 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1373__67
timestamp 1
transform 1 0 17020 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1374__68
timestamp 1
transform -1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1375__69
timestamp 1
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1376__70
timestamp 1
transform -1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1377__71
timestamp 1
transform -1 0 15916 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1378__72
timestamp 1
transform 1 0 16928 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1379__73
timestamp 1
transform -1 0 14720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1380__74
timestamp 1
transform -1 0 22448 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1381__75
timestamp 1
transform -1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1382__76
timestamp 1
transform 1 0 30360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1383__77
timestamp 1
transform -1 0 26772 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1384__78
timestamp 1
transform 1 0 24932 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1385__79
timestamp 1
transform 1 0 30912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1386__80
timestamp 1
transform 1 0 28612 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1387__81
timestamp 1
transform 1 0 28060 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1388__82
timestamp 1
transform -1 0 29532 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1389__83
timestamp 1
transform 1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1390__84
timestamp 1
transform 1 0 24012 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1391__85
timestamp 1
transform -1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1392__86
timestamp 1
transform -1 0 24104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1393__87
timestamp 1
transform 1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1394__88
timestamp 1
transform 1 0 19320 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1395__89
timestamp 1
transform -1 0 20056 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1396__90
timestamp 1
transform 1 0 19228 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1397__91
timestamp 1
transform 1 0 18308 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1398__92
timestamp 1
transform -1 0 18492 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1399__93
timestamp 1
transform -1 0 16560 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1400__94
timestamp 1
transform -1 0 16376 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1401__95
timestamp 1
transform -1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1402__96
timestamp 1
transform 1 0 13156 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1403__97
timestamp 1
transform -1 0 9660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1404__98
timestamp 1
transform -1 0 12512 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1405__99
timestamp 1
transform -1 0 9384 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1406__100
timestamp 1
transform -1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1407__101
timestamp 1
transform 1 0 6256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1408__102
timestamp 1
transform 1 0 6532 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1409__103
timestamp 1
transform -1 0 5704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1410__104
timestamp 1
transform -1 0 3956 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1411__105
timestamp 1
transform -1 0 3496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1412__106
timestamp 1
transform -1 0 2024 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1413__107
timestamp 1
transform -1 0 22632 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1414__108
timestamp 1
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1415__109
timestamp 1
transform -1 0 23736 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1416__110
timestamp 1
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1417__111
timestamp 1
transform -1 0 16468 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1418__112
timestamp 1
transform -1 0 20700 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1419__113
timestamp 1
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1420__114
timestamp 1
transform -1 0 19044 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1421__115
timestamp 1
transform -1 0 13340 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1422__116
timestamp 1
transform -1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1423__117
timestamp 1
transform -1 0 17480 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1424__118
timestamp 1
transform -1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1425__119
timestamp 1
transform -1 0 10764 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1426__120
timestamp 1
transform -1 0 16652 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1427__121
timestamp 1
transform 1 0 14996 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1428__122
timestamp 1
transform 1 0 13156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1429__123
timestamp 1
transform -1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1430__124
timestamp 1
transform 1 0 13708 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1431__125
timestamp 1
transform 1 0 14628 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1432__126
timestamp 1
transform 1 0 10212 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1433__127
timestamp 1
transform -1 0 19228 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1434__128
timestamp 1
transform -1 0 12236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1435__129
timestamp 1
transform -1 0 10304 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1436__130
timestamp 1
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1437__131
timestamp 1
transform 1 0 2024 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1438__132
timestamp 1
transform 1 0 5520 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1439__133
timestamp 1
transform -1 0 7912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1440__134
timestamp 1
transform -1 0 1656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1441__135
timestamp 1
transform -1 0 6164 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1442__136
timestamp 1
transform -1 0 2300 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1443__137
timestamp 1
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1444__138
timestamp 1
transform -1 0 2944 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1445__139
timestamp 1
transform -1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1446__140
timestamp 1
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1447__141
timestamp 1
transform 1 0 5244 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1448__142
timestamp 1
transform -1 0 2024 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1449__143
timestamp 1
transform 1 0 1656 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1450__144
timestamp 1
transform -1 0 2300 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1
transform 1 0 10580 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1
transform 1 0 18676 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1
transform 1 0 18676 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1
transform -1 0 17848 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1
transform 1 0 15364 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1
transform 1 0 12420 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1
transform -1 0 22724 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1
transform 1 0 24196 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1
transform 1 0 24748 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1
transform 1 0 24564 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1461_
timestamp 1
transform 1 0 27416 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1
transform 1 0 29532 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1
transform 1 0 29532 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1
transform -1 0 30728 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1
transform 1 0 28152 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1
transform 1 0 29532 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1
transform -1 0 30636 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1
transform 1 0 27140 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1
transform 1 0 25300 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1
transform 1 0 23828 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1471_
timestamp 1
transform 1 0 18952 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1472_
timestamp 1
transform 1 0 8740 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1473_
timestamp 1
transform -1 0 11500 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1474_
timestamp 1
transform 1 0 8924 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1475_
timestamp 1
transform -1 0 22724 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1476_
timestamp 1
transform -1 0 30820 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1477_
timestamp 1
transform -1 0 29348 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1478_
timestamp 1
transform -1 0 27968 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1479_
timestamp 1
transform -1 0 27876 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1480_
timestamp 1
transform -1 0 27324 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1481_
timestamp 1
transform -1 0 25852 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1482_
timestamp 1
transform -1 0 25668 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1483_
timestamp 1
transform -1 0 24196 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1484_
timestamp 1
transform 1 0 9936 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1485_
timestamp 1
transform 1 0 13524 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1486_
timestamp 1
transform 1 0 7268 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1487_
timestamp 1
transform -1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1488_
timestamp 1
transform 1 0 5244 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1489_
timestamp 1
transform 1 0 2484 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1490_
timestamp 1
transform -1 0 2484 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1491_
timestamp 1
transform 1 0 5980 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1492_
timestamp 1
transform 1 0 6256 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1493_
timestamp 1
transform 1 0 4140 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1494_
timestamp 1
transform 1 0 4232 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1495_
timestamp 1
transform 1 0 18676 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1496_
timestamp 1
transform 1 0 25760 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1497_
timestamp 1
transform 1 0 27416 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1498_
timestamp 1
transform -1 0 30360 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1499_
timestamp 1
transform -1 0 30820 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1500_
timestamp 1
transform -1 0 30636 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1501_
timestamp 1
transform 1 0 29164 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1502_
timestamp 1
transform 1 0 27416 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1503_
timestamp 1
transform 1 0 13524 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1504_
timestamp 1
transform 1 0 15456 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1505_
timestamp 1
transform 1 0 13340 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1506_
timestamp 1
transform 1 0 13892 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1507_
timestamp 1
transform 1 0 6532 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1508_
timestamp 1
transform 1 0 1932 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1509_
timestamp 1
transform -1 0 4692 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1510_
timestamp 1
transform 1 0 1932 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1511_
timestamp 1
transform 1 0 3404 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1512_
timestamp 1
transform 1 0 1656 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1513_
timestamp 1
transform 1 0 1656 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1514_
timestamp 1
transform 1 0 1656 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1515_
timestamp 1
transform 1 0 1932 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1516_
timestamp 1
transform 1 0 20608 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1517_
timestamp 1
transform 1 0 22724 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1518_
timestamp 1
transform 1 0 24196 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1519_
timestamp 1
transform 1 0 22080 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1520_
timestamp 1
transform 1 0 23460 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1521_
timestamp 1
transform 1 0 20700 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1522_
timestamp 1
transform 1 0 21712 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1
transform 1 0 23828 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1
transform 1 0 16836 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1
transform 1 0 16560 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1
transform -1 0 11684 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1
transform 1 0 21252 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1
transform 1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1
transform 1 0 14536 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1530_
timestamp 1
transform 1 0 16468 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1
transform 1 0 13984 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1
transform 1 0 21252 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1
transform 1 0 28612 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1534_
timestamp 1
transform -1 0 30544 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1535_
timestamp 1
transform 1 0 26404 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1536_
timestamp 1
transform 1 0 25208 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1537_
timestamp 1
transform -1 0 30912 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1538_
timestamp 1
transform 1 0 29256 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1539_
timestamp 1
transform -1 0 28980 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1540_
timestamp 1
transform -1 0 28796 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1541_
timestamp 1
transform -1 0 28520 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1542_
timestamp 1
transform 1 0 24288 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1543_
timestamp 1
transform 1 0 23920 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1544_
timestamp 1
transform 1 0 23736 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1545_
timestamp 1
transform 1 0 21252 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1546_
timestamp 1
transform 1 0 19688 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1547_
timestamp 1
transform 1 0 19688 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1548_
timestamp 1
transform 1 0 19504 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1549_
timestamp 1
transform 1 0 18676 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1550_
timestamp 1
transform -1 0 17940 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1551_
timestamp 1
transform 1 0 16192 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1552_
timestamp 1
transform 1 0 16008 0 1 1632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1553_
timestamp 1
transform 1 0 13340 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1554_
timestamp 1
transform 1 0 13340 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1555_
timestamp 1
transform 1 0 9292 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1556_
timestamp 1
transform 1 0 11868 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1557_
timestamp 1
transform 1 0 9384 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1558_
timestamp 1
transform 1 0 10948 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1559_
timestamp 1
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1560_
timestamp 1
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1561_
timestamp 1
transform 1 0 5336 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1562_
timestamp 1
transform 1 0 3680 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1563_
timestamp 1
transform 1 0 3128 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1564_
timestamp 1
transform 1 0 1656 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1565_
timestamp 1
transform 1 0 22172 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1566_
timestamp 1
transform 1 0 23828 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1567_
timestamp 1
transform 1 0 23000 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1568_
timestamp 1
transform 1 0 21252 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1569_
timestamp 1
transform 1 0 16100 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1570_
timestamp 1
transform -1 0 19964 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1571_
timestamp 1
transform 1 0 19136 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1572_
timestamp 1
transform 1 0 18676 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1573_
timestamp 1
transform 1 0 12604 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1574_
timestamp 1
transform 1 0 17940 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1575_
timestamp 1
transform 1 0 17112 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1576_
timestamp 1
transform -1 0 20884 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1577_
timestamp 1
transform 1 0 10396 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1578_
timestamp 1
transform 1 0 16100 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1579_
timestamp 1
transform -1 0 14996 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1580_
timestamp 1
transform 1 0 13524 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1
transform 1 0 11960 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1
transform 1 0 14444 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1
transform 1 0 14536 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1
transform 1 0 10488 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1
transform 1 0 18860 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1
transform 1 0 11868 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1
transform -1 0 10120 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1
transform 1 0 8372 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1
transform 1 0 2300 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1
transform 1 0 5796 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1
transform 1 0 7176 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1
transform 1 0 1656 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1
transform 1 0 1932 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1
transform 1 0 1656 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1
transform 1 0 2576 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1
transform 1 0 1104 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1
transform 1 0 1656 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1
transform 1 0 5520 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1
transform 1 0 1656 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1
transform 1 0 2024 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1
transform 1 0 1932 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1609_
timestamp 1
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1610_
timestamp 1
transform 1 0 8280 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1611_
timestamp 1
transform 1 0 8372 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1612_
timestamp 1
transform -1 0 6532 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1613_
timestamp 1
transform -1 0 6716 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1614_
timestamp 1
transform 1 0 12788 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1615_
timestamp 1
transform 1 0 12236 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1616_
timestamp 1
transform 1 0 11132 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1617_
timestamp 1
transform -1 0 12236 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1618_
timestamp 1
transform -1 0 10580 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 18124 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1
transform -1 0 6808 0 -1 9248
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1
transform -1 0 5704 0 -1 9248
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1
transform -1 0 11868 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1
transform 1 0 11592 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1
transform 1 0 6256 0 -1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1
transform -1 0 7452 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1
transform 1 0 12880 0 -1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1
transform -1 0 14536 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1
transform -1 0 20424 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1
transform 1 0 20608 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1
transform 1 0 26680 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1
transform 1 0 26404 0 -1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1
transform 1 0 21436 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1
transform 1 0 21252 0 -1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1
transform 1 0 26588 0 1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1
transform 1 0 26404 0 -1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  clkload0
timestamp 1
transform 1 0 5244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  clkload1
timestamp 1
transform 1 0 11040 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  clkload2
timestamp 1
transform 1 0 11592 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload3
timestamp 1
transform 1 0 7268 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload4
timestamp 1
transform -1 0 12880 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  clkload5
timestamp 1
transform 1 0 12972 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  clkload6
timestamp 1
transform -1 0 20424 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkload7
timestamp 1
transform 1 0 24656 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  clkload8
timestamp 1
transform 1 0 25300 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  clkload9
timestamp 1
transform -1 0 22264 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  clkload10
timestamp 1
transform 1 0 22264 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  clkload11
timestamp 1
transform 1 0 27600 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  clkload12
timestamp 1
transform 1 0 25668 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1
transform 1 0 13616 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout12
timestamp 1
transform 1 0 13524 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 1
transform -1 0 22908 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1
transform -1 0 21252 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1
transform -1 0 21160 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout16
timestamp 1
transform 1 0 26036 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1
transform 1 0 10304 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1
transform 1 0 25116 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1
transform -1 0 20516 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1
transform -1 0 23736 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1
transform -1 0 17388 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1
transform -1 0 24748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1
transform 1 0 22080 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1
transform 1 0 22724 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1
transform 1 0 20148 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1
transform -1 0 7636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1
transform -1 0 12328 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1
transform 1 0 18952 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1
transform -1 0 18860 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1
transform 1 0 13616 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1
transform 1 0 21712 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1
transform -1 0 14444 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1
transform 1 0 18216 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 1
transform 1 0 17848 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1
transform 1 0 16192 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1
transform 1 0 16560 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1
transform -1 0 21252 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout40
timestamp 1
transform -1 0 23276 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1
transform -1 0 21804 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1
transform -1 0 13524 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1
transform 1 0 13064 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 1
transform 1 0 10948 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1
transform -1 0 17020 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1
transform 1 0 16928 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1
transform -1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1
transform -1 0 12052 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout49
timestamp 1
transform -1 0 9384 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout50
timestamp 1
transform -1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout51
timestamp 1
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1
transform -1 0 6164 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 1
transform -1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 1
transform -1 0 17756 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 1
transform -1 0 19688 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 1
transform -1 0 22540 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp 1
transform -1 0 26772 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 1
transform 1 0 21804 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1
transform 1 0 30452 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1
transform 1 0 27784 0 -1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_97
timestamp 1
transform 1 0 9476 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_103
timestamp 1
transform 1 0 10028 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_118
timestamp 1636968456
transform 1 0 11408 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_130
timestamp 1
transform 1 0 12512 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1
transform 1 0 13248 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636968456
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636968456
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636968456
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_209
timestamp 1
transform 1 0 19780 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_217
timestamp 1
transform 1 0 20516 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1
transform 1 0 21068 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1
transform 1 0 23828 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_274
timestamp 1
transform 1 0 25760 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636968456
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636968456
transform 1 0 30084 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333
timestamp 1
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_93
timestamp 1
transform 1 0 9108 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1
transform 1 0 10948 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_122
timestamp 1
transform 1 0 11776 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_155
timestamp 1636968456
transform 1 0 14812 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_172
timestamp 1
transform 1 0 16376 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_189
timestamp 1636968456
transform 1 0 17940 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_201
timestamp 1
transform 1 0 19044 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_207
timestamp 1
transform 1 0 19596 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_241
timestamp 1
transform 1 0 22724 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_248
timestamp 1
transform 1 0 23368 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_295
timestamp 1636968456
transform 1 0 27692 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_307
timestamp 1636968456
transform 1 0 28796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_319
timestamp 1636968456
transform 1 0 29900 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_331
timestamp 1
transform 1 0 31004 0 -1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1
transform 1 0 8372 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_151
timestamp 1
transform 1 0 14444 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_160
timestamp 1
transform 1 0 15272 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_197
timestamp 1
transform 1 0 18676 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_203
timestamp 1
transform 1 0 19228 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_286
timestamp 1
transform 1 0 26864 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_304
timestamp 1
transform 1 0 28520 0 1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636968456
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636968456
transform 1 0 30084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 1
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_93
timestamp 1
transform 1 0 9108 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_118
timestamp 1
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_130
timestamp 1
transform 1 0 12512 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_161
timestamp 1
transform 1 0 15364 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 1
transform 1 0 16100 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_194
timestamp 1636968456
transform 1 0 18400 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_206
timestamp 1
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_235
timestamp 1
transform 1 0 22172 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_240
timestamp 1636968456
transform 1 0 22632 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_275
timestamp 1
transform 1 0 25852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_281
timestamp 1
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_307
timestamp 1636968456
transform 1 0 28796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_319
timestamp 1636968456
transform 1 0 29900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_331
timestamp 1
transform 1 0 31004 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1
transform 1 0 5428 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_61
timestamp 1
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_97
timestamp 1
transform 1 0 9476 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_101
timestamp 1
transform 1 0 9844 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_123
timestamp 1636968456
transform 1 0 11868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_135
timestamp 1
transform 1 0 12972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_149
timestamp 1636968456
transform 1 0 14260 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_161
timestamp 1
transform 1 0 15364 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_165
timestamp 1
transform 1 0 15732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_174
timestamp 1
transform 1 0 16560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp 1
transform 1 0 17572 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1
transform 1 0 18308 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_197
timestamp 1
transform 1 0 18676 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_243
timestamp 1
transform 1 0 22908 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_256
timestamp 1
transform 1 0 24104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_280
timestamp 1
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_315
timestamp 1636968456
transform 1 0 29532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_327
timestamp 1
transform 1 0 30636 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_27
timestamp 1
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_33
timestamp 1
transform 1 0 3588 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_48
timestamp 1
transform 1 0 4968 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_52
timestamp 1
transform 1 0 5336 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_90
timestamp 1
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_98
timestamp 1
transform 1 0 9568 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_129
timestamp 1636968456
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_141
timestamp 1636968456
transform 1 0 13524 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_153
timestamp 1636968456
transform 1 0 14628 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1
transform 1 0 15732 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_174
timestamp 1636968456
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_186
timestamp 1636968456
transform 1 0 17664 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_198
timestamp 1
transform 1 0 18768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_206
timestamp 1
transform 1 0 19504 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_212
timestamp 1
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_233
timestamp 1636968456
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_245
timestamp 1636968456
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_257
timestamp 1636968456
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_269
timestamp 1
transform 1 0 25300 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_277
timestamp 1
transform 1 0 26036 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636968456
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_313
timestamp 1636968456
transform 1 0 29348 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_325
timestamp 1
transform 1 0 30452 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_333
timestamp 1
transform 1 0 31188 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_15
timestamp 1
transform 1 0 1932 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_50
timestamp 1
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_92
timestamp 1636968456
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_104
timestamp 1
transform 1 0 10120 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_112
timestamp 1
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 1636968456
transform 1 0 11316 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1
transform 1 0 12420 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_157
timestamp 1636968456
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_169
timestamp 1
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_178
timestamp 1
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_182
timestamp 1
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_190
timestamp 1
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_213
timestamp 1
transform 1 0 20148 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_221
timestamp 1
transform 1 0 20884 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_241
timestamp 1
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_275
timestamp 1
transform 1 0 25852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_299
timestamp 1
transform 1 0 28060 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 1
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1
transform 1 0 828 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_11
timestamp 1
transform 1 0 1564 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_50
timestamp 1
transform 1 0 5152 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_64
timestamp 1
transform 1 0 6440 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_70
timestamp 1
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_78
timestamp 1
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_82
timestamp 1636968456
transform 1 0 8096 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_94
timestamp 1636968456
transform 1 0 9200 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_106
timestamp 1
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_116
timestamp 1636968456
transform 1 0 11224 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_128
timestamp 1
transform 1 0 12328 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_157
timestamp 1
transform 1 0 14996 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_197
timestamp 1
transform 1 0 18676 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_201
timestamp 1636968456
transform 1 0 19044 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_213
timestamp 1
transform 1 0 20148 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_241
timestamp 1
transform 1 0 22724 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_260
timestamp 1
transform 1 0 24472 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_268
timestamp 1
transform 1 0 25208 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 1
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_293
timestamp 1
transform 1 0 27508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_328
timestamp 1
transform 1 0 30728 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_334
timestamp 1
transform 1 0 31280 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 1
transform 1 0 828 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1
transform 1 0 3220 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_42
timestamp 1636968456
transform 1 0 4416 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_54
timestamp 1636968456
transform 1 0 5520 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_66
timestamp 1
transform 1 0 6624 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_74
timestamp 1
transform 1 0 7360 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_92
timestamp 1
transform 1 0 9016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_98
timestamp 1
transform 1 0 9568 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_123
timestamp 1
transform 1 0 11868 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_131
timestamp 1
transform 1 0 12604 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_146
timestamp 1
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_160
timestamp 1
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_175
timestamp 1
transform 1 0 16652 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_179
timestamp 1
transform 1 0 17020 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_183
timestamp 1
transform 1 0 17388 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_213
timestamp 1
transform 1 0 20148 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_219
timestamp 1
transform 1 0 20700 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636968456
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_265
timestamp 1
transform 1 0 24932 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_269
timestamp 1
transform 1 0 25300 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_291
timestamp 1
transform 1 0 27324 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_302
timestamp 1
transform 1 0 28336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_309
timestamp 1
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_317
timestamp 1
transform 1 0 29716 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_331
timestamp 1
transform 1 0 31004 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1
transform 1 0 828 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_11
timestamp 1
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_21
timestamp 1
transform 1 0 2484 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_32
timestamp 1636968456
transform 1 0 3496 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_44
timestamp 1636968456
transform 1 0 4600 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636968456
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1636968456
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_81
timestamp 1
transform 1 0 8004 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_101
timestamp 1
transform 1 0 9844 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_130
timestamp 1
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_160
timestamp 1
transform 1 0 15272 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636968456
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1636968456
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_193
timestamp 1
transform 1 0 18308 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_202
timestamp 1636968456
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_214
timestamp 1
transform 1 0 20240 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1
transform 1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_229
timestamp 1
transform 1 0 21620 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_237
timestamp 1
transform 1 0 22356 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_248
timestamp 1636968456
transform 1 0 23368 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_260
timestamp 1
transform 1 0 24472 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_268
timestamp 1
transform 1 0 25208 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_299
timestamp 1
transform 1 0 28060 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_303
timestamp 1
transform 1 0 28428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_327
timestamp 1
transform 1 0 30636 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_37
timestamp 1636968456
transform 1 0 3956 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_49
timestamp 1636968456
transform 1 0 5060 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_70
timestamp 1
transform 1 0 6992 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 1
transform 1 0 7820 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_93
timestamp 1
transform 1 0 9108 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_107
timestamp 1636968456
transform 1 0 10396 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_119
timestamp 1
transform 1 0 11500 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_128
timestamp 1636968456
transform 1 0 12328 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636968456
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1636968456
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1636968456
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1636968456
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_216
timestamp 1636968456
transform 1 0 20424 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_236
timestamp 1636968456
transform 1 0 22264 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_248
timestamp 1
transform 1 0 23368 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_253
timestamp 1
transform 1 0 23828 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_261
timestamp 1
transform 1 0 24564 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_309
timestamp 1
transform 1 0 28980 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_326
timestamp 1
transform 1 0 30544 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_334
timestamp 1
transform 1 0 31280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 1
transform 1 0 828 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_46
timestamp 1
transform 1 0 4784 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1
transform 1 0 5796 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_71
timestamp 1
transform 1 0 7084 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_86
timestamp 1
transform 1 0 8464 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_107
timestamp 1
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1
transform 1 0 10948 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_119
timestamp 1
transform 1 0 11500 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_123
timestamp 1
transform 1 0 11868 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_127
timestamp 1
transform 1 0 12236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_134
timestamp 1
transform 1 0 12880 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_150
timestamp 1
transform 1 0 14352 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_156
timestamp 1
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_177
timestamp 1
transform 1 0 16836 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_185
timestamp 1
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1
transform 1 0 20976 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_229
timestamp 1
transform 1 0 21620 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_252
timestamp 1636968456
transform 1 0 23736 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_264
timestamp 1
transform 1 0 24840 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_270
timestamp 1
transform 1 0 25392 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_297
timestamp 1
transform 1 0 27876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1
transform 1 0 30820 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_3
timestamp 1
transform 1 0 828 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1
transform 1 0 3956 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_47
timestamp 1
transform 1 0 4876 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_55
timestamp 1
transform 1 0 5612 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_67
timestamp 1
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_71
timestamp 1
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_184
timestamp 1
transform 1 0 17480 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_192
timestamp 1
transform 1 0 18216 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_240
timestamp 1636968456
transform 1 0 22632 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636968456
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1636968456
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_280
timestamp 1
transform 1 0 26312 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_285
timestamp 1636968456
transform 1 0 26772 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_297
timestamp 1
transform 1 0 27876 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_305
timestamp 1
transform 1 0 28612 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_312
timestamp 1636968456
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_324
timestamp 1
transform 1 0 30360 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_332
timestamp 1
transform 1 0 31096 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_15
timestamp 1
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_22
timestamp 1
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_26
timestamp 1636968456
transform 1 0 2944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_38
timestamp 1
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_42
timestamp 1
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp 1
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_61
timestamp 1
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_82
timestamp 1
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_93
timestamp 1
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_131
timestamp 1
transform 1 0 12604 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_152
timestamp 1
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_169
timestamp 1
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_177
timestamp 1636968456
transform 1 0 16836 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_189
timestamp 1
transform 1 0 17940 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1636968456
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_237
timestamp 1
transform 1 0 22356 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_281
timestamp 1
transform 1 0 26404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_290
timestamp 1
transform 1 0 27232 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_296
timestamp 1636968456
transform 1 0 27784 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_308
timestamp 1636968456
transform 1 0 28888 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_320
timestamp 1636968456
transform 1 0 29992 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_332
timestamp 1
transform 1 0 31096 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_15
timestamp 1
transform 1 0 1932 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_24
timestamp 1
transform 1 0 2760 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636968456
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_41
timestamp 1
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_48
timestamp 1
transform 1 0 4968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_54
timestamp 1
transform 1 0 5520 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_64
timestamp 1
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_73
timestamp 1
transform 1 0 7268 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_80
timestamp 1
transform 1 0 7912 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_96
timestamp 1636968456
transform 1 0 9384 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_108
timestamp 1636968456
transform 1 0 10488 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_127
timestamp 1636968456
transform 1 0 12236 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 1
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_150
timestamp 1636968456
transform 1 0 14352 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_162
timestamp 1
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_168
timestamp 1636968456
transform 1 0 16008 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_180
timestamp 1
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_188
timestamp 1
transform 1 0 17848 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_210
timestamp 1
transform 1 0 19872 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_218
timestamp 1
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_223
timestamp 1
transform 1 0 21068 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_231
timestamp 1
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_258
timestamp 1
transform 1 0 24288 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_290
timestamp 1
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_320
timestamp 1636968456
transform 1 0 29992 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_332
timestamp 1
transform 1 0 31096 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1
transform 1 0 828 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_11
timestamp 1
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_40
timestamp 1
transform 1 0 4232 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_44
timestamp 1
transform 1 0 4600 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_68
timestamp 1
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_78
timestamp 1636968456
transform 1 0 7728 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_90
timestamp 1
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_94
timestamp 1
transform 1 0 9200 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_98
timestamp 1
transform 1 0 9568 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1
transform 1 0 10948 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_128
timestamp 1636968456
transform 1 0 12328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_140
timestamp 1
transform 1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_151
timestamp 1
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1
transform 1 0 15732 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1636968456
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_184
timestamp 1
transform 1 0 17480 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_188
timestamp 1
transform 1 0 17848 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1636968456
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_217
timestamp 1
transform 1 0 20516 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1
transform 1 0 20976 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_251
timestamp 1
transform 1 0 23644 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_260
timestamp 1
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_270
timestamp 1
transform 1 0 25392 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_288
timestamp 1
transform 1 0 27048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_296
timestamp 1
transform 1 0 27784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_305
timestamp 1
transform 1 0 28612 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_324
timestamp 1
transform 1 0 30360 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_332
timestamp 1
transform 1 0 31096 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1
transform 1 0 828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_42
timestamp 1
transform 1 0 4416 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_50
timestamp 1
transform 1 0 5152 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_70
timestamp 1
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1
transform 1 0 7912 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_99
timestamp 1
transform 1 0 9660 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_149
timestamp 1
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_200
timestamp 1
transform 1 0 18952 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_208
timestamp 1
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1
transform 1 0 23552 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1
transform 1 0 23828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_262
timestamp 1
transform 1 0 24656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_293
timestamp 1
transform 1 0 27508 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_312
timestamp 1
transform 1 0 29256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_324
timestamp 1
transform 1 0 30360 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_332
timestamp 1
transform 1 0 31096 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1
transform 1 0 828 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_11
timestamp 1
transform 1 0 1564 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1636968456
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1
transform 1 0 5796 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_71
timestamp 1
transform 1 0 7084 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_104
timestamp 1
transform 1 0 10120 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_147
timestamp 1
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_151
timestamp 1
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1636968456
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_181
timestamp 1
transform 1 0 17204 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_195
timestamp 1
transform 1 0 18492 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_201
timestamp 1636968456
transform 1 0 19044 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_213
timestamp 1
transform 1 0 20148 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_221
timestamp 1
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_233
timestamp 1
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_243
timestamp 1636968456
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_255
timestamp 1636968456
transform 1 0 24012 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_284
timestamp 1
transform 1 0 26680 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_288
timestamp 1636968456
transform 1 0 27048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_300
timestamp 1
transform 1 0 28152 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_304
timestamp 1
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_332
timestamp 1
transform 1 0 31096 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636968456
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_15
timestamp 1
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_19
timestamp 1
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1636968456
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_41
timestamp 1
transform 1 0 4324 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_80
timestamp 1
transform 1 0 7912 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_102
timestamp 1
transform 1 0 9936 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_106
timestamp 1636968456
transform 1 0 10304 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_118
timestamp 1
transform 1 0 11408 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_149
timestamp 1
transform 1 0 14260 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_156
timestamp 1
transform 1 0 14904 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_162
timestamp 1
transform 1 0 15456 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1636968456
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_189
timestamp 1
transform 1 0 17940 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_213
timestamp 1
transform 1 0 20148 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_235
timestamp 1
transform 1 0 22172 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1
transform 1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_258
timestamp 1
transform 1 0 24288 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_266
timestamp 1
transform 1 0 25024 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_283
timestamp 1636968456
transform 1 0 26588 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_295
timestamp 1636968456
transform 1 0 27692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_309
timestamp 1
transform 1 0 28980 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_334
timestamp 1
transform 1 0 31280 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636968456
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 1
transform 1 0 1932 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_35
timestamp 1636968456
transform 1 0 3772 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_47
timestamp 1
transform 1 0 4876 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_73
timestamp 1636968456
transform 1 0 7268 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_96
timestamp 1
transform 1 0 9384 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_107
timestamp 1
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_122
timestamp 1636968456
transform 1 0 11776 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_134
timestamp 1636968456
transform 1 0 12880 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_146
timestamp 1636968456
transform 1 0 13984 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_158
timestamp 1
transform 1 0 15088 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_192
timestamp 1
transform 1 0 18216 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_208
timestamp 1636968456
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 1
transform 1 0 20792 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_230
timestamp 1
transform 1 0 21712 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_239
timestamp 1
transform 1 0 22540 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_265
timestamp 1
transform 1 0 24932 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_277
timestamp 1
transform 1 0 26036 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1636968456
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_293
timestamp 1
transform 1 0 27508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 1
transform 1 0 828 0 1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_45
timestamp 1636968456
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_57
timestamp 1
transform 1 0 5796 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_61
timestamp 1
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_67
timestamp 1
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_79
timestamp 1
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_101
timestamp 1
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_122
timestamp 1636968456
transform 1 0 11776 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_134
timestamp 1
transform 1 0 12880 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_148
timestamp 1
transform 1 0 14168 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_156
timestamp 1
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_197
timestamp 1
transform 1 0 18676 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_214
timestamp 1
transform 1 0 20240 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_246
timestamp 1
transform 1 0 23184 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_309
timestamp 1
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_3
timestamp 1
transform 1 0 828 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_9
timestamp 1
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1636968456
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 1
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_65
timestamp 1
transform 1 0 6532 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_79
timestamp 1
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_99
timestamp 1
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_122
timestamp 1
transform 1 0 11776 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_128
timestamp 1
transform 1 0 12328 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_160
timestamp 1
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1
transform 1 0 16100 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_173
timestamp 1
transform 1 0 16468 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_190
timestamp 1
transform 1 0 18032 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_194
timestamp 1
transform 1 0 18400 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp 1
transform 1 0 20792 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_225
timestamp 1
transform 1 0 21252 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_233
timestamp 1
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_239
timestamp 1
transform 1 0 22540 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_253
timestamp 1
transform 1 0 23828 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_257
timestamp 1636968456
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_269
timestamp 1
transform 1 0 25300 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1
transform 1 0 26036 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1636968456
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_293
timestamp 1
transform 1 0 27508 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_302
timestamp 1
transform 1 0 28336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_321
timestamp 1
transform 1 0 30084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_331
timestamp 1
transform 1 0 31004 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636968456
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_15
timestamp 1
transform 1 0 1932 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_19
timestamp 1
transform 1 0 2300 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 1
transform 1 0 2852 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636968456
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1636968456
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_53
timestamp 1
transform 1 0 5428 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_63
timestamp 1
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1
transform 1 0 7912 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1
transform 1 0 8372 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_93
timestamp 1
transform 1 0 9108 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_124
timestamp 1
transform 1 0 11960 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_133
timestamp 1
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_157
timestamp 1
transform 1 0 14996 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_165
timestamp 1
transform 1 0 15732 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_182
timestamp 1636968456
transform 1 0 17296 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_197
timestamp 1
transform 1 0 18676 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_216
timestamp 1
transform 1 0 20424 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_230
timestamp 1636968456
transform 1 0 21712 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_242
timestamp 1
transform 1 0 22816 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1
transform 1 0 23552 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1636968456
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1636968456
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1636968456
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1636968456
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_316
timestamp 1636968456
transform 1 0 29624 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_328
timestamp 1
transform 1 0 30728 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_334
timestamp 1
transform 1 0 31280 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636968456
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_15
timestamp 1
transform 1 0 1932 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_26
timestamp 1
transform 1 0 2944 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_38
timestamp 1636968456
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_50
timestamp 1
transform 1 0 5152 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_76
timestamp 1
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_84
timestamp 1
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_99
timestamp 1
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_104
timestamp 1
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_117
timestamp 1636968456
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_129
timestamp 1
transform 1 0 12420 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_141
timestamp 1
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_145
timestamp 1
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1
transform 1 0 16100 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1636968456
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_193
timestamp 1
transform 1 0 18308 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_199
timestamp 1
transform 1 0 18860 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_203
timestamp 1
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_217
timestamp 1
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_238
timestamp 1636968456
transform 1 0 22448 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_250
timestamp 1
transform 1 0 23552 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_266
timestamp 1
transform 1 0 25024 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_286
timestamp 1
transform 1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_305
timestamp 1
transform 1 0 28612 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_3
timestamp 1
transform 1 0 828 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1
transform 1 0 7820 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636968456
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_97
timestamp 1
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_118
timestamp 1
transform 1 0 11408 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_124
timestamp 1
transform 1 0 11960 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_192
timestamp 1
transform 1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1636968456
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_209
timestamp 1
transform 1 0 19780 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_224
timestamp 1
transform 1 0 21160 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_247
timestamp 1
transform 1 0 23276 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_285
timestamp 1
transform 1 0 26772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_298
timestamp 1
transform 1 0 27968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_314
timestamp 1
transform 1 0 29440 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_334
timestamp 1
transform 1 0 31280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1
transform 1 0 828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_11
timestamp 1
transform 1 0 1564 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_36
timestamp 1
transform 1 0 3864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_84
timestamp 1636968456
transform 1 0 8280 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_96
timestamp 1
transform 1 0 9384 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_104
timestamp 1
transform 1 0 10120 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_113
timestamp 1
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_122
timestamp 1
transform 1 0 11776 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_128
timestamp 1
transform 1 0 12328 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_140
timestamp 1
transform 1 0 13432 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_156
timestamp 1636968456
transform 1 0 14904 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_169
timestamp 1
transform 1 0 16100 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_178
timestamp 1
transform 1 0 16928 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_184
timestamp 1
transform 1 0 17480 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_196
timestamp 1
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_205
timestamp 1
transform 1 0 19412 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_213
timestamp 1
transform 1 0 20148 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_225
timestamp 1
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_245
timestamp 1
transform 1 0 23092 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_305
timestamp 1
transform 1 0 28612 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_333
timestamp 1
transform 1 0 31188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 1
transform 1 0 828 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_11
timestamp 1
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_16
timestamp 1
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_71
timestamp 1
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1636968456
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_112
timestamp 1
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_125
timestamp 1636968456
transform 1 0 12052 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1
transform 1 0 13524 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_162
timestamp 1
transform 1 0 15456 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_170
timestamp 1
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1636968456
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_209
timestamp 1
transform 1 0 19780 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_217
timestamp 1
transform 1 0 20516 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_225
timestamp 1
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 1
transform 1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_253
timestamp 1
transform 1 0 23828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_262
timestamp 1
transform 1 0 24656 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_272
timestamp 1
transform 1 0 25576 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_276
timestamp 1
transform 1 0 25944 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_285
timestamp 1
transform 1 0 26772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_294
timestamp 1
transform 1 0 27600 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_306
timestamp 1
transform 1 0 28704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_309
timestamp 1
transform 1 0 28980 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_324
timestamp 1
transform 1 0 30360 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_333
timestamp 1
transform 1 0 31188 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_44
timestamp 1
transform 1 0 4600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_69
timestamp 1
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_80
timestamp 1636968456
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_92
timestamp 1
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_117
timestamp 1
transform 1 0 11316 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_126
timestamp 1636968456
transform 1 0 12144 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_138
timestamp 1
transform 1 0 13248 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_146
timestamp 1
transform 1 0 13984 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_154
timestamp 1636968456
transform 1 0 14720 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_175
timestamp 1
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_210
timestamp 1
transform 1 0 19872 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_238
timestamp 1
transform 1 0 22448 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_243
timestamp 1636968456
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_260
timestamp 1
transform 1 0 24472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_292
timestamp 1
transform 1 0 27416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_299
timestamp 1
transform 1 0 28060 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_315
timestamp 1636968456
transform 1 0 29532 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_327
timestamp 1
transform 1 0 30636 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1
transform 1 0 828 0 1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_45
timestamp 1636968456
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_57
timestamp 1
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_65
timestamp 1
transform 1 0 6532 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_85
timestamp 1
transform 1 0 8372 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_91
timestamp 1
transform 1 0 8924 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_119
timestamp 1
transform 1 0 11500 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_127
timestamp 1
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_136
timestamp 1
transform 1 0 13064 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_158
timestamp 1
transform 1 0 15088 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_162
timestamp 1
transform 1 0 15456 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_176
timestamp 1
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_190
timestamp 1
transform 1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_216
timestamp 1
transform 1 0 20424 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_261
timestamp 1
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_279
timestamp 1
transform 1 0 26220 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_299
timestamp 1
transform 1 0 28060 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_322
timestamp 1636968456
transform 1 0 30176 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_334
timestamp 1
transform 1 0 31280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1
transform 1 0 828 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_48
timestamp 1
transform 1 0 4968 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 1
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_61
timestamp 1
transform 1 0 6164 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_89
timestamp 1
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636968456
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_125
timestamp 1
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_145
timestamp 1636968456
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_157
timestamp 1
transform 1 0 14996 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_184
timestamp 1
transform 1 0 17480 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_192
timestamp 1
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_243
timestamp 1
transform 1 0 22908 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_252
timestamp 1
transform 1 0 23736 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_256
timestamp 1
transform 1 0 24104 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_289
timestamp 1
transform 1 0 27140 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_332
timestamp 1
transform 1 0 31096 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1636968456
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_15
timestamp 1
transform 1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_19
timestamp 1
transform 1 0 2300 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_35
timestamp 1
transform 1 0 3772 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_42
timestamp 1636968456
transform 1 0 4416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_54
timestamp 1
transform 1 0 5520 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_62
timestamp 1
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1636968456
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_97
timestamp 1
transform 1 0 9476 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_111
timestamp 1636968456
transform 1 0 10764 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_123
timestamp 1
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_127
timestamp 1
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_152
timestamp 1
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_190
timestamp 1
transform 1 0 18032 0 1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1636968456
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_209
timestamp 1
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_220
timestamp 1
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_262
timestamp 1
transform 1 0 24656 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_285
timestamp 1
transform 1 0 26772 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_293
timestamp 1
transform 1 0 27508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_328
timestamp 1
transform 1 0 30728 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_334
timestamp 1
transform 1 0 31280 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636968456
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_31
timestamp 1
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_42
timestamp 1636968456
transform 1 0 4416 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_61
timestamp 1
transform 1 0 6164 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_71
timestamp 1
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_90
timestamp 1
transform 1 0 8832 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_96
timestamp 1
transform 1 0 9384 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_131
timestamp 1
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_140
timestamp 1
transform 1 0 13432 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_146
timestamp 1
transform 1 0 13984 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_152
timestamp 1
transform 1 0 14536 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_161
timestamp 1
transform 1 0 15364 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_183
timestamp 1636968456
transform 1 0 17388 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_195
timestamp 1636968456
transform 1 0 18492 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_207
timestamp 1
transform 1 0 19596 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_213
timestamp 1
transform 1 0 20148 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1
transform 1 0 20976 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_251
timestamp 1
transform 1 0 23644 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_257
timestamp 1
transform 1 0 24196 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_269
timestamp 1
transform 1 0 25300 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_277
timestamp 1
transform 1 0 26036 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1636968456
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_328
timestamp 1
transform 1 0 30728 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_334
timestamp 1
transform 1 0 31280 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1
transform 1 0 828 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_45
timestamp 1636968456
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_57
timestamp 1
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_71
timestamp 1
transform 1 0 7084 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_85
timestamp 1
transform 1 0 8372 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_93
timestamp 1
transform 1 0 9108 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_132
timestamp 1
transform 1 0 12696 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 1
transform 1 0 13524 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_197
timestamp 1
transform 1 0 18676 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_213
timestamp 1
transform 1 0 20148 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_219
timestamp 1
transform 1 0 20700 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_227
timestamp 1636968456
transform 1 0 21436 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_239
timestamp 1
transform 1 0 22540 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_253
timestamp 1
transform 1 0 23828 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_272
timestamp 1
transform 1 0 25576 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_288
timestamp 1
transform 1 0 27048 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_294
timestamp 1
transform 1 0 27600 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_323
timestamp 1636968456
transform 1 0 30268 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636968456
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_45
timestamp 1
transform 1 0 4692 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1
transform 1 0 5244 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_57
timestamp 1
transform 1 0 5796 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_65
timestamp 1
transform 1 0 6532 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_71
timestamp 1
transform 1 0 7084 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_77
timestamp 1636968456
transform 1 0 7636 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_89
timestamp 1636968456
transform 1 0 8740 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_101
timestamp 1
transform 1 0 9844 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_113
timestamp 1
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1636968456
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1636968456
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_149
timestamp 1
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_185
timestamp 1636968456
transform 1 0 17572 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_197
timestamp 1636968456
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_209
timestamp 1
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_215
timestamp 1
transform 1 0 20332 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_244
timestamp 1
transform 1 0 23000 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_252
timestamp 1
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_297
timestamp 1
transform 1 0 27876 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_301
timestamp 1
transform 1 0 28244 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_326
timestamp 1
transform 1 0 30544 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_334
timestamp 1
transform 1 0 31280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_3
timestamp 1
transform 1 0 828 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_11
timestamp 1
transform 1 0 1564 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_34
timestamp 1
transform 1 0 3680 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_44
timestamp 1636968456
transform 1 0 4600 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_56
timestamp 1
transform 1 0 5704 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_68
timestamp 1636968456
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_80
timestamp 1
transform 1 0 7912 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1
transform 1 0 8372 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_91
timestamp 1
transform 1 0 8924 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_95
timestamp 1636968456
transform 1 0 9292 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_107
timestamp 1
transform 1 0 10396 0 1 19040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_118
timestamp 1636968456
transform 1 0 11408 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_130
timestamp 1
transform 1 0 12512 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_141
timestamp 1
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_149
timestamp 1
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1
transform 1 0 17940 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1
transform 1 0 18492 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_197
timestamp 1
transform 1 0 18676 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_203
timestamp 1636968456
transform 1 0 19228 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_215
timestamp 1
transform 1 0 20332 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_235
timestamp 1
transform 1 0 22172 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_247
timestamp 1
transform 1 0 23276 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1
transform 1 0 23644 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_253
timestamp 1
transform 1 0 23828 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_283
timestamp 1
transform 1 0 26588 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_309
timestamp 1
transform 1 0 28980 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_329
timestamp 1
transform 1 0 30820 0 1 19040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1636968456
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_47
timestamp 1
transform 1 0 4876 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 1
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_65
timestamp 1
transform 1 0 6532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_69
timestamp 1
transform 1 0 6900 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_77
timestamp 1
transform 1 0 7636 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_88
timestamp 1
transform 1 0 8648 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1
transform 1 0 10212 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1
transform 1 0 10764 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_113
timestamp 1
transform 1 0 10948 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_122
timestamp 1636968456
transform 1 0 11776 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_134
timestamp 1
transform 1 0 12880 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_138
timestamp 1
transform 1 0 13248 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_187
timestamp 1
transform 1 0 17756 0 -1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_211
timestamp 1636968456
transform 1 0 19964 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_225
timestamp 1
transform 1 0 21252 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_229
timestamp 1
transform 1 0 21620 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_235
timestamp 1
transform 1 0 22172 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_257
timestamp 1
transform 1 0 24196 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_265
timestamp 1
transform 1 0 24932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_275
timestamp 1
transform 1 0 25852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1
transform 1 0 26220 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1636968456
transform 1 0 26404 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_300
timestamp 1
transform 1 0 28152 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_306
timestamp 1
transform 1 0 28704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_331
timestamp 1
transform 1 0 31004 0 -1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1636968456
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_15
timestamp 1
transform 1 0 1932 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_19
timestamp 1
transform 1 0 2300 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_29
timestamp 1
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_39
timestamp 1
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_70
timestamp 1
transform 1 0 6992 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_78
timestamp 1
transform 1 0 7728 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_89
timestamp 1
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_107
timestamp 1
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_128
timestamp 1
transform 1 0 12328 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_136
timestamp 1
transform 1 0 13064 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_160
timestamp 1
transform 1 0 15272 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_222
timestamp 1
transform 1 0 20976 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_230
timestamp 1
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_246
timestamp 1
transform 1 0 23184 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_253
timestamp 1
transform 1 0 23828 0 1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_291
timestamp 1636968456
transform 1 0 27324 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_303
timestamp 1
transform 1 0 28428 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1
transform 1 0 28796 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_331
timestamp 1
transform 1 0 31004 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_3
timestamp 1
transform 1 0 828 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_45
timestamp 1
transform 1 0 4692 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_51
timestamp 1
transform 1 0 5244 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_81
timestamp 1
transform 1 0 8004 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 1
transform 1 0 10948 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_137
timestamp 1
transform 1 0 13156 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_141
timestamp 1
transform 1 0 13524 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_145
timestamp 1636968456
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_157
timestamp 1
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_196
timestamp 1
transform 1 0 18584 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_216
timestamp 1
transform 1 0 20424 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1
transform 1 0 30820 0 -1 21216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636968456
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_15
timestamp 1
transform 1 0 1932 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_21
timestamp 1
transform 1 0 2484 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_33
timestamp 1
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1636968456
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_53
timestamp 1
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_57
timestamp 1
transform 1 0 5796 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_72
timestamp 1
transform 1 0 7176 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_91
timestamp 1
transform 1 0 8924 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_109
timestamp 1
transform 1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_113
timestamp 1
transform 1 0 10948 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_125
timestamp 1
transform 1 0 12052 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_130
timestamp 1
transform 1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_136
timestamp 1
transform 1 0 13064 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1636968456
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_153
timestamp 1
transform 1 0 14628 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_161
timestamp 1
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_165
timestamp 1
transform 1 0 15732 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_169
timestamp 1
transform 1 0 16100 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_181
timestamp 1636968456
transform 1 0 17204 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1
transform 1 0 18308 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_197
timestamp 1
transform 1 0 18676 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_210
timestamp 1636968456
transform 1 0 19872 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_222
timestamp 1
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_225
timestamp 1
transform 1 0 21252 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_232
timestamp 1636968456
transform 1 0 21896 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1
transform 1 0 23000 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_256
timestamp 1
transform 1 0 24104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_262
timestamp 1
transform 1 0 24656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_268
timestamp 1
transform 1 0 25208 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_281
timestamp 1
transform 1 0 26404 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_304
timestamp 1
transform 1 0 28520 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_319
timestamp 1636968456
transform 1 0 29900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_331
timestamp 1
transform 1 0 31004 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 21988 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 10120 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 5704 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 21344 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 25208 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform 1 0 6164 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 27324 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 28152 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 18400 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform 1 0 29900 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 10856 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 29256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 8280 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 14260 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 14260 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 28428 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform 1 0 7176 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform 1 0 28980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 14536 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 29808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform 1 0 26404 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform 1 0 30636 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 31004 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 23368 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 25576 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 22448 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 30820 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform 1 0 29256 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 31372 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 28612 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform 1 0 14076 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 30452 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 19688 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 28888 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform 1 0 11408 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 26772 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 7268 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform 1 0 30636 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 30452 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform -1 0 24472 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 3864 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform -1 0 4140 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform 1 0 3220 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform 1 0 3220 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 8004 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 28704 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 3036 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform -1 0 23460 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 3956 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 3128 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform -1 0 25852 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1
transform 1 0 28980 0 1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 28520 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 28244 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 26036 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 26312 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 25760 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 25208 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 24656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform -1 0 24104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform -1 0 21896 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap17
timestamp 1
transform -1 0 10212 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_61
timestamp 1
transform -1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_62
timestamp 1
transform -1 0 8924 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_63
timestamp 1
transform -1 0 7544 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_64
timestamp 1
transform -1 0 13064 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_65
timestamp 1
transform -1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_66
timestamp 1
transform -1 0 12052 0 1 21216
box -38 -48 314 592
<< labels >>
flabel metal4 s 4316 496 4636 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12090 496 12410 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19864 496 20184 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27638 496 27958 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11430 496 11750 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19204 496 19524 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26978 496 27298 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 29318 22104 29378 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 28214 22104 28274 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 27662 22104 27722 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 27110 22104 27170 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 26006 22104 26066 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 25454 22104 25514 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 24902 22104 24962 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 23798 22104 23858 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 23246 22104 23306 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 22694 22104 22754 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 21590 22104 21650 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 21038 22104 21098 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 20486 22104 20546 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 19382 22104 19442 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 9998 22104 10058 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal4 s 9446 22104 9506 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal4 s 8342 22104 8402 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal4 s 7790 22104 7850 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal4 s 7238 22104 7298 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal4 s 6134 22104 6194 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal4 s 14414 22104 14474 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal output
flabel metal4 s 13862 22104 13922 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal output
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal output
flabel metal4 s 12758 22104 12818 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal output
flabel metal4 s 12206 22104 12266 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal output
flabel metal4 s 11654 22104 11714 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal output
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal output
flabel metal4 s 10550 22104 10610 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal output
flabel metal4 s 18830 22104 18890 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal output
flabel metal4 s 18278 22104 18338 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal output
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal output
flabel metal4 s 17174 22104 17234 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal output
flabel metal4 s 16622 22104 16682 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal output
flabel metal4 s 16070 22104 16130 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal output
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal output
flabel metal4 s 14966 22104 15026 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
