VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 73.150 BY 33.600 ;
  OBS
      LAYER met1 ;
        RECT 0.000 33.250 8.050 33.600 ;
      LAYER met1 ;
        RECT 8.050 33.250 11.550 33.600 ;
      LAYER met1 ;
        RECT 11.550 33.250 73.150 33.600 ;
        RECT 0.000 32.900 6.650 33.250 ;
      LAYER met1 ;
        RECT 6.650 32.900 12.950 33.250 ;
      LAYER met1 ;
        RECT 12.950 32.900 73.150 33.250 ;
        RECT 0.000 32.550 5.600 32.900 ;
      LAYER met1 ;
        RECT 5.600 32.550 13.650 32.900 ;
      LAYER met1 ;
        RECT 13.650 32.550 73.150 32.900 ;
        RECT 0.000 32.200 4.900 32.550 ;
      LAYER met1 ;
        RECT 4.900 32.200 14.350 32.550 ;
      LAYER met1 ;
        RECT 14.350 32.200 48.650 32.550 ;
      LAYER met1 ;
        RECT 48.650 32.200 49.350 32.550 ;
      LAYER met1 ;
        RECT 49.350 32.200 53.200 32.550 ;
      LAYER met1 ;
        RECT 53.200 32.200 53.550 32.550 ;
      LAYER met1 ;
        RECT 53.550 32.200 57.400 32.550 ;
      LAYER met1 ;
        RECT 57.400 32.200 57.750 32.550 ;
      LAYER met1 ;
        RECT 57.750 32.200 73.150 32.550 ;
        RECT 0.000 31.850 4.550 32.200 ;
      LAYER met1 ;
        RECT 4.550 31.850 8.750 32.200 ;
      LAYER met1 ;
        RECT 8.750 31.850 10.850 32.200 ;
      LAYER met1 ;
        RECT 10.850 31.850 15.050 32.200 ;
      LAYER met1 ;
        RECT 15.050 31.850 47.600 32.200 ;
      LAYER met1 ;
        RECT 47.600 31.850 50.050 32.200 ;
      LAYER met1 ;
        RECT 50.050 31.850 52.500 32.200 ;
      LAYER met1 ;
        RECT 52.500 31.850 54.250 32.200 ;
      LAYER met1 ;
        RECT 54.250 31.850 56.000 32.200 ;
      LAYER met1 ;
        RECT 56.000 31.850 58.450 32.200 ;
      LAYER met1 ;
        RECT 58.450 31.850 60.550 32.200 ;
      LAYER met1 ;
        RECT 60.550 31.850 63.000 32.200 ;
      LAYER met1 ;
        RECT 63.000 31.850 73.150 32.200 ;
        RECT 0.000 31.500 3.850 31.850 ;
      LAYER met1 ;
        RECT 3.850 31.500 7.000 31.850 ;
      LAYER met1 ;
        RECT 7.000 31.500 12.250 31.850 ;
      LAYER met1 ;
        RECT 12.250 31.500 15.400 31.850 ;
      LAYER met1 ;
        RECT 15.400 31.500 47.600 31.850 ;
      LAYER met1 ;
        RECT 47.600 31.500 48.300 31.850 ;
      LAYER met1 ;
        RECT 48.300 31.500 49.350 31.850 ;
      LAYER met1 ;
        RECT 49.350 31.500 50.400 31.850 ;
      LAYER met1 ;
        RECT 50.400 31.500 52.150 31.850 ;
      LAYER met1 ;
        RECT 52.150 31.500 52.850 31.850 ;
      LAYER met1 ;
        RECT 52.850 31.500 53.900 31.850 ;
        RECT 0.000 31.150 3.500 31.500 ;
      LAYER met1 ;
        RECT 3.500 31.150 6.300 31.500 ;
      LAYER met1 ;
        RECT 6.300 31.150 13.300 31.500 ;
      LAYER met1 ;
        RECT 13.300 31.150 16.100 31.500 ;
      LAYER met1 ;
        RECT 16.100 31.150 49.700 31.500 ;
      LAYER met1 ;
        RECT 49.700 31.150 50.400 31.500 ;
      LAYER met1 ;
        RECT 50.400 31.150 51.800 31.500 ;
        RECT 0.000 30.800 3.150 31.150 ;
      LAYER met1 ;
        RECT 3.150 30.800 5.600 31.150 ;
      LAYER met1 ;
        RECT 5.600 30.800 14.000 31.150 ;
      LAYER met1 ;
        RECT 14.000 30.800 16.450 31.150 ;
      LAYER met1 ;
        RECT 16.450 30.800 50.050 31.150 ;
      LAYER met1 ;
        RECT 50.050 30.800 50.750 31.150 ;
      LAYER met1 ;
        RECT 50.750 30.800 51.800 31.150 ;
        RECT 0.000 30.450 2.800 30.800 ;
      LAYER met1 ;
        RECT 2.800 30.450 4.900 30.800 ;
      LAYER met1 ;
        RECT 4.900 30.450 14.350 30.800 ;
      LAYER met1 ;
        RECT 14.350 30.450 16.800 30.800 ;
      LAYER met1 ;
        RECT 16.800 30.450 49.700 30.800 ;
        RECT 0.000 30.100 2.450 30.450 ;
      LAYER met1 ;
        RECT 2.450 30.100 4.550 30.450 ;
      LAYER met1 ;
        RECT 4.550 30.100 15.050 30.450 ;
      LAYER met1 ;
        RECT 15.050 30.100 17.150 30.450 ;
      LAYER met1 ;
        RECT 17.150 30.100 49.700 30.450 ;
      LAYER met1 ;
        RECT 49.700 30.100 50.400 30.800 ;
      LAYER met1 ;
        RECT 0.000 29.750 2.100 30.100 ;
      LAYER met1 ;
        RECT 2.100 29.750 4.200 30.100 ;
      LAYER met1 ;
        RECT 4.200 29.750 15.400 30.100 ;
      LAYER met1 ;
        RECT 15.400 29.750 17.500 30.100 ;
      LAYER met1 ;
        RECT 0.000 29.050 1.750 29.750 ;
      LAYER met1 ;
        RECT 1.750 29.400 3.850 29.750 ;
      LAYER met1 ;
        RECT 3.850 29.400 15.750 29.750 ;
      LAYER met1 ;
        RECT 15.750 29.400 17.500 29.750 ;
      LAYER met1 ;
        RECT 17.500 29.400 49.350 30.100 ;
      LAYER met1 ;
        RECT 49.350 29.750 50.400 30.100 ;
      LAYER met1 ;
        RECT 50.400 29.750 51.800 30.800 ;
      LAYER met1 ;
        RECT 49.350 29.400 50.050 29.750 ;
      LAYER met1 ;
        RECT 50.050 29.400 51.800 29.750 ;
      LAYER met1 ;
        RECT 1.750 29.050 11.550 29.400 ;
      LAYER met1 ;
        RECT 11.550 29.050 16.100 29.400 ;
      LAYER met1 ;
        RECT 16.100 29.050 17.850 29.400 ;
      LAYER met1 ;
        RECT 17.850 29.050 49.000 29.400 ;
      LAYER met1 ;
        RECT 49.000 29.050 49.700 29.400 ;
      LAYER met1 ;
        RECT 49.700 29.050 51.800 29.400 ;
        RECT 0.000 28.700 1.400 29.050 ;
      LAYER met1 ;
        RECT 1.400 28.700 11.550 29.050 ;
      LAYER met1 ;
        RECT 0.000 28.000 1.050 28.700 ;
      LAYER met1 ;
        RECT 1.050 28.000 11.550 28.700 ;
      LAYER met1 ;
        RECT 11.550 28.350 16.450 29.050 ;
      LAYER met1 ;
        RECT 16.450 28.350 18.200 29.050 ;
      LAYER met1 ;
        RECT 18.200 28.700 22.750 29.050 ;
      LAYER met1 ;
        RECT 22.750 28.700 25.200 29.050 ;
      LAYER met1 ;
        RECT 25.200 28.700 31.850 29.050 ;
      LAYER met1 ;
        RECT 31.850 28.700 34.650 29.050 ;
      LAYER met1 ;
        RECT 34.650 28.700 48.650 29.050 ;
      LAYER met1 ;
        RECT 48.650 28.700 49.350 29.050 ;
      LAYER met1 ;
        RECT 49.350 28.700 51.800 29.050 ;
        RECT 18.200 28.350 22.050 28.700 ;
      LAYER met1 ;
        RECT 22.050 28.350 25.200 28.700 ;
      LAYER met1 ;
        RECT 25.200 28.350 31.150 28.700 ;
      LAYER met1 ;
        RECT 31.150 28.350 35.700 28.700 ;
      LAYER met1 ;
        RECT 35.700 28.350 48.300 28.700 ;
      LAYER met1 ;
        RECT 48.300 28.350 49.000 28.700 ;
      LAYER met1 ;
        RECT 49.000 28.350 51.800 28.700 ;
        RECT 0.000 26.950 0.700 28.000 ;
      LAYER met1 ;
        RECT 0.700 26.950 11.550 28.000 ;
      LAYER met1 ;
        RECT 11.550 27.650 16.800 28.350 ;
      LAYER met1 ;
        RECT 16.800 27.650 18.550 28.350 ;
      LAYER met1 ;
        RECT 18.550 28.000 21.700 28.350 ;
      LAYER met1 ;
        RECT 21.700 28.000 25.200 28.350 ;
      LAYER met1 ;
        RECT 25.200 28.000 30.800 28.350 ;
      LAYER met1 ;
        RECT 30.800 28.000 32.900 28.350 ;
      LAYER met1 ;
        RECT 32.900 28.000 33.950 28.350 ;
      LAYER met1 ;
        RECT 33.950 28.000 36.050 28.350 ;
      LAYER met1 ;
        RECT 36.050 28.000 47.950 28.350 ;
      LAYER met1 ;
        RECT 47.950 28.000 48.650 28.350 ;
      LAYER met1 ;
        RECT 48.650 28.000 51.800 28.350 ;
      LAYER met1 ;
        RECT 51.800 28.000 52.500 31.500 ;
      LAYER met1 ;
        RECT 52.500 31.150 53.900 31.500 ;
      LAYER met1 ;
        RECT 53.900 31.150 54.600 31.850 ;
      LAYER met1 ;
        RECT 54.600 31.500 56.000 31.850 ;
      LAYER met1 ;
        RECT 56.000 31.500 56.700 31.850 ;
      LAYER met1 ;
        RECT 56.700 31.500 57.750 31.850 ;
      LAYER met1 ;
        RECT 57.750 31.500 58.800 31.850 ;
      LAYER met1 ;
        RECT 58.800 31.500 60.550 31.850 ;
      LAYER met1 ;
        RECT 60.550 31.500 61.250 31.850 ;
      LAYER met1 ;
        RECT 61.250 31.500 73.150 31.850 ;
        RECT 54.600 31.150 58.100 31.500 ;
      LAYER met1 ;
        RECT 58.100 31.150 59.150 31.500 ;
      LAYER met1 ;
        RECT 52.500 30.100 54.250 31.150 ;
        RECT 52.500 29.400 52.850 30.100 ;
      LAYER met1 ;
        RECT 52.850 29.400 53.900 30.100 ;
      LAYER met1 ;
        RECT 53.900 29.400 54.250 30.100 ;
        RECT 52.500 28.350 54.250 29.400 ;
      LAYER met1 ;
        RECT 54.250 28.350 54.950 31.150 ;
      LAYER met1 ;
        RECT 54.950 30.450 58.450 31.150 ;
      LAYER met1 ;
        RECT 58.450 30.450 59.150 31.150 ;
      LAYER met1 ;
        RECT 59.150 30.450 60.550 31.500 ;
      LAYER met1 ;
        RECT 60.550 30.450 60.900 31.500 ;
      LAYER met1 ;
        RECT 60.900 30.450 73.150 31.500 ;
        RECT 54.950 29.750 58.100 30.450 ;
      LAYER met1 ;
        RECT 58.100 29.750 58.800 30.450 ;
      LAYER met1 ;
        RECT 58.800 29.750 60.550 30.450 ;
      LAYER met1 ;
        RECT 60.550 30.100 62.650 30.450 ;
      LAYER met1 ;
        RECT 62.650 30.100 73.150 30.450 ;
      LAYER met1 ;
        RECT 60.550 29.750 60.900 30.100 ;
      LAYER met1 ;
        RECT 60.900 29.750 61.950 30.100 ;
      LAYER met1 ;
        RECT 61.950 29.750 63.000 30.100 ;
      LAYER met1 ;
        RECT 63.000 29.750 73.150 30.100 ;
        RECT 54.950 29.400 57.750 29.750 ;
      LAYER met1 ;
        RECT 57.750 29.400 58.450 29.750 ;
      LAYER met1 ;
        RECT 58.450 29.400 62.300 29.750 ;
      LAYER met1 ;
        RECT 62.300 29.400 63.350 29.750 ;
      LAYER met1 ;
        RECT 54.950 29.050 57.400 29.400 ;
      LAYER met1 ;
        RECT 57.400 29.050 58.100 29.400 ;
      LAYER met1 ;
        RECT 58.100 29.050 62.650 29.400 ;
        RECT 54.950 28.700 57.050 29.050 ;
      LAYER met1 ;
        RECT 57.050 28.700 57.750 29.050 ;
      LAYER met1 ;
        RECT 57.750 28.700 62.650 29.050 ;
        RECT 54.950 28.350 56.700 28.700 ;
      LAYER met1 ;
        RECT 56.700 28.350 57.400 28.700 ;
      LAYER met1 ;
        RECT 57.400 28.350 62.650 28.700 ;
        RECT 52.500 28.000 53.900 28.350 ;
      LAYER met1 ;
        RECT 53.900 28.000 54.950 28.350 ;
      LAYER met1 ;
        RECT 54.950 28.000 56.350 28.350 ;
      LAYER met1 ;
        RECT 56.350 28.000 57.050 28.350 ;
      LAYER met1 ;
        RECT 57.050 28.000 62.650 28.350 ;
      LAYER met1 ;
        RECT 62.650 28.000 63.350 29.400 ;
      LAYER met1 ;
        RECT 63.350 28.000 73.150 29.750 ;
        RECT 18.550 27.650 21.000 28.000 ;
      LAYER met1 ;
        RECT 21.000 27.650 25.200 28.000 ;
      LAYER met1 ;
        RECT 25.200 27.650 30.450 28.000 ;
      LAYER met1 ;
        RECT 30.450 27.650 32.200 28.000 ;
      LAYER met1 ;
        RECT 11.550 26.950 17.150 27.650 ;
      LAYER met1 ;
        RECT 17.150 26.950 18.900 27.650 ;
      LAYER met1 ;
        RECT 0.000 25.900 5.950 26.950 ;
        RECT 0.000 25.550 0.350 25.900 ;
      LAYER met1 ;
        RECT 0.350 25.550 1.750 25.900 ;
        RECT 0.000 25.200 1.750 25.550 ;
      LAYER met1 ;
        RECT 1.750 25.200 5.950 25.900 ;
      LAYER met1 ;
        RECT 0.000 22.750 1.400 25.200 ;
      LAYER met1 ;
        RECT 1.400 22.750 5.950 25.200 ;
      LAYER met1 ;
        RECT 5.950 24.850 8.750 26.950 ;
      LAYER met1 ;
        RECT 8.750 26.250 17.500 26.950 ;
      LAYER met1 ;
        RECT 17.500 26.600 18.900 26.950 ;
      LAYER met1 ;
        RECT 18.900 26.600 20.650 27.650 ;
      LAYER met1 ;
        RECT 20.650 27.300 22.050 27.650 ;
      LAYER met1 ;
        RECT 22.050 27.300 22.750 27.650 ;
      LAYER met1 ;
        RECT 20.650 26.950 21.350 27.300 ;
      LAYER met1 ;
        RECT 21.350 26.950 22.750 27.300 ;
      LAYER met1 ;
        RECT 20.650 26.600 21.000 26.950 ;
      LAYER met1 ;
        RECT 21.000 26.600 22.750 26.950 ;
      LAYER met1 ;
        RECT 17.500 26.250 19.250 26.600 ;
      LAYER met1 ;
        RECT 8.750 24.850 17.850 26.250 ;
      LAYER met1 ;
        RECT 17.850 24.850 19.250 26.250 ;
      LAYER met1 ;
        RECT 19.250 24.850 22.750 26.600 ;
      LAYER met1 ;
        RECT 0.000 22.050 1.750 22.750 ;
      LAYER met1 ;
        RECT 0.000 20.650 0.350 22.050 ;
      LAYER met1 ;
        RECT 0.350 21.350 1.750 22.050 ;
      LAYER met1 ;
        RECT 1.750 21.350 5.950 22.750 ;
      LAYER met1 ;
        RECT 5.950 22.050 16.100 24.850 ;
      LAYER met1 ;
        RECT 16.100 22.050 17.850 24.850 ;
      LAYER met1 ;
        RECT 17.850 23.100 19.600 24.850 ;
      LAYER met1 ;
        RECT 19.600 23.100 22.750 24.850 ;
      LAYER met1 ;
        RECT 0.350 20.650 2.100 21.350 ;
      LAYER met1 ;
        RECT 0.000 19.950 0.700 20.650 ;
      LAYER met1 ;
        RECT 0.700 20.300 2.100 20.650 ;
      LAYER met1 ;
        RECT 2.100 20.300 5.950 21.350 ;
      LAYER met1 ;
        RECT 5.950 20.300 8.750 22.050 ;
      LAYER met1 ;
        RECT 8.750 20.300 10.500 22.050 ;
      LAYER met1 ;
        RECT 0.700 19.950 2.450 20.300 ;
      LAYER met1 ;
        RECT 0.000 19.250 1.050 19.950 ;
      LAYER met1 ;
        RECT 1.050 19.600 2.450 19.950 ;
      LAYER met1 ;
        RECT 2.450 19.600 10.500 20.300 ;
      LAYER met1 ;
        RECT 1.050 19.250 2.800 19.600 ;
      LAYER met1 ;
        RECT 2.800 19.250 10.500 19.600 ;
        RECT 0.000 18.550 1.400 19.250 ;
      LAYER met1 ;
        RECT 1.400 18.550 3.150 19.250 ;
      LAYER met1 ;
        RECT 3.150 18.550 10.500 19.250 ;
        RECT 0.000 18.200 1.750 18.550 ;
      LAYER met1 ;
        RECT 1.750 18.200 3.500 18.550 ;
      LAYER met1 ;
        RECT 3.500 18.200 10.500 18.550 ;
        RECT 0.000 17.500 2.100 18.200 ;
      LAYER met1 ;
        RECT 2.100 17.850 3.850 18.200 ;
      LAYER met1 ;
        RECT 3.850 17.850 10.500 18.200 ;
      LAYER met1 ;
        RECT 2.100 17.500 4.200 17.850 ;
      LAYER met1 ;
        RECT 4.200 17.500 10.500 17.850 ;
        RECT 0.000 17.150 2.450 17.500 ;
      LAYER met1 ;
        RECT 2.450 17.150 4.550 17.500 ;
      LAYER met1 ;
        RECT 4.550 17.150 10.500 17.500 ;
        RECT 0.000 16.800 2.800 17.150 ;
      LAYER met1 ;
        RECT 2.800 16.800 5.250 17.150 ;
      LAYER met1 ;
        RECT 5.250 16.800 10.500 17.150 ;
        RECT 0.000 16.450 3.150 16.800 ;
      LAYER met1 ;
        RECT 3.150 16.450 5.600 16.800 ;
      LAYER met1 ;
        RECT 5.600 16.450 10.500 16.800 ;
        RECT 0.000 16.100 3.500 16.450 ;
      LAYER met1 ;
        RECT 3.500 16.100 6.650 16.450 ;
      LAYER met1 ;
        RECT 6.650 16.100 10.500 16.450 ;
        RECT 0.000 15.750 4.200 16.100 ;
      LAYER met1 ;
        RECT 4.200 15.750 7.350 16.100 ;
      LAYER met1 ;
        RECT 7.350 15.750 10.500 16.100 ;
      LAYER met1 ;
        RECT 10.500 15.750 13.300 22.050 ;
      LAYER met1 ;
        RECT 13.300 21.700 17.850 22.050 ;
      LAYER met1 ;
        RECT 17.850 21.700 19.250 23.100 ;
      LAYER met1 ;
        RECT 13.300 20.650 17.500 21.700 ;
      LAYER met1 ;
        RECT 17.500 21.000 19.250 21.700 ;
      LAYER met1 ;
        RECT 19.250 21.000 22.750 23.100 ;
      LAYER met1 ;
        RECT 17.500 20.650 18.900 21.000 ;
      LAYER met1 ;
        RECT 13.300 19.950 17.150 20.650 ;
      LAYER met1 ;
        RECT 17.150 19.950 18.900 20.650 ;
      LAYER met1 ;
        RECT 18.900 19.950 22.750 21.000 ;
        RECT 13.300 19.250 16.800 19.950 ;
      LAYER met1 ;
        RECT 16.800 19.250 18.550 19.950 ;
      LAYER met1 ;
        RECT 18.550 19.600 22.750 19.950 ;
      LAYER met1 ;
        RECT 22.750 19.600 25.200 27.650 ;
      LAYER met1 ;
        RECT 25.200 27.300 30.100 27.650 ;
      LAYER met1 ;
        RECT 30.100 27.300 32.200 27.650 ;
      LAYER met1 ;
        RECT 32.200 27.300 34.300 28.000 ;
      LAYER met1 ;
        RECT 34.300 27.650 36.400 28.000 ;
      LAYER met1 ;
        RECT 36.400 27.650 47.600 28.000 ;
      LAYER met1 ;
        RECT 47.600 27.650 48.650 28.000 ;
      LAYER met1 ;
        RECT 48.650 27.650 52.150 28.000 ;
      LAYER met1 ;
        RECT 52.150 27.650 52.850 28.000 ;
      LAYER met1 ;
        RECT 52.850 27.650 53.900 28.000 ;
      LAYER met1 ;
        RECT 53.900 27.650 54.600 28.000 ;
      LAYER met1 ;
        RECT 54.600 27.650 56.000 28.000 ;
      LAYER met1 ;
        RECT 56.000 27.650 57.050 28.000 ;
      LAYER met1 ;
        RECT 57.050 27.650 60.200 28.000 ;
      LAYER met1 ;
        RECT 60.200 27.650 60.550 28.000 ;
      LAYER met1 ;
        RECT 60.550 27.650 61.950 28.000 ;
      LAYER met1 ;
        RECT 61.950 27.650 63.000 28.000 ;
      LAYER met1 ;
        RECT 63.000 27.650 73.150 28.000 ;
      LAYER met1 ;
        RECT 34.300 27.300 36.750 27.650 ;
      LAYER met1 ;
        RECT 36.750 27.300 47.600 27.650 ;
      LAYER met1 ;
        RECT 47.600 27.300 50.750 27.650 ;
      LAYER met1 ;
        RECT 50.750 27.300 52.500 27.650 ;
      LAYER met1 ;
        RECT 52.500 27.300 54.250 27.650 ;
      LAYER met1 ;
        RECT 54.250 27.300 56.000 27.650 ;
      LAYER met1 ;
        RECT 56.000 27.300 59.150 27.650 ;
      LAYER met1 ;
        RECT 59.150 27.300 60.200 27.650 ;
      LAYER met1 ;
        RECT 60.200 27.300 62.650 27.650 ;
      LAYER met1 ;
        RECT 62.650 27.300 73.150 27.650 ;
        RECT 25.200 26.600 29.750 27.300 ;
      LAYER met1 ;
        RECT 29.750 26.600 32.200 27.300 ;
      LAYER met1 ;
        RECT 32.200 26.600 34.650 27.300 ;
      LAYER met1 ;
        RECT 34.650 26.950 36.750 27.300 ;
      LAYER met1 ;
        RECT 36.750 26.950 52.850 27.300 ;
      LAYER met1 ;
        RECT 52.850 26.950 53.550 27.300 ;
      LAYER met1 ;
        RECT 53.550 26.950 60.900 27.300 ;
      LAYER met1 ;
        RECT 60.900 26.950 61.950 27.300 ;
      LAYER met1 ;
        RECT 61.950 26.950 73.150 27.300 ;
        RECT 25.200 25.200 29.400 26.600 ;
      LAYER met1 ;
        RECT 29.400 25.200 31.850 26.600 ;
      LAYER met1 ;
        RECT 25.200 22.750 29.050 25.200 ;
      LAYER met1 ;
        RECT 29.050 22.750 31.850 25.200 ;
      LAYER met1 ;
        RECT 25.200 21.350 29.400 22.750 ;
      LAYER met1 ;
        RECT 29.400 21.350 31.850 22.750 ;
      LAYER met1 ;
        RECT 25.200 20.300 29.750 21.350 ;
      LAYER met1 ;
        RECT 29.750 21.000 31.850 21.350 ;
      LAYER met1 ;
        RECT 31.850 21.000 34.650 26.600 ;
      LAYER met1 ;
        RECT 34.650 25.900 37.100 26.950 ;
      LAYER met1 ;
        RECT 37.100 25.900 73.150 26.950 ;
      LAYER met1 ;
        RECT 34.650 22.050 37.450 25.900 ;
      LAYER met1 ;
        RECT 37.450 24.500 73.150 25.900 ;
        RECT 37.450 24.150 52.500 24.500 ;
      LAYER met1 ;
        RECT 52.500 24.150 53.900 24.500 ;
      LAYER met1 ;
        RECT 53.900 24.150 67.550 24.500 ;
      LAYER met1 ;
        RECT 67.550 24.150 68.600 24.500 ;
      LAYER met1 ;
        RECT 68.600 24.150 73.150 24.500 ;
        RECT 37.450 23.800 40.600 24.150 ;
      LAYER met1 ;
        RECT 40.600 23.800 43.750 24.150 ;
      LAYER met1 ;
        RECT 43.750 23.800 46.550 24.150 ;
      LAYER met1 ;
        RECT 46.550 23.800 49.350 24.150 ;
      LAYER met1 ;
        RECT 49.350 23.800 51.450 24.150 ;
      LAYER met1 ;
        RECT 51.450 23.800 54.950 24.150 ;
      LAYER met1 ;
        RECT 54.950 23.800 56.700 24.150 ;
      LAYER met1 ;
        RECT 56.700 23.800 60.200 24.150 ;
      LAYER met1 ;
        RECT 60.200 23.800 66.150 24.150 ;
      LAYER met1 ;
        RECT 66.150 23.800 69.650 24.150 ;
      LAYER met1 ;
        RECT 69.650 23.800 73.150 24.150 ;
        RECT 37.450 23.450 41.300 23.800 ;
      LAYER met1 ;
        RECT 41.300 23.450 43.050 23.800 ;
      LAYER met1 ;
        RECT 43.050 23.450 47.250 23.800 ;
      LAYER met1 ;
        RECT 47.250 23.450 48.650 23.800 ;
      LAYER met1 ;
        RECT 48.650 23.450 51.100 23.800 ;
      LAYER met1 ;
        RECT 51.100 23.450 52.500 23.800 ;
      LAYER met1 ;
        RECT 52.500 23.450 53.200 23.800 ;
      LAYER met1 ;
        RECT 53.200 23.450 55.300 23.800 ;
      LAYER met1 ;
        RECT 55.300 23.450 57.400 23.800 ;
      LAYER met1 ;
        RECT 57.400 23.450 59.500 23.800 ;
      LAYER met1 ;
        RECT 59.500 23.450 65.450 23.800 ;
      LAYER met1 ;
        RECT 65.450 23.450 70.350 23.800 ;
      LAYER met1 ;
        RECT 70.350 23.450 73.150 23.800 ;
        RECT 37.450 22.400 41.650 23.450 ;
      LAYER met1 ;
        RECT 41.650 23.100 42.700 23.450 ;
      LAYER met1 ;
        RECT 42.700 23.100 47.250 23.450 ;
      LAYER met1 ;
        RECT 47.250 23.100 48.300 23.450 ;
      LAYER met1 ;
        RECT 48.300 23.100 50.750 23.450 ;
      LAYER met1 ;
        RECT 50.750 23.100 51.800 23.450 ;
      LAYER met1 ;
        RECT 51.800 23.100 53.900 23.450 ;
      LAYER met1 ;
        RECT 53.900 23.100 55.300 23.450 ;
      LAYER met1 ;
        RECT 55.300 23.100 57.750 23.450 ;
      LAYER met1 ;
        RECT 41.650 22.400 43.050 23.100 ;
      LAYER met1 ;
        RECT 43.050 22.400 47.250 23.100 ;
      LAYER met1 ;
        RECT 47.250 22.400 47.950 23.100 ;
      LAYER met1 ;
        RECT 47.950 22.750 50.750 23.100 ;
      LAYER met1 ;
        RECT 50.750 22.750 51.450 23.100 ;
      LAYER met1 ;
        RECT 51.450 22.750 54.250 23.100 ;
      LAYER met1 ;
        RECT 54.250 22.750 54.950 23.100 ;
      LAYER met1 ;
        RECT 54.950 22.750 57.750 23.100 ;
        RECT 37.450 22.050 42.000 22.400 ;
      LAYER met1 ;
        RECT 34.650 21.000 37.100 22.050 ;
      LAYER met1 ;
        RECT 37.100 21.350 42.000 22.050 ;
      LAYER met1 ;
        RECT 42.000 21.350 43.400 22.400 ;
      LAYER met1 ;
        RECT 43.400 21.700 46.900 22.400 ;
      LAYER met1 ;
        RECT 46.900 22.050 47.950 22.400 ;
      LAYER met1 ;
        RECT 47.950 22.050 50.400 22.750 ;
      LAYER met1 ;
        RECT 50.400 22.050 51.450 22.750 ;
      LAYER met1 ;
        RECT 51.450 22.050 57.750 22.750 ;
      LAYER met1 ;
        RECT 46.900 21.700 47.600 22.050 ;
      LAYER met1 ;
        RECT 43.400 21.350 46.550 21.700 ;
        RECT 37.100 21.000 42.350 21.350 ;
      LAYER met1 ;
        RECT 29.750 20.300 32.200 21.000 ;
      LAYER met1 ;
        RECT 32.200 20.300 34.650 21.000 ;
      LAYER met1 ;
        RECT 34.650 20.300 36.750 21.000 ;
      LAYER met1 ;
        RECT 36.750 20.650 42.350 21.000 ;
      LAYER met1 ;
        RECT 42.350 20.650 43.750 21.350 ;
      LAYER met1 ;
        RECT 43.750 20.650 46.550 21.350 ;
      LAYER met1 ;
        RECT 46.550 21.000 47.600 21.700 ;
      LAYER met1 ;
        RECT 47.600 21.350 50.400 22.050 ;
      LAYER met1 ;
        RECT 50.400 21.700 51.800 22.050 ;
      LAYER met1 ;
        RECT 51.800 21.700 57.750 22.050 ;
      LAYER met1 ;
        RECT 50.400 21.350 52.150 21.700 ;
      LAYER met1 ;
        RECT 52.150 21.350 57.750 21.700 ;
        RECT 47.600 21.000 50.750 21.350 ;
      LAYER met1 ;
        RECT 50.750 21.000 52.850 21.350 ;
      LAYER met1 ;
        RECT 52.850 21.000 57.750 21.350 ;
      LAYER met1 ;
        RECT 46.550 20.650 47.250 21.000 ;
      LAYER met1 ;
        RECT 47.250 20.650 50.750 21.000 ;
      LAYER met1 ;
        RECT 50.750 20.650 53.200 21.000 ;
      LAYER met1 ;
        RECT 53.200 20.650 57.750 21.000 ;
        RECT 36.750 20.300 42.700 20.650 ;
      LAYER met1 ;
        RECT 42.700 20.300 43.750 20.650 ;
      LAYER met1 ;
        RECT 43.750 20.300 46.200 20.650 ;
        RECT 25.200 19.950 30.100 20.300 ;
      LAYER met1 ;
        RECT 30.100 19.950 32.200 20.300 ;
      LAYER met1 ;
        RECT 32.200 19.950 34.300 20.300 ;
      LAYER met1 ;
        RECT 34.300 19.950 36.400 20.300 ;
      LAYER met1 ;
        RECT 36.400 19.950 42.700 20.300 ;
        RECT 25.200 19.600 30.450 19.950 ;
      LAYER met1 ;
        RECT 30.450 19.600 32.550 19.950 ;
      LAYER met1 ;
        RECT 32.550 19.600 34.300 19.950 ;
      LAYER met1 ;
        RECT 34.300 19.600 36.050 19.950 ;
      LAYER met1 ;
        RECT 36.050 19.600 42.700 19.950 ;
      LAYER met1 ;
        RECT 42.700 19.600 44.100 20.300 ;
      LAYER met1 ;
        RECT 44.100 19.600 46.200 20.300 ;
      LAYER met1 ;
        RECT 46.200 19.950 47.250 20.650 ;
      LAYER met1 ;
        RECT 47.250 20.300 51.450 20.650 ;
      LAYER met1 ;
        RECT 51.450 20.300 53.900 20.650 ;
      LAYER met1 ;
        RECT 53.900 20.300 57.750 20.650 ;
        RECT 47.250 19.950 51.800 20.300 ;
      LAYER met1 ;
        RECT 51.800 19.950 54.600 20.300 ;
      LAYER met1 ;
        RECT 54.600 19.950 57.750 20.300 ;
      LAYER met1 ;
        RECT 46.200 19.600 46.900 19.950 ;
      LAYER met1 ;
        RECT 46.900 19.600 52.500 19.950 ;
      LAYER met1 ;
        RECT 52.500 19.600 54.950 19.950 ;
      LAYER met1 ;
        RECT 54.950 19.600 57.750 19.950 ;
        RECT 18.550 19.250 20.650 19.600 ;
        RECT 13.300 18.900 16.450 19.250 ;
      LAYER met1 ;
        RECT 16.450 18.900 18.200 19.250 ;
      LAYER met1 ;
        RECT 18.200 18.900 20.650 19.250 ;
      LAYER met1 ;
        RECT 20.650 18.900 26.950 19.600 ;
      LAYER met1 ;
        RECT 26.950 19.250 30.800 19.600 ;
      LAYER met1 ;
        RECT 30.800 19.250 33.250 19.600 ;
      LAYER met1 ;
        RECT 33.250 19.250 33.600 19.600 ;
      LAYER met1 ;
        RECT 33.600 19.250 35.700 19.600 ;
      LAYER met1 ;
        RECT 35.700 19.250 43.050 19.600 ;
        RECT 26.950 18.900 31.150 19.250 ;
      LAYER met1 ;
        RECT 31.150 18.900 35.350 19.250 ;
      LAYER met1 ;
        RECT 35.350 18.900 43.050 19.250 ;
        RECT 13.300 18.550 16.100 18.900 ;
      LAYER met1 ;
        RECT 16.100 18.550 17.850 18.900 ;
      LAYER met1 ;
        RECT 17.850 18.550 32.200 18.900 ;
      LAYER met1 ;
        RECT 32.200 18.550 34.300 18.900 ;
      LAYER met1 ;
        RECT 34.300 18.550 43.050 18.900 ;
      LAYER met1 ;
        RECT 43.050 18.550 44.450 19.600 ;
      LAYER met1 ;
        RECT 44.450 18.550 45.850 19.600 ;
      LAYER met1 ;
        RECT 45.850 18.900 46.900 19.600 ;
      LAYER met1 ;
        RECT 46.900 19.250 53.200 19.600 ;
      LAYER met1 ;
        RECT 53.200 19.250 55.300 19.600 ;
      LAYER met1 ;
        RECT 55.300 19.250 57.750 19.600 ;
        RECT 46.900 18.900 53.900 19.250 ;
      LAYER met1 ;
        RECT 53.900 18.900 55.650 19.250 ;
        RECT 45.850 18.550 46.550 18.900 ;
      LAYER met1 ;
        RECT 46.550 18.550 54.250 18.900 ;
      LAYER met1 ;
        RECT 54.250 18.550 55.650 18.900 ;
      LAYER met1 ;
        RECT 13.300 18.200 15.750 18.550 ;
      LAYER met1 ;
        RECT 15.750 18.200 17.850 18.550 ;
      LAYER met1 ;
        RECT 17.850 18.200 43.400 18.550 ;
        RECT 13.300 17.850 15.400 18.200 ;
      LAYER met1 ;
        RECT 15.400 17.850 17.500 18.200 ;
      LAYER met1 ;
        RECT 17.500 17.850 43.400 18.200 ;
      LAYER met1 ;
        RECT 43.400 17.850 44.800 18.550 ;
      LAYER met1 ;
        RECT 13.300 17.500 15.050 17.850 ;
      LAYER met1 ;
        RECT 15.050 17.500 17.150 17.850 ;
      LAYER met1 ;
        RECT 17.150 17.500 43.750 17.850 ;
      LAYER met1 ;
        RECT 43.750 17.500 44.800 17.850 ;
      LAYER met1 ;
        RECT 44.800 17.500 45.500 18.550 ;
      LAYER met1 ;
        RECT 45.500 18.200 46.550 18.550 ;
      LAYER met1 ;
        RECT 46.550 18.200 54.600 18.550 ;
      LAYER met1 ;
        RECT 54.600 18.200 55.650 18.550 ;
      LAYER met1 ;
        RECT 55.650 18.200 57.750 19.250 ;
      LAYER met1 ;
        RECT 45.500 17.500 46.200 18.200 ;
      LAYER met1 ;
        RECT 46.200 17.850 54.600 18.200 ;
      LAYER met1 ;
        RECT 54.600 17.850 56.000 18.200 ;
      LAYER met1 ;
        RECT 56.000 17.850 57.750 18.200 ;
        RECT 13.300 17.150 14.700 17.500 ;
      LAYER met1 ;
        RECT 14.700 17.150 16.800 17.500 ;
      LAYER met1 ;
        RECT 16.800 17.150 43.750 17.500 ;
      LAYER met1 ;
        RECT 43.750 17.150 46.200 17.500 ;
      LAYER met1 ;
        RECT 46.200 17.150 50.400 17.850 ;
      LAYER met1 ;
        RECT 50.400 17.500 50.750 17.850 ;
      LAYER met1 ;
        RECT 50.750 17.500 54.600 17.850 ;
      LAYER met1 ;
        RECT 50.400 17.150 51.100 17.500 ;
      LAYER met1 ;
        RECT 51.100 17.150 54.600 17.500 ;
        RECT 13.300 16.800 14.350 17.150 ;
      LAYER met1 ;
        RECT 14.350 16.800 16.450 17.150 ;
      LAYER met1 ;
        RECT 16.450 16.800 43.750 17.150 ;
      LAYER met1 ;
        RECT 43.750 16.800 45.850 17.150 ;
      LAYER met1 ;
        RECT 0.000 15.400 4.550 15.750 ;
      LAYER met1 ;
        RECT 4.550 15.400 13.300 15.750 ;
      LAYER met1 ;
        RECT 13.300 15.400 14.000 16.800 ;
      LAYER met1 ;
        RECT 14.000 16.450 16.100 16.800 ;
      LAYER met1 ;
        RECT 16.100 16.450 44.100 16.800 ;
      LAYER met1 ;
        RECT 14.000 16.100 15.750 16.450 ;
      LAYER met1 ;
        RECT 15.750 16.100 44.100 16.450 ;
      LAYER met1 ;
        RECT 44.100 16.100 45.850 16.800 ;
      LAYER met1 ;
        RECT 45.850 16.100 50.400 17.150 ;
      LAYER met1 ;
        RECT 50.400 16.800 51.450 17.150 ;
      LAYER met1 ;
        RECT 51.450 16.800 54.600 17.150 ;
      LAYER met1 ;
        RECT 54.600 16.800 55.650 17.850 ;
      LAYER met1 ;
        RECT 55.650 16.800 57.750 17.850 ;
      LAYER met1 ;
        RECT 50.400 16.450 51.800 16.800 ;
      LAYER met1 ;
        RECT 51.800 16.450 54.250 16.800 ;
      LAYER met1 ;
        RECT 54.250 16.450 55.300 16.800 ;
      LAYER met1 ;
        RECT 55.300 16.450 57.750 16.800 ;
      LAYER met1 ;
        RECT 57.750 16.450 59.150 23.450 ;
      LAYER met1 ;
        RECT 59.150 23.100 65.100 23.450 ;
      LAYER met1 ;
        RECT 65.100 23.100 66.500 23.450 ;
      LAYER met1 ;
        RECT 66.500 23.100 68.600 23.450 ;
      LAYER met1 ;
        RECT 68.600 23.100 70.000 23.450 ;
      LAYER met1 ;
        RECT 59.150 22.400 64.750 23.100 ;
      LAYER met1 ;
        RECT 64.750 22.750 66.150 23.100 ;
      LAYER met1 ;
        RECT 66.150 22.750 68.950 23.100 ;
      LAYER met1 ;
        RECT 68.950 22.750 70.000 23.100 ;
      LAYER met1 ;
        RECT 70.000 22.750 73.150 23.450 ;
      LAYER met1 ;
        RECT 64.750 22.400 65.800 22.750 ;
      LAYER met1 ;
        RECT 65.800 22.400 73.150 22.750 ;
        RECT 59.150 22.050 64.400 22.400 ;
      LAYER met1 ;
        RECT 64.400 22.050 65.450 22.400 ;
      LAYER met1 ;
        RECT 59.150 21.000 64.050 22.050 ;
      LAYER met1 ;
        RECT 64.050 21.700 65.450 22.050 ;
      LAYER met1 ;
        RECT 65.450 21.700 73.150 22.400 ;
      LAYER met1 ;
        RECT 64.050 21.000 65.100 21.700 ;
      LAYER met1 ;
        RECT 59.150 18.200 63.700 21.000 ;
      LAYER met1 ;
        RECT 63.700 18.200 65.100 21.000 ;
      LAYER met1 ;
        RECT 65.100 18.200 73.150 21.700 ;
        RECT 59.150 17.500 64.050 18.200 ;
      LAYER met1 ;
        RECT 64.050 17.500 65.450 18.200 ;
      LAYER met1 ;
        RECT 65.450 17.500 73.150 18.200 ;
        RECT 59.150 16.800 62.650 17.500 ;
      LAYER met1 ;
        RECT 62.650 16.800 63.000 17.500 ;
      LAYER met1 ;
        RECT 63.000 16.800 64.400 17.500 ;
      LAYER met1 ;
        RECT 64.400 17.150 65.800 17.500 ;
      LAYER met1 ;
        RECT 65.800 17.150 73.150 17.500 ;
      LAYER met1 ;
        RECT 64.400 16.800 66.150 17.150 ;
      LAYER met1 ;
        RECT 66.150 16.800 69.650 17.150 ;
      LAYER met1 ;
        RECT 69.650 16.800 70.350 17.150 ;
      LAYER met1 ;
        RECT 70.350 16.800 73.150 17.150 ;
        RECT 59.150 16.450 62.300 16.800 ;
      LAYER met1 ;
        RECT 62.300 16.450 63.000 16.800 ;
      LAYER met1 ;
        RECT 63.000 16.450 64.750 16.800 ;
      LAYER met1 ;
        RECT 64.750 16.450 66.500 16.800 ;
      LAYER met1 ;
        RECT 66.500 16.450 68.950 16.800 ;
      LAYER met1 ;
        RECT 68.950 16.450 70.000 16.800 ;
      LAYER met1 ;
        RECT 70.000 16.450 73.150 16.800 ;
      LAYER met1 ;
        RECT 50.400 16.100 52.500 16.450 ;
      LAYER met1 ;
        RECT 52.500 16.100 53.550 16.450 ;
      LAYER met1 ;
        RECT 53.550 16.100 54.950 16.450 ;
      LAYER met1 ;
        RECT 54.950 16.100 57.750 16.450 ;
      LAYER met1 ;
        RECT 57.750 16.100 59.500 16.450 ;
      LAYER met1 ;
        RECT 59.500 16.100 61.950 16.450 ;
      LAYER met1 ;
        RECT 61.950 16.100 63.000 16.450 ;
      LAYER met1 ;
        RECT 63.000 16.100 65.100 16.450 ;
      LAYER met1 ;
        RECT 65.100 16.100 67.550 16.450 ;
      LAYER met1 ;
        RECT 67.550 16.100 67.900 16.450 ;
      LAYER met1 ;
        RECT 67.900 16.100 69.650 16.450 ;
      LAYER met1 ;
        RECT 69.650 16.100 73.150 16.450 ;
      LAYER met1 ;
        RECT 14.000 15.750 15.400 16.100 ;
      LAYER met1 ;
        RECT 15.400 15.750 44.450 16.100 ;
      LAYER met1 ;
        RECT 44.450 15.750 45.500 16.100 ;
      LAYER met1 ;
        RECT 45.500 15.750 50.750 16.100 ;
      LAYER met1 ;
        RECT 50.750 15.750 54.600 16.100 ;
      LAYER met1 ;
        RECT 54.600 15.750 57.050 16.100 ;
      LAYER met1 ;
        RECT 57.050 15.750 63.000 16.100 ;
      LAYER met1 ;
        RECT 63.000 15.750 65.450 16.100 ;
      LAYER met1 ;
        RECT 65.450 15.750 68.950 16.100 ;
      LAYER met1 ;
        RECT 68.950 15.750 73.150 16.100 ;
      LAYER met1 ;
        RECT 14.000 15.400 14.700 15.750 ;
      LAYER met1 ;
        RECT 14.700 15.400 44.450 15.750 ;
      LAYER met1 ;
        RECT 44.450 15.400 45.150 15.750 ;
      LAYER met1 ;
        RECT 45.150 15.400 51.450 15.750 ;
      LAYER met1 ;
        RECT 51.450 15.400 53.900 15.750 ;
      LAYER met1 ;
        RECT 53.900 15.400 56.700 15.750 ;
      LAYER met1 ;
        RECT 56.700 15.400 62.650 15.750 ;
      LAYER met1 ;
        RECT 62.650 15.400 66.150 15.750 ;
      LAYER met1 ;
        RECT 66.150 15.400 68.600 15.750 ;
      LAYER met1 ;
        RECT 68.600 15.400 73.150 15.750 ;
        RECT 0.000 15.050 5.250 15.400 ;
      LAYER met1 ;
        RECT 5.250 15.050 13.300 15.400 ;
      LAYER met1 ;
        RECT 0.000 14.700 5.950 15.050 ;
      LAYER met1 ;
        RECT 5.950 14.700 13.300 15.050 ;
      LAYER met1 ;
        RECT 13.300 14.700 73.150 15.400 ;
        RECT 0.000 14.350 7.000 14.700 ;
      LAYER met1 ;
        RECT 7.000 14.350 12.600 14.700 ;
      LAYER met1 ;
        RECT 12.600 14.350 73.150 14.700 ;
        RECT 0.000 14.000 8.750 14.350 ;
      LAYER met1 ;
        RECT 8.750 14.000 10.850 14.350 ;
      LAYER met1 ;
        RECT 10.850 14.000 73.150 14.350 ;
        RECT 0.000 13.650 28.350 14.000 ;
      LAYER met1 ;
        RECT 28.350 13.650 31.150 14.000 ;
      LAYER met1 ;
        RECT 0.000 11.550 28.000 13.650 ;
      LAYER met1 ;
        RECT 28.000 12.950 31.150 13.650 ;
      LAYER met1 ;
        RECT 31.150 12.950 43.750 14.000 ;
      LAYER met1 ;
        RECT 28.000 11.550 29.050 12.950 ;
      LAYER met1 ;
        RECT 29.050 11.900 30.450 12.950 ;
      LAYER met1 ;
        RECT 30.450 11.900 31.150 12.950 ;
      LAYER met1 ;
        RECT 29.050 11.550 30.100 11.900 ;
      LAYER met1 ;
        RECT 30.100 11.550 31.150 11.900 ;
      LAYER met1 ;
        RECT 0.000 11.200 1.750 11.550 ;
      LAYER met1 ;
        RECT 1.750 11.200 6.300 11.550 ;
      LAYER met1 ;
        RECT 6.300 11.200 7.350 11.550 ;
        RECT 0.000 10.150 1.400 11.200 ;
      LAYER met1 ;
        RECT 1.400 10.150 6.650 11.200 ;
      LAYER met1 ;
        RECT 6.650 10.150 7.350 11.200 ;
      LAYER met1 ;
        RECT 7.350 10.150 12.250 11.550 ;
      LAYER met1 ;
        RECT 12.250 10.150 12.950 11.550 ;
      LAYER met1 ;
        RECT 12.950 11.200 14.000 11.550 ;
      LAYER met1 ;
        RECT 14.000 11.200 28.000 11.550 ;
        RECT 0.000 6.300 4.900 10.150 ;
        RECT 0.000 3.150 1.400 6.300 ;
      LAYER met1 ;
        RECT 1.400 4.550 2.800 6.300 ;
      LAYER met1 ;
        RECT 2.800 4.550 4.900 6.300 ;
      LAYER met1 ;
        RECT 4.900 4.550 6.300 10.150 ;
      LAYER met1 ;
        RECT 6.300 6.300 7.350 10.150 ;
      LAYER met1 ;
        RECT 7.350 7.700 8.750 10.150 ;
      LAYER met1 ;
        RECT 8.750 7.700 12.950 10.150 ;
      LAYER met1 ;
        RECT 12.950 8.750 14.350 11.200 ;
      LAYER met1 ;
        RECT 14.350 10.850 16.800 11.200 ;
      LAYER met1 ;
        RECT 16.800 10.850 17.500 11.200 ;
      LAYER met1 ;
        RECT 17.500 10.850 28.000 11.200 ;
      LAYER met1 ;
        RECT 28.000 10.850 31.150 11.550 ;
      LAYER met1 ;
        RECT 14.350 10.500 16.450 10.850 ;
      LAYER met1 ;
        RECT 16.450 10.500 17.850 10.850 ;
      LAYER met1 ;
        RECT 14.350 10.150 16.100 10.500 ;
      LAYER met1 ;
        RECT 16.100 10.150 17.850 10.500 ;
      LAYER met1 ;
        RECT 17.850 10.150 28.000 10.850 ;
        RECT 14.350 9.800 15.750 10.150 ;
      LAYER met1 ;
        RECT 15.750 9.800 17.500 10.150 ;
      LAYER met1 ;
        RECT 17.500 9.800 28.000 10.150 ;
        RECT 14.350 9.450 15.400 9.800 ;
      LAYER met1 ;
        RECT 15.400 9.450 17.150 9.800 ;
      LAYER met1 ;
        RECT 17.150 9.450 28.000 9.800 ;
        RECT 14.350 9.100 15.050 9.450 ;
      LAYER met1 ;
        RECT 15.050 9.100 16.800 9.450 ;
      LAYER met1 ;
        RECT 16.800 9.100 28.000 9.450 ;
      LAYER met1 ;
        RECT 28.000 9.100 29.050 10.850 ;
      LAYER met1 ;
        RECT 29.050 10.500 30.100 10.850 ;
      LAYER met1 ;
        RECT 30.100 10.500 31.150 10.850 ;
      LAYER met1 ;
        RECT 29.050 9.100 30.450 10.500 ;
      LAYER met1 ;
        RECT 30.450 9.100 31.150 10.500 ;
      LAYER met1 ;
        RECT 31.150 9.100 31.500 12.950 ;
      LAYER met1 ;
        RECT 31.500 12.600 32.200 12.950 ;
      LAYER met1 ;
        RECT 32.200 12.600 33.950 12.950 ;
      LAYER met1 ;
        RECT 33.950 12.600 34.300 12.950 ;
      LAYER met1 ;
        RECT 34.300 12.600 35.000 12.950 ;
      LAYER met1 ;
        RECT 31.500 12.250 32.550 12.600 ;
      LAYER met1 ;
        RECT 32.550 12.250 33.600 12.600 ;
      LAYER met1 ;
        RECT 31.500 11.550 32.900 12.250 ;
      LAYER met1 ;
        RECT 32.900 11.550 33.600 12.250 ;
      LAYER met1 ;
        RECT 31.500 10.850 33.250 11.550 ;
      LAYER met1 ;
        RECT 33.250 10.850 33.600 11.550 ;
      LAYER met1 ;
        RECT 33.600 10.850 34.650 12.600 ;
        RECT 31.500 9.100 32.200 10.850 ;
      LAYER met1 ;
        RECT 32.200 10.500 32.550 10.850 ;
      LAYER met1 ;
        RECT 32.550 10.500 34.650 10.850 ;
      LAYER met1 ;
        RECT 32.200 10.150 32.900 10.500 ;
      LAYER met1 ;
        RECT 32.900 10.150 34.650 10.500 ;
      LAYER met1 ;
        RECT 32.200 9.450 33.250 10.150 ;
      LAYER met1 ;
        RECT 33.250 9.450 34.650 10.150 ;
      LAYER met1 ;
        RECT 32.200 9.100 33.600 9.450 ;
      LAYER met1 ;
        RECT 33.600 9.100 34.650 9.450 ;
      LAYER met1 ;
        RECT 34.650 9.100 35.000 12.600 ;
      LAYER met1 ;
        RECT 35.000 12.250 35.700 12.950 ;
      LAYER met1 ;
        RECT 35.700 12.250 37.100 12.950 ;
      LAYER met1 ;
        RECT 35.000 11.900 36.050 12.250 ;
      LAYER met1 ;
        RECT 36.050 11.900 37.100 12.250 ;
      LAYER met1 ;
        RECT 35.000 11.200 36.400 11.900 ;
      LAYER met1 ;
        RECT 36.400 11.200 37.100 11.900 ;
      LAYER met1 ;
        RECT 35.000 10.850 36.750 11.200 ;
      LAYER met1 ;
        RECT 36.750 10.850 37.100 11.200 ;
      LAYER met1 ;
        RECT 37.100 10.850 37.800 12.950 ;
      LAYER met1 ;
        RECT 37.800 12.600 38.500 12.950 ;
      LAYER met1 ;
        RECT 38.500 12.600 40.950 12.950 ;
      LAYER met1 ;
        RECT 40.950 12.600 43.750 12.950 ;
      LAYER met1 ;
        RECT 35.000 9.100 35.700 10.850 ;
      LAYER met1 ;
        RECT 35.700 10.500 36.050 10.850 ;
      LAYER met1 ;
        RECT 36.050 10.500 37.800 10.850 ;
      LAYER met1 ;
        RECT 35.700 9.800 36.400 10.500 ;
      LAYER met1 ;
        RECT 36.400 9.800 37.800 10.500 ;
      LAYER met1 ;
        RECT 35.700 9.450 36.750 9.800 ;
      LAYER met1 ;
        RECT 36.750 9.450 37.800 9.800 ;
      LAYER met1 ;
        RECT 35.700 9.100 37.100 9.450 ;
      LAYER met1 ;
        RECT 37.100 9.100 37.800 9.450 ;
      LAYER met1 ;
        RECT 37.800 9.100 38.150 12.600 ;
      LAYER met1 ;
        RECT 38.150 11.900 41.300 12.600 ;
        RECT 38.150 11.200 38.850 11.900 ;
      LAYER met1 ;
        RECT 38.850 11.200 40.250 11.900 ;
      LAYER met1 ;
        RECT 40.250 11.200 41.300 11.900 ;
        RECT 38.150 10.500 41.300 11.200 ;
      LAYER met1 ;
        RECT 41.300 10.500 43.750 12.600 ;
      LAYER met1 ;
        RECT 38.150 10.150 39.200 10.500 ;
      LAYER met1 ;
        RECT 39.200 10.150 43.750 10.500 ;
      LAYER met1 ;
        RECT 38.150 9.800 38.850 10.150 ;
      LAYER met1 ;
        RECT 38.850 9.800 43.750 10.150 ;
      LAYER met1 ;
        RECT 38.150 9.100 41.300 9.800 ;
      LAYER met1 ;
        RECT 41.300 9.100 43.750 9.800 ;
      LAYER met1 ;
        RECT 43.750 9.100 44.450 14.000 ;
      LAYER met1 ;
        RECT 44.450 12.950 73.150 14.000 ;
        RECT 44.450 12.600 45.150 12.950 ;
      LAYER met1 ;
        RECT 45.150 12.600 47.950 12.950 ;
      LAYER met1 ;
        RECT 44.450 10.500 44.800 12.600 ;
      LAYER met1 ;
        RECT 44.800 11.900 47.950 12.600 ;
      LAYER met1 ;
        RECT 47.950 11.900 48.650 12.950 ;
      LAYER met1 ;
        RECT 48.650 12.600 51.100 12.950 ;
      LAYER met1 ;
        RECT 51.100 12.600 52.150 12.950 ;
      LAYER met1 ;
        RECT 52.150 12.600 54.600 12.950 ;
      LAYER met1 ;
        RECT 54.600 12.600 55.300 12.950 ;
      LAYER met1 ;
        RECT 55.300 12.600 58.100 12.950 ;
        RECT 48.650 11.900 51.450 12.600 ;
      LAYER met1 ;
        RECT 51.450 11.900 51.800 12.600 ;
      LAYER met1 ;
        RECT 51.800 11.900 54.600 12.600 ;
        RECT 44.800 11.200 45.850 11.900 ;
      LAYER met1 ;
        RECT 45.850 11.200 50.400 11.900 ;
      LAYER met1 ;
        RECT 50.400 11.200 51.450 11.900 ;
      LAYER met1 ;
        RECT 51.450 11.200 53.900 11.900 ;
      LAYER met1 ;
        RECT 53.900 11.200 54.600 11.900 ;
        RECT 44.800 10.500 47.950 11.200 ;
      LAYER met1 ;
        RECT 44.450 9.800 47.250 10.500 ;
      LAYER met1 ;
        RECT 47.250 9.800 47.950 10.500 ;
      LAYER met1 ;
        RECT 44.450 9.100 44.800 9.800 ;
      LAYER met1 ;
        RECT 44.800 9.100 47.950 9.800 ;
      LAYER met1 ;
        RECT 47.950 9.100 48.300 11.200 ;
      LAYER met1 ;
        RECT 48.300 10.850 51.450 11.200 ;
      LAYER met1 ;
        RECT 51.450 10.850 51.800 11.200 ;
      LAYER met1 ;
        RECT 51.800 10.850 54.600 11.200 ;
        RECT 48.300 10.500 54.600 10.850 ;
        RECT 48.300 9.800 49.000 10.500 ;
      LAYER met1 ;
        RECT 49.000 9.800 50.400 10.500 ;
      LAYER met1 ;
        RECT 50.400 9.800 52.500 10.500 ;
      LAYER met1 ;
        RECT 52.500 9.800 53.900 10.500 ;
      LAYER met1 ;
        RECT 53.900 9.800 54.600 10.500 ;
        RECT 48.300 9.100 54.600 9.800 ;
      LAYER met1 ;
        RECT 54.600 9.100 54.950 12.600 ;
      LAYER met1 ;
        RECT 54.950 11.900 58.100 12.600 ;
      LAYER met1 ;
        RECT 58.100 11.900 73.150 12.950 ;
      LAYER met1 ;
        RECT 54.950 9.800 56.000 11.900 ;
      LAYER met1 ;
        RECT 56.000 9.800 73.150 11.900 ;
      LAYER met1 ;
        RECT 54.950 9.100 58.100 9.800 ;
      LAYER met1 ;
        RECT 58.100 9.100 73.150 9.800 ;
        RECT 14.350 8.750 14.700 9.100 ;
      LAYER met1 ;
        RECT 14.700 8.750 16.450 9.100 ;
        RECT 12.950 8.400 16.450 8.750 ;
      LAYER met1 ;
        RECT 16.450 8.400 73.150 9.100 ;
      LAYER met1 ;
        RECT 12.950 8.050 16.100 8.400 ;
      LAYER met1 ;
        RECT 16.100 8.050 73.150 8.400 ;
      LAYER met1 ;
        RECT 12.950 7.700 15.750 8.050 ;
      LAYER met1 ;
        RECT 15.750 7.700 73.150 8.050 ;
      LAYER met1 ;
        RECT 7.350 6.300 12.250 7.700 ;
      LAYER met1 ;
        RECT 6.300 4.550 10.850 6.300 ;
      LAYER met1 ;
        RECT 10.850 4.550 12.250 6.300 ;
        RECT 1.400 3.150 6.300 4.550 ;
      LAYER met1 ;
        RECT 6.300 3.150 7.350 4.550 ;
      LAYER met1 ;
        RECT 7.350 3.150 12.250 4.550 ;
      LAYER met1 ;
        RECT 12.250 3.150 12.950 7.700 ;
      LAYER met1 ;
        RECT 12.950 7.000 15.400 7.700 ;
      LAYER met1 ;
        RECT 15.400 7.000 73.150 7.700 ;
      LAYER met1 ;
        RECT 12.950 6.300 15.750 7.000 ;
      LAYER met1 ;
        RECT 15.750 6.650 73.150 7.000 ;
        RECT 15.750 6.300 30.800 6.650 ;
      LAYER met1 ;
        RECT 12.950 5.950 16.100 6.300 ;
      LAYER met1 ;
        RECT 16.100 5.950 30.800 6.300 ;
      LAYER met1 ;
        RECT 30.800 5.950 33.950 6.650 ;
        RECT 12.950 3.150 14.350 5.950 ;
      LAYER met1 ;
        RECT 14.350 5.600 14.700 5.950 ;
      LAYER met1 ;
        RECT 14.700 5.600 16.450 5.950 ;
      LAYER met1 ;
        RECT 16.450 5.600 30.800 5.950 ;
        RECT 14.350 5.250 15.050 5.600 ;
      LAYER met1 ;
        RECT 15.050 5.250 16.800 5.600 ;
      LAYER met1 ;
        RECT 16.800 5.250 30.800 5.600 ;
        RECT 14.350 4.900 15.400 5.250 ;
      LAYER met1 ;
        RECT 15.400 4.900 17.150 5.250 ;
      LAYER met1 ;
        RECT 17.150 4.900 30.800 5.250 ;
        RECT 14.350 4.550 15.750 4.900 ;
      LAYER met1 ;
        RECT 15.750 4.550 17.500 4.900 ;
      LAYER met1 ;
        RECT 17.500 4.550 30.800 4.900 ;
      LAYER met1 ;
        RECT 30.800 4.550 31.850 5.950 ;
      LAYER met1 ;
        RECT 31.850 4.550 33.250 5.950 ;
      LAYER met1 ;
        RECT 33.250 4.550 33.950 5.950 ;
      LAYER met1 ;
        RECT 33.950 5.600 54.250 6.650 ;
      LAYER met1 ;
        RECT 54.250 5.600 55.300 6.650 ;
      LAYER met1 ;
        RECT 14.350 4.200 16.100 4.550 ;
      LAYER met1 ;
        RECT 16.100 4.200 17.850 4.550 ;
      LAYER met1 ;
        RECT 14.350 3.850 16.450 4.200 ;
      LAYER met1 ;
        RECT 16.450 3.850 17.850 4.200 ;
      LAYER met1 ;
        RECT 14.350 3.500 16.800 3.850 ;
      LAYER met1 ;
        RECT 16.800 3.500 17.850 3.850 ;
      LAYER met1 ;
        RECT 17.850 3.500 30.800 4.550 ;
      LAYER met1 ;
        RECT 30.800 3.850 33.950 4.550 ;
      LAYER met1 ;
        RECT 33.950 3.850 34.300 5.600 ;
      LAYER met1 ;
        RECT 34.300 4.900 37.450 5.600 ;
        RECT 30.800 3.500 33.250 3.850 ;
      LAYER met1 ;
        RECT 14.350 3.150 30.800 3.500 ;
        RECT 0.000 2.100 30.800 3.150 ;
      LAYER met1 ;
        RECT 30.800 2.100 31.850 3.500 ;
      LAYER met1 ;
        RECT 31.850 3.150 32.200 3.500 ;
      LAYER met1 ;
        RECT 32.200 3.150 33.250 3.500 ;
      LAYER met1 ;
        RECT 33.250 3.150 34.300 3.850 ;
        RECT 31.850 2.800 32.550 3.150 ;
      LAYER met1 ;
        RECT 32.550 2.800 33.600 3.150 ;
      LAYER met1 ;
        RECT 33.600 2.800 34.300 3.150 ;
      LAYER met1 ;
        RECT 34.300 2.800 35.000 4.900 ;
      LAYER met1 ;
        RECT 35.000 2.800 36.400 4.900 ;
      LAYER met1 ;
        RECT 36.400 2.800 37.450 4.900 ;
      LAYER met1 ;
        RECT 37.450 3.150 37.800 5.600 ;
      LAYER met1 ;
        RECT 37.800 4.900 40.600 5.600 ;
      LAYER met1 ;
        RECT 40.600 4.900 41.300 5.600 ;
      LAYER met1 ;
        RECT 41.300 4.900 44.100 5.600 ;
        RECT 37.800 4.200 38.500 4.900 ;
      LAYER met1 ;
        RECT 38.500 4.550 43.050 4.900 ;
      LAYER met1 ;
        RECT 43.050 4.550 44.100 4.900 ;
      LAYER met1 ;
        RECT 38.500 4.200 43.400 4.550 ;
      LAYER met1 ;
        RECT 43.400 4.200 44.100 4.550 ;
        RECT 37.800 3.850 40.600 4.200 ;
      LAYER met1 ;
        RECT 40.600 3.850 40.950 4.200 ;
      LAYER met1 ;
        RECT 40.950 3.850 44.100 4.200 ;
        RECT 37.800 3.150 44.100 3.850 ;
      LAYER met1 ;
        RECT 37.450 2.800 39.900 3.150 ;
      LAYER met1 ;
        RECT 39.900 2.800 42.000 3.150 ;
      LAYER met1 ;
        RECT 42.000 2.800 43.400 3.150 ;
      LAYER met1 ;
        RECT 43.400 2.800 44.100 3.150 ;
      LAYER met1 ;
        RECT 31.850 2.450 32.900 2.800 ;
      LAYER met1 ;
        RECT 32.900 2.450 33.950 2.800 ;
      LAYER met1 ;
        RECT 31.850 2.100 33.250 2.450 ;
      LAYER met1 ;
        RECT 33.250 2.100 33.950 2.450 ;
      LAYER met1 ;
        RECT 33.950 2.100 34.300 2.800 ;
      LAYER met1 ;
        RECT 34.300 2.100 37.450 2.800 ;
      LAYER met1 ;
        RECT 37.450 2.100 37.800 2.800 ;
      LAYER met1 ;
        RECT 37.800 2.100 44.100 2.800 ;
      LAYER met1 ;
        RECT 44.100 2.100 44.450 5.600 ;
      LAYER met1 ;
        RECT 44.450 2.800 45.150 5.600 ;
      LAYER met1 ;
        RECT 45.150 2.800 47.600 5.600 ;
        RECT 0.000 1.750 31.150 2.100 ;
      LAYER met1 ;
        RECT 31.150 1.750 31.500 2.100 ;
      LAYER met1 ;
        RECT 31.500 1.750 34.300 2.100 ;
      LAYER met1 ;
        RECT 34.300 1.750 37.100 2.100 ;
      LAYER met1 ;
        RECT 37.100 1.750 37.800 2.100 ;
      LAYER met1 ;
        RECT 37.800 1.750 40.600 2.100 ;
      LAYER met1 ;
        RECT 40.600 1.750 41.300 2.100 ;
      LAYER met1 ;
        RECT 41.300 1.750 43.750 2.100 ;
      LAYER met1 ;
        RECT 43.750 1.750 44.450 2.100 ;
      LAYER met1 ;
        RECT 44.450 1.750 47.250 2.800 ;
      LAYER met1 ;
        RECT 47.250 2.100 47.600 2.800 ;
      LAYER met1 ;
        RECT 47.600 2.100 48.300 5.600 ;
      LAYER met1 ;
        RECT 48.300 2.100 48.650 5.600 ;
      LAYER met1 ;
        RECT 48.650 5.250 49.700 5.600 ;
      LAYER met1 ;
        RECT 49.700 5.250 51.100 5.600 ;
      LAYER met1 ;
        RECT 48.650 4.550 50.050 5.250 ;
      LAYER met1 ;
        RECT 50.050 4.550 51.100 5.250 ;
      LAYER met1 ;
        RECT 48.650 4.200 50.400 4.550 ;
      LAYER met1 ;
        RECT 50.400 4.200 51.100 4.550 ;
      LAYER met1 ;
        RECT 48.650 3.850 50.750 4.200 ;
      LAYER met1 ;
        RECT 50.750 3.850 51.100 4.200 ;
      LAYER met1 ;
        RECT 51.100 3.850 51.800 5.600 ;
        RECT 48.650 2.100 49.700 3.850 ;
      LAYER met1 ;
        RECT 49.700 3.150 50.050 3.850 ;
      LAYER met1 ;
        RECT 50.050 3.150 51.800 3.850 ;
      LAYER met1 ;
        RECT 49.700 2.800 50.400 3.150 ;
      LAYER met1 ;
        RECT 50.400 2.800 51.800 3.150 ;
      LAYER met1 ;
        RECT 49.700 2.100 50.750 2.800 ;
      LAYER met1 ;
        RECT 50.750 2.100 51.800 2.800 ;
      LAYER met1 ;
        RECT 47.250 1.750 47.950 2.100 ;
      LAYER met1 ;
        RECT 47.950 1.750 48.300 2.100 ;
      LAYER met1 ;
        RECT 48.300 1.750 49.000 2.100 ;
      LAYER met1 ;
        RECT 49.000 1.750 49.350 2.100 ;
      LAYER met1 ;
        RECT 49.350 1.750 51.100 2.100 ;
      LAYER met1 ;
        RECT 51.100 1.750 51.800 2.100 ;
      LAYER met1 ;
        RECT 51.800 1.750 52.150 5.600 ;
      LAYER met1 ;
        RECT 52.150 4.900 55.300 5.600 ;
        RECT 52.150 2.800 52.850 4.900 ;
      LAYER met1 ;
        RECT 52.850 2.800 54.250 4.900 ;
      LAYER met1 ;
        RECT 54.250 2.800 55.300 4.900 ;
        RECT 52.150 2.100 55.300 2.800 ;
      LAYER met1 ;
        RECT 55.300 2.100 73.150 6.650 ;
      LAYER met1 ;
        RECT 52.150 1.750 54.950 2.100 ;
      LAYER met1 ;
        RECT 54.950 1.750 73.150 2.100 ;
        RECT 0.000 0.000 73.150 1.750 ;
  END
END my_logo
END LIBRARY

