* NGSPICE file created from tt_um_jimktrains_vslc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt tt_um_jimktrains_vslc VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_0_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1270_ _1516_/Q _1270_/B VGND VGND VPWR VPWR _1270_/X sky130_fd_sc_hd__and2b_1
Xwire18 wire18/A VGND VGND VPWR VPWR wire18/X sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0985_ _1622_/Q _0985_/B VGND VGND VPWR VPWR _0986_/B sky130_fd_sc_hd__xnor2_1
X_1606_ _1606_/CLK _1606_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
X_1537_ _1541_/CLK input5/X VGND VGND VPWR VPWR _1537_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1450__86 _1454__90/A VGND VGND VPWR VPWR _1602_/CLK sky130_fd_sc_hd__inv_2
X_0770_ hold18/A VGND VGND VPWR VPWR _0770_/Y sky130_fd_sc_hd__inv_2
X_1253_ hold57/A hold51/A _1547_/Q VGND VGND VPWR VPWR _1253_/X sky130_fd_sc_hd__mux2_1
X_1322_ _1519_/Q _1322_/B VGND VGND VPWR VPWR _1322_/X sky130_fd_sc_hd__or2_1
X_1184_ hold42/X _1550_/Q _1184_/S VGND VGND VPWR VPWR _1550_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1372__8/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0968_ _0940_/A _1624_/Q _0963_/Y wire17/X _1149_/A VGND VGND VPWR VPWR _0969_/B
+ sky130_fd_sc_hd__a32o_1
X_0899_ hold36/A _0984_/B _1030_/B VGND VGND VPWR VPWR _0899_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ _0831_/B _0822_/B _0822_/C _0832_/C VGND VGND VPWR VPWR _0825_/C sky130_fd_sc_hd__or4_1
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1236_ _1236_/A _1236_/B _1236_/C _1130_/D VGND VGND VPWR VPWR _1236_/X sky130_fd_sc_hd__or4b_1
X_1305_ _1178_/S _1304_/X _1303_/X _1276_/X VGND VGND VPWR VPWR _1305_/X sky130_fd_sc_hd__a211o_1
X_1167_ _1201_/B _1352_/A uo_out[6] VGND VGND VPWR VPWR _1167_/X sky130_fd_sc_hd__a21o_1
X_1098_ _1577_/Q _1104_/B VGND VGND VPWR VPWR _1098_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1420__56 clkload6/A VGND VGND VPWR VPWR _1572_/CLK sky130_fd_sc_hd__inv_2
X_1021_ hold29/A _1592_/Q _1593_/Q _1594_/Q VGND VGND VPWR VPWR _1023_/D sky130_fd_sc_hd__and4_1
X_0805_ hold37/A _1655_/Q VGND VGND VPWR VPWR _0823_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1219_ _1581_/Q _0766_/Y _1217_/X _1218_/X VGND VGND VPWR VPWR _1221_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1570_ _1570_/CLK _1570_/D VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1004_ _1614_/Q _1004_/B VGND VGND VPWR VPWR _1005_/B sky130_fd_sc_hd__or2_1
X_1368__4 _1533_/CLK VGND VGND VPWR VPWR _1511_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ _1622_/CLK _1622_/D VGND VGND VPWR VPWR _1622_/Q sky130_fd_sc_hd__dfxtp_1
X_1553_ _1553_/CLK _1553_/D VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfxtp_1
X_1456__92 clkload9/A VGND VGND VPWR VPWR _1608_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1490__126 clkload2/A VGND VGND VPWR VPWR _1642_/CLK sky130_fd_sc_hd__inv_2
Xwire19 wire19/A VGND VGND VPWR VPWR wire19/X sky130_fd_sc_hd__buf_2
X_0984_ _1030_/B _0984_/B VGND VGND VPWR VPWR _0984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1536_ _1541_/CLK input4/X VGND VGND VPWR VPWR _1536_/Q sky130_fd_sc_hd__dfxtp_1
X_1605_ _1605_/CLK _1605_/D VGND VGND VPWR VPWR _1605_/Q sky130_fd_sc_hd__dfxtp_1
X_1381__17 clkload13/A VGND VGND VPWR VPWR _1524_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1321_ _1521_/Q _1345_/A2 _1320_/X _1336_/C1 VGND VGND VPWR VPWR _1521_/D sky130_fd_sc_hd__o211a_1
X_1252_ hold45/A hold56/A _1547_/Q VGND VGND VPWR VPWR _1252_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1183_ _1188_/A hold55/X _1184_/S VGND VGND VPWR VPWR _1551_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_6_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0967_ _0971_/A _0967_/B VGND VGND VPWR VPWR _1625_/D sky130_fd_sc_hd__and2_1
X_1426__62 clkload2/A VGND VGND VPWR VPWR _1578_/CLK sky130_fd_sc_hd__inv_2
X_1519_ _1519_/CLK _1519_/D VGND VGND VPWR VPWR _1519_/Q sky130_fd_sc_hd__dfxtp_1
X_0898_ _1248_/A _0897_/X _1030_/A VGND VGND VPWR VPWR _0984_/B sky130_fd_sc_hd__a21boi_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0821_ _0757_/Y _1655_/Q _1611_/Q _0807_/B VGND VGND VPWR VPWR _0832_/C sky130_fd_sc_hd__a2bb2o_1
X_1496__132 clkload10/A VGND VGND VPWR VPWR _1648_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1166_ _1201_/B _1352_/A VGND VGND VPWR VPWR _1166_/Y sky130_fd_sc_hd__nand2_1
X_1235_ _1235_/A _1235_/B VGND VGND VPWR VPWR _1236_/C sky130_fd_sc_hd__nor2_1
X_1304_ hold52/A hold46/A _1339_/S VGND VGND VPWR VPWR _1304_/X sky130_fd_sc_hd__mux2_1
X_1097_ _1076_/A _1089_/X _1096_/X _0845_/A VGND VGND VPWR VPWR _1578_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1020_ hold29/A _1592_/Q _1593_/Q VGND VGND VPWR VPWR _1057_/A sky130_fd_sc_hd__nand3_1
Xclkbuf_4_11_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload10/A sky130_fd_sc_hd__clkbuf_8
X_0804_ _1619_/Q hold20/A VGND VGND VPWR VPWR _0832_/A sky130_fd_sc_hd__and2b_1
X_1149_ _1149_/A _1349_/B VGND VGND VPWR VPWR _1358_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1218_ _1581_/Q _0766_/Y _1136_/A _1580_/Q VGND VGND VPWR VPWR _1218_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1003_ _1615_/Q _1002_/X _1019_/C _0993_/B VGND VGND VPWR VPWR _1615_/D sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1387__23 _1372__8/A VGND VGND VPWR VPWR _1530_/CLK sky130_fd_sc_hd__inv_2
X_1621_ _1621_/CLK _1621_/D VGND VGND VPWR VPWR _1621_/Q sky130_fd_sc_hd__dfxtp_1
X_1552_ _1552_/CLK hold13/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1370__6 _1533_/CLK VGND VGND VPWR VPWR _1513_/CLK sky130_fd_sc_hd__inv_2
X_0983_ _1621_/Q _0983_/B VGND VGND VPWR VPWR _0985_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1535_ _1541_/CLK input3/X VGND VGND VPWR VPWR _1535_/Q sky130_fd_sc_hd__dfxtp_1
X_1604_ _1604_/CLK _1604_/D VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ _1340_/A1 _1319_/X _1318_/X _1344_/C1 VGND VGND VPWR VPWR _1320_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1182_ hold54/A hold12/X _1184_/S VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__mux2_1
X_1251_ _1251_/A _1251_/B _1251_/C VGND VGND VPWR VPWR _1532_/D sky130_fd_sc_hd__and3_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1441__77 clkload1/A VGND VGND VPWR VPWR _1593_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_6_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0966_ _0940_/A _1625_/Q _0963_/Y wire17/X _1201_/B VGND VGND VPWR VPWR _0967_/B
+ sky130_fd_sc_hd__a32o_1
X_0897_ _0897_/A _0897_/B _0896_/X VGND VGND VPWR VPWR _0897_/X sky130_fd_sc_hd__or3b_1
X_1518_ _1518_/CLK _1518_/D VGND VGND VPWR VPWR _1518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ _0834_/A _0834_/B _0834_/C VGND VGND VPWR VPWR _0822_/C sky130_fd_sc_hd__or3_1
X_1303_ hold52/A _0913_/Y _1333_/B1 _1302_/X VGND VGND VPWR VPWR _1303_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1234_ _1234_/A _1234_/B VGND VGND VPWR VPWR _1236_/B sky130_fd_sc_hd__and2_1
X_1165_ uo_out[7] _1179_/S _1164_/X _1161_/X _1180_/A VGND VGND VPWR VPWR _1557_/D
+ sky130_fd_sc_hd__o221a_1
X_1096_ _1578_/Q _1104_/B VGND VGND VPWR VPWR _1096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0949_ _0956_/A _0949_/B VGND VGND VPWR VPWR _1633_/D sky130_fd_sc_hd__and2_1
XFILLER_0_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1504__140 clkload8/A VGND VGND VPWR VPWR _1656_/CLK sky130_fd_sc_hd__inv_2
X_0803_ _1648_/Q _1610_/Q VGND VGND VPWR VPWR _0834_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1411__47 clkload0/A VGND VGND VPWR VPWR _1563_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1148_ _1162_/A _1148_/B _1162_/B _1162_/C VGND VGND VPWR VPWR _1148_/X sky130_fd_sc_hd__or4bb_1
X_1079_ _1076_/A _1192_/A _1078_/X _1117_/C1 VGND VGND VPWR VPWR _1586_/D sky130_fd_sc_hd__o211a_1
X_1217_ _1214_/X _1215_/X _1216_/X VGND VGND VPWR VPWR _1217_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1002_ _1614_/Q _1004_/B VGND VGND VPWR VPWR _1002_/X sky130_fd_sc_hd__and2_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload9/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ _1620_/CLK _1620_/D VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
X_1551_ _1551_/CLK _1551_/D VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1447__83 _1454__90/A VGND VGND VPWR VPWR _1599_/CLK sky130_fd_sc_hd__inv_2
X_0982_ _0983_/B VGND VGND VPWR VPWR _0982_/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1534_ _1541_/CLK input2/X VGND VGND VPWR VPWR _1534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1603_ _1603_/CLK _1603_/D VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1181_ _1546_/Q hold3/X _1184_/S VGND VGND VPWR VPWR _1553_/D sky130_fd_sc_hd__mux2_1
X_1250_ _1676_/A _0826_/X _0984_/B _1248_/X VGND VGND VPWR VPWR _1251_/C sky130_fd_sc_hd__o211ai_1
XFILLER_0_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0896_ _0888_/X _0891_/X _0896_/C _0896_/D VGND VGND VPWR VPWR _0896_/X sky130_fd_sc_hd__and4bb_1
X_0965_ _0971_/A _0965_/B VGND VGND VPWR VPWR _1626_/D sky130_fd_sc_hd__and2_1
X_1517_ _1517_/CLK _1517_/D VGND VGND VPWR VPWR _1517_/Q sky130_fd_sc_hd__dfxtp_1
X_1480__116 clkload9/A VGND VGND VPWR VPWR _1632_/CLK sky130_fd_sc_hd__inv_2
X_1417__53 clkload6/A VGND VGND VPWR VPWR _1569_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1302_ hold46/A _1322_/B VGND VGND VPWR VPWR _1302_/X sky130_fd_sc_hd__or2_1
X_1233_ hold54/X _1130_/D _1232_/X _1199_/A VGND VGND VPWR VPWR _1545_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1164_ _1260_/A _1342_/C1 _1179_/S VGND VGND VPWR VPWR _1164_/X sky130_fd_sc_hd__a21bo_1
X_1095_ _1162_/B _1089_/X _1094_/X _0971_/A VGND VGND VPWR VPWR _1579_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0948_ _0955_/A1 _1633_/Q _0945_/Y _0945_/B _1148_/B VGND VGND VPWR VPWR _0949_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0879_ _0876_/Y _0877_/X _0878_/X _0875_/X VGND VGND VPWR VPWR _0879_/X sky130_fd_sc_hd__a211o_1
X_0802_ _0802_/A _1651_/Q VGND VGND VPWR VPWR _0830_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1216_ _1580_/Q _1136_/A _0768_/Y _1579_/Q VGND VGND VPWR VPWR _1216_/X sky130_fd_sc_hd__a22o_1
X_1147_ _1149_/A _1349_/B VGND VGND VPWR VPWR _1147_/Y sky130_fd_sc_hd__nand2_1
X_1078_ _1260_/A _1086_/B VGND VGND VPWR VPWR _1078_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
X_1486__122 clkload2/A VGND VGND VPWR VPWR _1638_/CLK sky130_fd_sc_hd__inv_2
Xhold33 hold58/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1001_ _1613_/Q _1612_/Q _1008_/B VGND VGND VPWR VPWR _1004_/B sky130_fd_sc_hd__and3_1
XFILLER_0_12_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1378__14 _1541_/CLK VGND VGND VPWR VPWR _1521_/CLK sky130_fd_sc_hd__inv_2
X_1550_ _1550_/CLK _1550_/D VGND VGND VPWR VPWR _1550_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1462__98 clkload9/A VGND VGND VPWR VPWR _1614_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ hold24/A _1619_/Q hold48/A _0981_/D VGND VGND VPWR VPWR _0983_/B sky130_fd_sc_hd__and4_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1602_ _1602_/CLK _1602_/D VGND VGND VPWR VPWR _1602_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1533_ _1533_/CLK _1533_/D VGND VGND VPWR VPWR _1533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ _1180_/A _1180_/B VGND VGND VPWR VPWR _1554_/D sky130_fd_sc_hd__and2_1
X_0964_ _0940_/A _1626_/Q _0963_/Y wire17/X _1260_/A VGND VGND VPWR VPWR _0965_/B
+ sky130_fd_sc_hd__a32o_1
X_1516_ _1516_/CLK _1516_/D VGND VGND VPWR VPWR _1516_/Q sky130_fd_sc_hd__dfxtp_1
X_0895_ _0757_/Y _1637_/Q _0776_/Y _1621_/Q _0894_/Y VGND VGND VPWR VPWR _0896_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1432__68 clkload10/A VGND VGND VPWR VPWR _1584_/CLK sky130_fd_sc_hd__inv_2
X_1232_ _1203_/Y _1221_/X _1226_/Y _1230_/X _1231_/Y VGND VGND VPWR VPWR _1232_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1301_ hold52/X _1275_/Y _1300_/X _1336_/C1 VGND VGND VPWR VPWR _1525_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ _1260_/A _1339_/S _1061_/Y _1162_/X VGND VGND VPWR VPWR _1179_/S sky130_fd_sc_hd__o211a_2
X_1094_ _1579_/Q _1104_/B VGND VGND VPWR VPWR _1094_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ _0956_/A _0947_/B VGND VGND VPWR VPWR _1634_/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ _1622_/Q _1642_/Q VGND VGND VPWR VPWR _0878_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 clkload0/A VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_6
XPHY_EDGE_ROW_28_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0801_ _1650_/Q _1612_/Q VGND VGND VPWR VPWR _0823_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1215_ _1579_/Q _0768_/Y _1139_/A _1578_/Q VGND VGND VPWR VPWR _1215_/X sky130_fd_sc_hd__o22a_1
X_1146_ _1146_/A _1146_/B VGND VGND VPWR VPWR _1558_/D sky130_fd_sc_hd__nor2_1
X_1077_ _1162_/B _1192_/A _1076_/X _1117_/C1 VGND VGND VPWR VPWR _1587_/D sky130_fd_sc_hd__o211a_1
X_1402__38 clkload6/A VGND VGND VPWR VPWR _1554_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1000_ _1612_/Q _1611_/Q _1010_/B VGND VGND VPWR VPWR _1006_/B sky130_fd_sc_hd__and3_1
XFILLER_0_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1129_ _1199_/A _1130_/D VGND VGND VPWR VPWR _1184_/S sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1393__29 clkload4/A VGND VGND VPWR VPWR _1545_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _1619_/Q hold48/A _0981_/D VGND VGND VPWR VPWR _0980_/X sky130_fd_sc_hd__and3_1
X_1438__74 _1372__8/A VGND VGND VPWR VPWR _1590_/CLK sky130_fd_sc_hd__inv_2
X_1601_ _1601_/CLK _1601_/D VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1532_ _1532_/CLK _1532_/D VGND VGND VPWR VPWR _1676_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0894_ _1619_/Q _1639_/Q VGND VGND VPWR VPWR _0894_/Y sky130_fd_sc_hd__xnor2_1
X_0963_ _0963_/A wire17/A VGND VGND VPWR VPWR _0963_/Y sky130_fd_sc_hd__nor2_1
X_1515_ _1515_/CLK _1515_/D VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1408__44 clkload3/A VGND VGND VPWR VPWR _1560_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1231_ _1257_/B _1231_/B VGND VGND VPWR VPWR _1231_/Y sky130_fd_sc_hd__nor2_1
X_1162_ _1162_/A _1162_/B _1162_/C VGND VGND VPWR VPWR _1162_/X sky130_fd_sc_hd__or3_1
X_1300_ _1159_/Y _1299_/X _1298_/X _1276_/X VGND VGND VPWR VPWR _1300_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1093_ _1072_/A _1089_/X _1092_/X _0971_/A VGND VGND VPWR VPWR _1580_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_22_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0877_ _1608_/Q _1628_/Q VGND VGND VPWR VPWR _0877_/X sky130_fd_sc_hd__or2_1
X_0946_ _0955_/A1 _1634_/Q _0945_/Y _0945_/B _1162_/A VGND VGND VPWR VPWR _0947_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload1 clkload1/A VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_4
XFILLER_0_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0800_ hold48/A _1656_/Q VGND VGND VPWR VPWR _0835_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470__106 clkload1/A VGND VGND VPWR VPWR _1622_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ _1211_/X _1212_/X _1213_/X VGND VGND VPWR VPWR _1214_/X sky130_fd_sc_hd__a21o_1
X_1145_ _1086_/B _1184_/S _1558_/Q VGND VGND VPWR VPWR _1146_/B sky130_fd_sc_hd__o21ba_1
X_1076_ _1076_/A _1086_/B VGND VGND VPWR VPWR _1076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0929_ _1639_/Q _1251_/A _0940_/C VGND VGND VPWR VPWR _0929_/X sky130_fd_sc_hd__and3_1
X_1399__35 clkload3/A VGND VGND VPWR VPWR _1551_/CLK sky130_fd_sc_hd__inv_2
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
X_1373__9 _1533_/CLK VGND VGND VPWR VPWR _1516_/CLK sky130_fd_sc_hd__inv_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1128_ _1234_/B _1235_/A _1127_/X VGND VGND VPWR VPWR _1130_/D sky130_fd_sc_hd__o21ai_4
X_1059_ hold29/X _1592_/Q _1058_/Y VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1476__112 clkload10/A VGND VGND VPWR VPWR _1628_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1453__89 _1454__90/A VGND VGND VPWR VPWR _1605_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1531_ _1531_/CLK _1531_/D VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
X_1600_ _1600_/CLK _1600_/D VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0893_ _0762_/Y _1629_/Q _1640_/Q _0817_/A _0892_/X VGND VGND VPWR VPWR _0896_/C
+ sky130_fd_sc_hd__o221a_1
X_0962_ _1162_/B _1076_/A _1346_/C _1346_/D VGND VGND VPWR VPWR wire17/A sky130_fd_sc_hd__nor4_1
X_1514_ _1514_/CLK _1514_/D VGND VGND VPWR VPWR uo_out[3] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout60 _1331_/C1 VGND VGND VPWR VPWR _1336_/C1 sky130_fd_sc_hd__buf_2
X_1423__59 clkload3/A VGND VGND VPWR VPWR _1575_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1161_ _1080_/A _1147_/Y _1157_/X _1178_/S _1160_/X VGND VGND VPWR VPWR _1161_/X
+ sky130_fd_sc_hd__o311a_1
X_1230_ _1066_/X _1187_/A _1189_/B _1234_/A _1188_/A VGND VGND VPWR VPWR _1230_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1092_ _1580_/Q _1104_/B VGND VGND VPWR VPWR _1092_/X sky130_fd_sc_hd__or2_1
X_0876_ _1608_/Q _1628_/Q VGND VGND VPWR VPWR _0876_/Y sky130_fd_sc_hd__nand2_1
X_0945_ _0963_/A _0945_/B VGND VGND VPWR VPWR _0945_/Y sky130_fd_sc_hd__nor2_2
X_1359_ _1358_/A _1358_/B uo_out[0] VGND VGND VPWR VPWR _1359_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clkload2/A VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_4
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1213_ _1578_/Q _1139_/A _0770_/Y _1577_/Q VGND VGND VPWR VPWR _1213_/X sky130_fd_sc_hd__a22o_1
X_1144_ hold33/X _1146_/A VGND VGND VPWR VPWR _1559_/D sky130_fd_sc_hd__xor2_1
X_1075_ _1072_/A _1192_/A _1074_/X _1117_/C1 VGND VGND VPWR VPWR _1588_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_7_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0928_ _0926_/X _0927_/X _0855_/A VGND VGND VPWR VPWR _1640_/D sky130_fd_sc_hd__o21a_1
X_0859_ _0956_/A _0859_/B VGND VGND VPWR VPWR _1652_/D sky130_fd_sc_hd__and2_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
X_1493__129 clkload8/A VGND VGND VPWR VPWR _1645_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1127_ hold38/A _1548_/Q _1547_/Q VGND VGND VPWR VPWR _1127_/X sky130_fd_sc_hd__or3_2
X_1459__95 clkload9/A VGND VGND VPWR VPWR _1611_/CLK sky130_fd_sc_hd__inv_2
X_1058_ hold29/A _1592_/Q _1060_/B VGND VGND VPWR VPWR _1058_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ _1676_/A VGND VGND VPWR VPWR uio_out[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1499__135 clkload8/A VGND VGND VPWR VPWR _1651_/CLK sky130_fd_sc_hd__inv_2
X_1530_ _1530_/CLK _1530_/D VGND VGND VPWR VPWR _1530_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1429__65 clkload2/A VGND VGND VPWR VPWR _1581_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1659_ _1659_/CLK _1659_/D VGND VGND VPWR VPWR _1659_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0961_ _1159_/B _1072_/A VGND VGND VPWR VPWR _1346_/D sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0892_ _0760_/Y _1634_/Q _0775_/Y hold48/A VGND VGND VPWR VPWR _0892_/X sky130_fd_sc_hd__o22a_1
X_1513_ _1513_/CLK _1513_/D VGND VGND VPWR VPWR uo_out[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout61 _1331_/C1 VGND VGND VPWR VPWR _1351_/A sky130_fd_sc_hd__buf_2
Xfanout50 hold2/A VGND VGND VPWR VPWR _1188_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1160_ _1201_/B _1149_/A _1349_/B uo_out[7] VGND VGND VPWR VPWR _1160_/X sky130_fd_sc_hd__a31o_1
X_1091_ _1159_/B _1089_/X _1090_/X _0845_/A VGND VGND VPWR VPWR _1581_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0944_ _0944_/A _1107_/B VGND VGND VPWR VPWR _0945_/B sky130_fd_sc_hd__nor2_4
X_0875_ _0802_/A _1633_/Q _1634_/Q _0760_/Y _0874_/X VGND VGND VPWR VPWR _0875_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1358_ _1358_/A _1358_/B VGND VGND VPWR VPWR _1358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1289_ hold39/A hold41/A _1334_/S VGND VGND VPWR VPWR _1289_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload3 clkload3/A VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_21_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1212_ _1577_/Q _0770_/Y _0771_/Y _1576_/Q VGND VGND VPWR VPWR _1212_/X sky130_fd_sc_hd__o22a_1
X_1143_ _1143_/A _1143_/B VGND VGND VPWR VPWR _1560_/D sky130_fd_sc_hd__nor2_1
X_1074_ _1162_/B _1086_/B VGND VGND VPWR VPWR _1074_/X sky130_fd_sc_hd__or2_1
X_0927_ _1162_/B _0941_/B VGND VGND VPWR VPWR _0927_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0789_ hold29/A _1592_/Q _1593_/Q _1594_/Q _1623_/Q _1624_/Q VGND VGND VPWR VPWR
+ _0789_/X sky130_fd_sc_hd__mux4_1
X_0858_ _0955_/A1 _1652_/Q _0857_/Y wire19/X _1159_/B VGND VGND VPWR VPWR _0859_/B
+ sky130_fd_sc_hd__a32o_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ _1234_/B _1235_/A VGND VGND VPWR VPWR _1126_/Y sky130_fd_sc_hd__nor2_1
X_1057_ _1057_/A _1060_/B _1057_/C VGND VGND VPWR VPWR _1593_/D sky130_fd_sc_hd__and3_1
XFILLER_0_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1501__137 clkload2/A VGND VGND VPWR VPWR _1653_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_34_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_1675_ _1675_/A VGND VGND VPWR VPWR uio_out[6] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _1159_/B _1107_/X _1108_/X _1117_/C1 VGND VGND VPWR VPWR _1573_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1374__10 _1533_/CLK VGND VGND VPWR VPWR _1517_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1658_ _1658_/CLK _1658_/D VGND VGND VPWR VPWR _1658_/Q sky130_fd_sc_hd__dfxtp_1
X_1589_ _1589_/CLK _1589_/D VGND VGND VPWR VPWR _1589_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1466__102 clkload7/A VGND VGND VPWR VPWR _1618_/CLK sky130_fd_sc_hd__inv_2
X_1507__143 clkload2/A VGND VGND VPWR VPWR _1659_/CLK sky130_fd_sc_hd__inv_2
X_0960_ _0960_/A _0960_/B VGND VGND VPWR VPWR _1627_/D sky130_fd_sc_hd__nand2_1
X_1512_ _1512_/CLK _1512_/D VGND VGND VPWR VPWR uo_out[1] sky130_fd_sc_hd__dfxtp_4
X_0891_ _0817_/A _1640_/Q _0889_/X _0890_/Y hold36/A VGND VGND VPWR VPWR _0891_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout62 fanout63/X VGND VGND VPWR VPWR _1331_/C1 sky130_fd_sc_hd__clkbuf_2
Xfanout51 fanout63/X VGND VGND VPWR VPWR _0855_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 _1586_/Q VGND VGND VPWR VPWR _1162_/C sky130_fd_sc_hd__buf_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ _1581_/Q _1104_/B VGND VGND VPWR VPWR _1090_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0874_ _1611_/Q hold6/A VGND VGND VPWR VPWR _0874_/X sky130_fd_sc_hd__xor2_1
Xclkload10 clkload10/A VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_4
XFILLER_0_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0943_ hold55/A _1550_/Q VGND VGND VPWR VPWR _1107_/B sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1357_ _1157_/X _1355_/Y _1356_/X _1351_/A VGND VGND VPWR VPWR _1512_/D sky130_fd_sc_hd__o211a_1
X_1288_ hold39/A _1342_/A2 _1342_/C1 _1287_/X VGND VGND VPWR VPWR _1288_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload4 clkload4/A VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_4
XFILLER_0_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1211_ _1576_/Q _0771_/Y _1208_/Y _1210_/Y _1209_/X VGND VGND VPWR VPWR _1211_/X
+ sky130_fd_sc_hd__a221o_1
X_1142_ hold58/X _1146_/A hold19/X VGND VGND VPWR VPWR _1143_/B sky130_fd_sc_hd__a21oi_1
X_1073_ _1159_/B _1192_/A _1072_/X _1117_/C1 VGND VGND VPWR VPWR _1589_/D sky130_fd_sc_hd__o211a_1
X_0926_ _0940_/A _1640_/Q _0940_/C VGND VGND VPWR VPWR _0926_/X sky130_fd_sc_hd__and3_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0857_ _0963_/A wire19/X VGND VGND VPWR VPWR _0857_/Y sky130_fd_sc_hd__nor2_2
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ _1625_/Q _0785_/X _1626_/Q VGND VGND VPWR VPWR _0788_/Y sky130_fd_sc_hd__a21boi_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ _1546_/Q hold54/A VGND VGND VPWR VPWR _1235_/A sky130_fd_sc_hd__or2_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ hold29/A _1592_/Q _1593_/Q VGND VGND VPWR VPWR _1057_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0909_ _1260_/A _1530_/Q _0908_/X _0963_/A VGND VGND VPWR VPWR _0910_/C sky130_fd_sc_hd__o31ai_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1674_ hold8/A VGND VGND VPWR VPWR uio_out[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ hold47/X _1122_/B VGND VGND VPWR VPWR _1108_/X sky130_fd_sc_hd__or2_1
X_1039_ _1028_/B _1051_/B _1039_/C VGND VGND VPWR VPWR _1602_/D sky130_fd_sc_hd__and3b_1
X_1483__119 clkload1/A VGND VGND VPWR VPWR _1635_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1657_ _1657_/CLK _1657_/D VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfxtp_1
X_1588_ _1588_/CLK _1588_/D VGND VGND VPWR VPWR _1588_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0890_ _1616_/Q _1636_/Q VGND VGND VPWR VPWR _0890_/Y sky130_fd_sc_hd__nand2_1
X_1434__70 clkload5/A VGND VGND VPWR VPWR _1586_/CLK sky130_fd_sc_hd__inv_2
X_1511_ _1511_/CLK _1511_/D VGND VGND VPWR VPWR uo_out[0] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_10_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1489__125 clkload2/A VGND VGND VPWR VPWR _1641_/CLK sky130_fd_sc_hd__inv_2
Xfanout63 input1/X VGND VGND VPWR VPWR fanout63/X sky130_fd_sc_hd__clkbuf_2
Xfanout41 _1348_/D VGND VGND VPWR VPWR _1260_/A sky130_fd_sc_hd__buf_2
Xfanout52 fanout63/X VGND VGND VPWR VPWR _0845_/A sky130_fd_sc_hd__clkbuf_2
Xfanout30 _1643_/Q VGND VGND VPWR VPWR _0923_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload11 _1372__8/A VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_16
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ _0940_/X _0941_/X _0855_/A VGND VGND VPWR VPWR _1635_/D sky130_fd_sc_hd__o21a_1
X_0873_ hold48/A _0775_/Y _0776_/Y _1621_/Q VGND VGND VPWR VPWR _0873_/X sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1356_ _1355_/A _1358_/B uo_out[1] VGND VGND VPWR VPWR _1356_/X sky130_fd_sc_hd__a21o_1
X_1287_ hold41/A _1337_/B VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__or2_1
Xclkload5 clkload5/A VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_21_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1404__40 clkload6/A VGND VGND VPWR VPWR _1556_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1072_ _1072_/A _1086_/B VGND VGND VPWR VPWR _1072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1141_ _1141_/A _1141_/B VGND VGND VPWR VPWR _1561_/D sky130_fd_sc_hd__nor2_1
X_1210_ hold35/A _1558_/Q VGND VGND VPWR VPWR _1210_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0787_ _1625_/Q _0787_/B VGND VGND VPWR VPWR _0787_/Y sky130_fd_sc_hd__nand2b_1
X_0925_ _0923_/X _0924_/X _0845_/A VGND VGND VPWR VPWR _1641_/D sky130_fd_sc_hd__o21a_1
X_0856_ _1107_/A hold55/A _1550_/Q VGND VGND VPWR VPWR wire19/A sky130_fd_sc_hd__nor3b_1
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1339_ _1518_/Q _1516_/Q _1339_/S VGND VGND VPWR VPWR _1339_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1124_ hold42/A _1188_/A VGND VGND VPWR VPWR _1234_/B sky130_fd_sc_hd__and2b_1
X_1055_ _1023_/D _1060_/B _1055_/C VGND VGND VPWR VPWR _1594_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1395__31 clkload4/A VGND VGND VPWR VPWR _1547_/CLK sky130_fd_sc_hd__inv_2
X_0839_ _0923_/A _1659_/Q _0836_/Y _0836_/A _1148_/B VGND VGND VPWR VPWR _0840_/B
+ sky130_fd_sc_hd__a32o_1
X_0908_ _1162_/A _1346_/C _1148_/B _1162_/B VGND VGND VPWR VPWR _0908_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1673_ hold11/A VGND VGND VPWR VPWR uio_out[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1038_ hold31/A hold5/A _1045_/A _1602_/Q VGND VGND VPWR VPWR _1039_/C sky130_fd_sc_hd__a31o_1
X_1107_ _1107_/A _1107_/B VGND VGND VPWR VPWR _1107_/X sky130_fd_sc_hd__or2_2
XFILLER_0_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1656_ _1656_/CLK _1656_/D VGND VGND VPWR VPWR _1656_/Q sky130_fd_sc_hd__dfxtp_1
X_1587_ _1587_/CLK _1587_/D VGND VGND VPWR VPWR _1587_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1510_ _1510_/CLK _1510_/D VGND VGND VPWR VPWR _1675_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1639_ _1639_/CLK _1639_/D VGND VGND VPWR VPWR _1639_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout20 _1084_/B VGND VGND VPWR VPWR _1192_/A sky130_fd_sc_hd__clkbuf_4
Xfanout42 _1585_/Q VGND VGND VPWR VPWR _1348_/D sky130_fd_sc_hd__clkbuf_4
Xfanout53 fanout63/X VGND VGND VPWR VPWR _0971_/A sky130_fd_sc_hd__clkbuf_2
Xfanout31 _1643_/Q VGND VGND VPWR VPWR _0955_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ _0941_/A _0941_/B VGND VGND VPWR VPWR _0941_/X sky130_fd_sc_hd__and2_1
XFILLER_0_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload12 _1533_/CLK VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_12
X_0872_ _0956_/A _0872_/B VGND VGND VPWR VPWR _1645_/D sky130_fd_sc_hd__and2_1
X_1355_ _1355_/A _1358_/B VGND VGND VPWR VPWR _1355_/Y sky130_fd_sc_hd__nand2_1
X_1286_ hold39/X _1345_/A2 _1285_/X _1336_/C1 VGND VGND VPWR VPWR _1528_/D sky130_fd_sc_hd__o211a_1
Xclkload6 clkload6/A VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_21_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ _1187_/A _1234_/A _1066_/X VGND VGND VPWR VPWR _1084_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ hold18/X _1143_/A VGND VGND VPWR VPWR _1141_/B sky130_fd_sc_hd__nor2_1
X_0924_ _1072_/A _0941_/B VGND VGND VPWR VPWR _0924_/X sky130_fd_sc_hd__and2_1
X_0786_ hold14/A hold31/A hold5/A _1602_/Q _1623_/Q _1624_/Q VGND VGND VPWR VPWR _0787_/B
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0855_ _0855_/A _0855_/B VGND VGND VPWR VPWR _1653_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1338_ _1518_/Q _1342_/A2 _1342_/C1 _1337_/X VGND VGND VPWR VPWR _1338_/X sky130_fd_sc_hd__o211a_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ _1260_/A _1176_/A _1530_/Q VGND VGND VPWR VPWR _1270_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1123_ _1349_/B _1107_/X _1122_/X _1199_/A VGND VGND VPWR VPWR _1566_/D sky130_fd_sc_hd__o211a_1
X_1054_ hold29/A _1592_/Q _1593_/Q _1594_/Q VGND VGND VPWR VPWR _1055_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0907_ _1260_/A _1346_/C _1339_/S _0903_/X VGND VGND VPWR VPWR _0910_/B sky130_fd_sc_hd__or4b_1
X_0838_ _0855_/A _0838_/B VGND VGND VPWR VPWR _1660_/D sky130_fd_sc_hd__and2_1
X_0769_ hold34/X VGND VGND VPWR VPWR _1139_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1672_ _1672_/A VGND VGND VPWR VPWR uio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1106_ _1107_/A _1107_/B VGND VGND VPWR VPWR _1122_/B sky130_fd_sc_hd__nor2_1
X_1037_ _1037_/A _1037_/B VGND VGND VPWR VPWR _1603_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1455__91 clkload9/A VGND VGND VPWR VPWR _1607_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380__16 clkload13/A VGND VGND VPWR VPWR _1523_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1655_ _1655_/CLK _1655_/D VGND VGND VPWR VPWR _1655_/Q sky130_fd_sc_hd__dfxtp_1
X_1586_ _1586_/CLK _1586_/D VGND VGND VPWR VPWR _1586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1473__109 _1454__90/A VGND VGND VPWR VPWR _1625_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1425__61 clkload0/A VGND VGND VPWR VPWR _1577_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1638_ _1638_/CLK _1638_/D VGND VGND VPWR VPWR _1638_/Q sky130_fd_sc_hd__dfxtp_1
X_1569_ _1569_/CLK _1569_/D VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfxtp_1
Xfanout21 _1339_/S VGND VGND VPWR VPWR _1334_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout54 _1259_/C1 VGND VGND VPWR VPWR _1199_/A sky130_fd_sc_hd__clkbuf_4
Xfanout43 _1176_/A VGND VGND VPWR VPWR _1201_/B sky130_fd_sc_hd__clkbuf_4
Xfanout32 _1643_/Q VGND VGND VPWR VPWR _0959_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0940_ _0940_/A _1635_/Q _0940_/C VGND VGND VPWR VPWR _0940_/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload13 clkload13/A VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0871_ _0955_/A1 _1645_/Q _0857_/Y wire19/X _1264_/B VGND VGND VPWR VPWR _0872_/B
+ sky130_fd_sc_hd__a32o_1
X_1354_ _1157_/X _1352_/Y _1353_/X _1351_/A VGND VGND VPWR VPWR _1513_/D sky130_fd_sc_hd__o211a_1
X_1285_ _1340_/A1 _1284_/X _1283_/X _1344_/C1 VGND VGND VPWR VPWR _1285_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload7 clkload7/A VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_16
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1495__131 clkload10/A VGND VGND VPWR VPWR _1647_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1070_ _1187_/A _1234_/A _1066_/X VGND VGND VPWR VPWR _1086_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0854_ _0923_/A _1653_/Q _0836_/Y _0836_/A _0941_/A VGND VGND VPWR VPWR _0855_/B
+ sky130_fd_sc_hd__a32o_1
X_0923_ _0923_/A _1641_/Q _0940_/C VGND VGND VPWR VPWR _0923_/X sky130_fd_sc_hd__and3_1
X_1479__115 clkload10/A VGND VGND VPWR VPWR _1631_/CLK sky130_fd_sc_hd__inv_2
X_0785_ hold25/A hold4/A _1605_/Q hold1/A _1623_/Q _1624_/Q VGND VGND VPWR VPWR _0785_/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1337_ _1516_/Q _1337_/B VGND VGND VPWR VPWR _1337_/X sky130_fd_sc_hd__or2_1
X_1268_ _1516_/Q _1348_/C _1260_/Y _1267_/X _1342_/C1 VGND VGND VPWR VPWR _1268_/X
+ sky130_fd_sc_hd__a221o_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1199_ _1199_/A _1199_/B VGND VGND VPWR VPWR _1199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1122_ hold45/X _1122_/B VGND VGND VPWR VPWR _1122_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1053_ hold15/X _1023_/D _1052_/Y VGND VGND VPWR VPWR _1595_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0906_ _1162_/A _1072_/A _0906_/C VGND VGND VPWR VPWR _0906_/X sky130_fd_sc_hd__or3_1
X_0837_ _0923_/A _1660_/Q _0836_/Y _0836_/A _1159_/B VGND VGND VPWR VPWR _0838_/B
+ sky130_fd_sc_hd__a32o_1
X_0768_ hold21/A VGND VGND VPWR VPWR _0768_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1386__22 clkload13/A VGND VGND VPWR VPWR _1529_/CLK sky130_fd_sc_hd__inv_2
X_1671_ hold17/A VGND VGND VPWR VPWR uio_oe[7] sky130_fd_sc_hd__buf_2
XFILLER_0_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ _0941_/A _1089_/X _1104_/X _0971_/A VGND VGND VPWR VPWR _1574_/D sky130_fd_sc_hd__o211a_1
X_1036_ hold25/X _1028_/B _1051_/B VGND VGND VPWR VPWR _1037_/B sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1654_ _1654_/CLK _1654_/D VGND VGND VPWR VPWR _1654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1585_ _1585_/CLK _1585_/D VGND VGND VPWR VPWR _1585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _1016_/B _1019_/B _1019_/C VGND VGND VPWR VPWR _1607_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1637_ _1637_/CLK _1637_/D VGND VGND VPWR VPWR _1637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1440__76 clkload1/A VGND VGND VPWR VPWR _1592_/CLK sky130_fd_sc_hd__inv_2
X_1568_ _1568_/CLK _1568_/D VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__dfxtp_1
Xfanout55 _1259_/C1 VGND VGND VPWR VPWR _1117_/C1 sky130_fd_sc_hd__buf_2
Xfanout22 _0906_/X VGND VGND VPWR VPWR _1339_/S sky130_fd_sc_hd__buf_2
Xfanout33 _1159_/B VGND VGND VPWR VPWR _1162_/A sky130_fd_sc_hd__buf_2
Xfanout11 _0984_/Y VGND VGND VPWR VPWR _1009_/C sky130_fd_sc_hd__clkbuf_2
Xfanout44 _1584_/Q VGND VGND VPWR VPWR _1176_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0870_ _0960_/A _0870_/B VGND VGND VPWR VPWR _1646_/D sky130_fd_sc_hd__nand2_1
Xclkload14 _1541_/CLK VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__inv_16
X_1353_ _1352_/A _1358_/B uo_out[2] VGND VGND VPWR VPWR _1353_/X sky130_fd_sc_hd__a21o_1
X_1284_ hold32/A hold44/A _1334_/S VGND VGND VPWR VPWR _1284_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ _1611_/Q _1010_/B VGND VGND VPWR VPWR _1008_/B sky130_fd_sc_hd__and2_1
Xclkload8 clkload8/A VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_8
XFILLER_0_1_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0922_ _0920_/X _0921_/X _0855_/A VGND VGND VPWR VPWR _1642_/D sky130_fd_sc_hd__o21a_1
X_0853_ _0855_/A _0853_/B VGND VGND VPWR VPWR _1654_/D sky130_fd_sc_hd__and2_1
X_1410__46 clkload0/A VGND VGND VPWR VPWR _1562_/CLK sky130_fd_sc_hd__inv_2
X_0784_ hold55/A _1550_/Q _1107_/A VGND VGND VPWR VPWR _0836_/A sky130_fd_sc_hd__nor3_4
XFILLER_0_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 rst_n VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
X_1267_ _1334_/S _1267_/B _1267_/C VGND VGND VPWR VPWR _1267_/X sky130_fd_sc_hd__and3_1
X_1198_ _1548_/Q _1199_/B _1197_/Y VGND VGND VPWR VPWR _1548_/D sky130_fd_sc_hd__a21o_1
X_1336_ _1518_/Q _1345_/A2 _1335_/X _1336_/C1 VGND VGND VPWR VPWR _1518_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ _1149_/A _1107_/X _1120_/X _1199_/A VGND VGND VPWR VPWR _1567_/D sky130_fd_sc_hd__o211a_1
X_1052_ hold15/A _1023_/D _1060_/B VGND VGND VPWR VPWR _1052_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0905_ _1162_/A _1148_/B _0906_/C VGND VGND VPWR VPWR _1348_/C sky130_fd_sc_hd__nor3_1
XFILLER_0_3_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0767_ hold27/X VGND VGND VPWR VPWR _1136_/A sky130_fd_sc_hd__inv_2
X_0836_ _0836_/A _0963_/A VGND VGND VPWR VPWR _0836_/Y sky130_fd_sc_hd__nor2_2
X_1319_ _1522_/Q _1520_/Q _1334_/S VGND VGND VPWR VPWR _1319_/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1670_ hold17/A VGND VGND VPWR VPWR uio_oe[6] sky130_fd_sc_hd__buf_2
X_1035_ hold4/X _1037_/A _1034_/Y VGND VGND VPWR VPWR _1604_/D sky130_fd_sc_hd__a21oi_1
X_1104_ hold35/X _1104_/B VGND VGND VPWR VPWR _1104_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ _0835_/A _0831_/C _0834_/D _0831_/D VGND VGND VPWR VPWR _0822_/B sky130_fd_sc_hd__or4_1
X_1446__82 _1454__90/A VGND VGND VPWR VPWR _1598_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1653_ _1653_/CLK _1653_/D VGND VGND VPWR VPWR _1653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1584_ _1584_/CLK _1584_/D VGND VGND VPWR VPWR _1584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ _1607_/Q _1030_/A VGND VGND VPWR VPWR _1019_/B sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_14_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1567_ _1567_/CLK _1567_/D VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__dfxtp_1
X_1636_ _1636_/CLK _1636_/D VGND VGND VPWR VPWR _1636_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout56 _1259_/C1 VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__clkbuf_2
X_1416__52 clkload6/A VGND VGND VPWR VPWR _1568_/CLK sky130_fd_sc_hd__inv_2
Xfanout34 _1589_/Q VGND VGND VPWR VPWR _1159_/B sky130_fd_sc_hd__buf_2
Xfanout12 _0984_/Y VGND VGND VPWR VPWR _1019_/C sky130_fd_sc_hd__buf_1
Xfanout45 _1349_/A VGND VGND VPWR VPWR _1149_/A sky130_fd_sc_hd__clkbuf_4
Xfanout23 _1178_/S VGND VGND VPWR VPWR _1340_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1352_ _1352_/A _1358_/B VGND VGND VPWR VPWR _1352_/Y sky130_fd_sc_hd__nand2_1
X_1283_ hold32/A _1342_/A2 _1333_/B1 _1282_/X VGND VGND VPWR VPWR _1283_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0998_ _1610_/Q _1030_/A _0998_/C VGND VGND VPWR VPWR _1010_/B sky130_fd_sc_hd__and3_1
Xclkload9 clkload9/A VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_6
X_1619_ _1619_/CLK _1619_/D VGND VGND VPWR VPWR _1619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0921_ _1159_/B _0941_/B VGND VGND VPWR VPWR _0921_/X sky130_fd_sc_hd__and2_1
XFILLER_0_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0852_ _0923_/A _1654_/Q _0836_/Y _0836_/A _1149_/A VGND VGND VPWR VPWR _0853_/B
+ sky130_fd_sc_hd__a32o_1
X_0783_ hold12/A _0901_/A hold3/A VGND VGND VPWR VPWR _1107_/A sky130_fd_sc_hd__or3b_4
X_1335_ _1340_/A1 _1334_/X _1333_/X _1344_/C1 VGND VGND VPWR VPWR _1335_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_1_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 ui_in[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1266_ _1536_/Q _1352_/A _1265_/X _1176_/A _1348_/D VGND VGND VPWR VPWR _1267_/C
+ sky130_fd_sc_hd__a2111o_1
X_1197_ _1199_/A _1197_/B VGND VGND VPWR VPWR _1197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1120_ hold56/X _1122_/B VGND VGND VPWR VPWR _1120_/X sky130_fd_sc_hd__or2_1
X_1485__121 clkload1/A VGND VGND VPWR VPWR _1637_/CLK sky130_fd_sc_hd__inv_2
X_1051_ _1022_/X _1051_/B _1051_/C VGND VGND VPWR VPWR _1596_/D sky130_fd_sc_hd__and3b_1
X_0904_ _1346_/A _1076_/A VGND VGND VPWR VPWR _0906_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0835_ _0835_/A _0835_/B _0835_/C _0835_/D VGND VGND VPWR VPWR _1248_/A sky130_fd_sc_hd__or4_1
X_0766_ hold9/A VGND VGND VPWR VPWR _0766_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1318_ _1522_/Q _0913_/Y _1342_/C1 _1317_/X VGND VGND VPWR VPWR _1318_/X sky130_fd_sc_hd__o211a_1
X_1249_ _0984_/B _1248_/X _1676_/A VGND VGND VPWR VPWR _1251_/B sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_19_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1469__105 clkload1/A VGND VGND VPWR VPWR _1621_/CLK sky130_fd_sc_hd__inv_2
X_1377__13 _1541_/CLK VGND VGND VPWR VPWR _1520_/CLK sky130_fd_sc_hd__inv_2
X_1034_ hold4/X _1037_/A _1051_/B VGND VGND VPWR VPWR _1034_/Y sky130_fd_sc_hd__o21ai_1
X_1103_ _1149_/A _1089_/X _1102_/X _0971_/A VGND VGND VPWR VPWR _1575_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_33_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0818_ _0818_/A _0833_/B _0833_/C _0832_/B VGND VGND VPWR VPWR _0825_/B sky130_fd_sc_hd__or4_1
X_1369__5 _1533_/CLK VGND VGND VPWR VPWR _1512_/CLK sky130_fd_sc_hd__inv_2
X_1461__97 clkload9/A VGND VGND VPWR VPWR _1613_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1652_ _1652_/CLK _1652_/D VGND VGND VPWR VPWR _1652_/Q sky130_fd_sc_hd__dfxtp_1
X_1583_ _1583_/CLK _1583_/D VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1017_ _1014_/B _1017_/B _1019_/C VGND VGND VPWR VPWR _1608_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1566_ _1566_/CLK _1566_/D VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
X_1635_ _1635_/CLK _1635_/D VGND VGND VPWR VPWR _1635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout57 fanout63/X VGND VGND VPWR VPWR _1259_/C1 sky130_fd_sc_hd__clkbuf_2
Xfanout24 _1159_/Y VGND VGND VPWR VPWR _1178_/S sky130_fd_sc_hd__clkbuf_4
Xfanout13 _1276_/X VGND VGND VPWR VPWR _1344_/C1 sky130_fd_sc_hd__buf_2
Xfanout46 hold26/A VGND VGND VPWR VPWR _1349_/A sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_24_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout35 _1072_/A VGND VGND VPWR VPWR _1148_/B sky130_fd_sc_hd__buf_2
XFILLER_0_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1431__67 clkload10/A VGND VGND VPWR VPWR _1583_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1351_ _1351_/A _1351_/B VGND VGND VPWR VPWR _1514_/D sky130_fd_sc_hd__and2_1
X_1282_ hold44/A _1337_/B VGND VGND VPWR VPWR _1282_/X sky130_fd_sc_hd__or2_1
X_1618_ _1618_/CLK _1618_/D VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_2
X_0997_ _1030_/A _0998_/C VGND VGND VPWR VPWR _1012_/B sky130_fd_sc_hd__and2_1
X_1549_ _1549_/CLK _1549_/D VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0920_ _0940_/A _1642_/Q _0940_/C VGND VGND VPWR VPWR _0920_/X sky130_fd_sc_hd__and3_1
X_0782_ hold38/A _1548_/Q _1547_/Q VGND VGND VPWR VPWR _0901_/A sky130_fd_sc_hd__nand3_1
X_0851_ _0956_/A _0851_/B VGND VGND VPWR VPWR _1655_/D sky130_fd_sc_hd__and2_1
X_1265_ _1534_/Q _1358_/A _1355_/A _1535_/Q _1264_/X VGND VGND VPWR VPWR _1265_/X
+ sky130_fd_sc_hd__a221o_1
X_1334_ _1519_/Q _1517_/Q _1334_/S VGND VGND VPWR VPWR _1334_/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 ui_in[1] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
X_1196_ _1127_/X _1193_/B _1195_/Y _1199_/A VGND VGND VPWR VPWR _1549_/D sky130_fd_sc_hd__o211ai_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1401__37 clkload4/A VGND VGND VPWR VPWR _1553_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1050_ hold15/A _1023_/D _1596_/Q VGND VGND VPWR VPWR _1051_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0834_ _0834_/A _0834_/B _0834_/C _0834_/D VGND VGND VPWR VPWR _0835_/D sky130_fd_sc_hd__or4_1
X_0903_ _1162_/A _1148_/B _1530_/Q _1162_/B VGND VGND VPWR VPWR _0903_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0765_ _1264_/B VGND VGND VPWR VPWR _1084_/A sky130_fd_sc_hd__inv_2
X_1317_ _1520_/Q _1322_/B VGND VGND VPWR VPWR _1317_/X sky130_fd_sc_hd__or2_1
X_1248_ _1248_/A _1248_/B _1248_/C _1248_/D VGND VGND VPWR VPWR _1248_/X sky130_fd_sc_hd__or4_1
X_1179_ uo_out[4] _1178_/X _1179_/S VGND VGND VPWR VPWR _1180_/B sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1392__28 clkload4/A VGND VGND VPWR VPWR _1544_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1102_ hold53/X _1104_/B VGND VGND VPWR VPWR _1102_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1033_ _1029_/X _1051_/B _1033_/C VGND VGND VPWR VPWR _1605_/D sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_16_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0817_ _0817_/A _1658_/Q VGND VGND VPWR VPWR _0832_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_3_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1437__73 clkload5/A VGND VGND VPWR VPWR _1589_/CLK sky130_fd_sc_hd__inv_2
X_1651_ _1651_/CLK _1651_/D VGND VGND VPWR VPWR _1651_/Q sky130_fd_sc_hd__dfxtp_1
X_1582_ _1582_/CLK _1582_/D VGND VGND VPWR VPWR _1582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1016_ _1608_/Q _1016_/B VGND VGND VPWR VPWR _1017_/B sky130_fd_sc_hd__or2_1
X_1371__7 _1533_/CLK VGND VGND VPWR VPWR _1514_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ _1634_/CLK _1634_/D VGND VGND VPWR VPWR _1634_/Q sky130_fd_sc_hd__dfxtp_1
X_1565_ _1565_/CLK hold10/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout47 _0941_/A VGND VGND VPWR VPWR _1349_/B sky130_fd_sc_hd__buf_2
Xfanout14 _1275_/Y VGND VGND VPWR VPWR _1345_/A2 sky130_fd_sc_hd__buf_2
Xfanout25 _1342_/C1 VGND VGND VPWR VPWR _1333_/B1 sky130_fd_sc_hd__buf_2
Xfanout58 _1331_/C1 VGND VGND VPWR VPWR _0956_/A sky130_fd_sc_hd__clkbuf_2
Xfanout36 _1588_/Q VGND VGND VPWR VPWR _1072_/A sky130_fd_sc_hd__buf_2
X_1407__43 clkload3/A VGND VGND VPWR VPWR _1559_/CLK sky130_fd_sc_hd__inv_2
X_1350_ uo_out[3] _1157_/X _1350_/S VGND VGND VPWR VPWR _1351_/B sky130_fd_sc_hd__mux2_1
X_1281_ hold32/X _1345_/A2 _1280_/X _1336_/C1 VGND VGND VPWR VPWR _1529_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_25_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0996_ _1608_/Q _1607_/Q _1030_/A VGND VGND VPWR VPWR _1014_/B sky130_fd_sc_hd__and3_1
X_1617_ _1617_/CLK _1617_/D VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
X_1548_ _1548_/CLK _1548_/D VGND VGND VPWR VPWR _1548_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0850_ _0955_/A1 _1655_/Q _0836_/Y _0836_/A _1176_/A VGND VGND VPWR VPWR _0851_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 ui_in[2] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
X_1264_ _1349_/A _1264_/B _1537_/Q VGND VGND VPWR VPWR _1264_/X sky130_fd_sc_hd__and3_1
X_1333_ _1519_/Q _1342_/A2 _1333_/B1 _1332_/X VGND VGND VPWR VPWR _1333_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1195_ hold38/X _1197_/B VGND VGND VPWR VPWR _1195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0979_ hold48/X _0981_/D VGND VGND VPWR VPWR _0979_/Y sky130_fd_sc_hd__nand2_1
X_1398__34 clkload4/A VGND VGND VPWR VPWR _1550_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0833_ _0833_/A _0833_/B _0833_/C _0833_/D VGND VGND VPWR VPWR _0835_/C sky130_fd_sc_hd__or4_1
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0902_ _0944_/A hold55/A _1550_/Q VGND VGND VPWR VPWR _1346_/C sky130_fd_sc_hd__or3b_2
X_0764_ _1349_/A VGND VGND VPWR VPWR _1082_/A sky130_fd_sc_hd__inv_2
X_1178_ _0941_/A _1177_/X _1178_/S VGND VGND VPWR VPWR _1178_/X sky130_fd_sc_hd__mux2_1
X_1316_ _1522_/Q _1275_/Y _1315_/X _1336_/C1 VGND VGND VPWR VPWR _1522_/D sky130_fd_sc_hd__o211a_1
X_1247_ _1653_/Q _1658_/Q _1659_/Q _1660_/Q VGND VGND VPWR VPWR _1248_/D sky130_fd_sc_hd__or4_1
XFILLER_0_34_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1032_ hold25/A hold4/A _1028_/B _1605_/Q VGND VGND VPWR VPWR _1033_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1101_ _1201_/B _1089_/X _1100_/X _0971_/A VGND VGND VPWR VPWR _1576_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0816_ _1607_/Q _0777_/Y _1652_/Q _0760_/Y VGND VGND VPWR VPWR _0833_/C sky130_fd_sc_hd__o22ai_1
X_1475__111 clkload10/A VGND VGND VPWR VPWR _1627_/CLK sky130_fd_sc_hd__inv_2
X_1452__88 _1454__90/A VGND VGND VPWR VPWR _1604_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ _1650_/CLK _1650_/D VGND VGND VPWR VPWR _1650_/Q sky130_fd_sc_hd__dfxtp_1
X_1581_ _1581_/CLK _1581_/D VGND VGND VPWR VPWR _1581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ _1012_/B _1015_/B _1019_/C VGND VGND VPWR VPWR _1609_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_8_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1564_ _1564_/CLK _1564_/D VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfxtp_1
X_1633_ _1633_/CLK _1633_/D VGND VGND VPWR VPWR _1633_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_18_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout26 _1158_/X VGND VGND VPWR VPWR _1342_/C1 sky130_fd_sc_hd__clkbuf_2
Xfanout15 _1060_/B VGND VGND VPWR VPWR _1051_/B sky130_fd_sc_hd__clkbuf_2
Xfanout37 _1346_/A VGND VGND VPWR VPWR _1162_/B sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout48 _1264_/B VGND VGND VPWR VPWR _0941_/A sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_32_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout59 _1331_/C1 VGND VGND VPWR VPWR _0960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1422__58 clkload3/A VGND VGND VPWR VPWR _1574_/CLK sky130_fd_sc_hd__inv_2
X_1280_ _1340_/A1 _1279_/X _1278_/X _1344_/C1 VGND VGND VPWR VPWR _1280_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ _1607_/Q _1030_/A VGND VGND VPWR VPWR _1016_/B sky130_fd_sc_hd__and2_1
X_1547_ _1547_/CLK _1547_/D VGND VGND VPWR VPWR _1547_/Q sky130_fd_sc_hd__dfxtp_2
X_1616_ _1616_/CLK _1616_/D VGND VGND VPWR VPWR _1616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0780_ _1653_/Q VGND VGND VPWR VPWR _0780_/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 ui_in[3] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
X_1263_ _1539_/Q _1355_/A _1261_/X _1262_/X VGND VGND VPWR VPWR _1267_/B sky130_fd_sc_hd__a211o_1
X_1194_ _1548_/Q _1199_/B VGND VGND VPWR VPWR _1197_/B sky130_fd_sc_hd__or2_1
X_1332_ _1517_/Q _1337_/B VGND VGND VPWR VPWR _1332_/X sky130_fd_sc_hd__or2_1
X_0978_ _0981_/D VGND VGND VPWR VPWR _0978_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0763_ _1176_/A VGND VGND VPWR VPWR _1080_/A sky130_fd_sc_hd__inv_2
X_1492__128 clkload1/A VGND VGND VPWR VPWR _1644_/CLK sky130_fd_sc_hd__inv_2
X_0832_ _0832_/A _0832_/B _0832_/C _0832_/D VGND VGND VPWR VPWR _0833_/D sky130_fd_sc_hd__or4_1
X_0901_ _0901_/A hold3/A hold12/A VGND VGND VPWR VPWR _0944_/A sky130_fd_sc_hd__or3b_4
X_1315_ _1340_/A1 _1314_/X _1313_/X _1344_/C1 VGND VGND VPWR VPWR _1315_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1177_ _1157_/X uo_out[4] _1177_/S VGND VGND VPWR VPWR _1177_/X sky130_fd_sc_hd__mux2_1
X_1246_ _1650_/Q _1651_/Q _1652_/Q _1246_/D VGND VGND VPWR VPWR _1248_/C sky130_fd_sc_hd__or4_1
X_1458__94 clkload9/A VGND VGND VPWR VPWR _1610_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_9_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload8/A sky130_fd_sc_hd__clkbuf_8
X_1031_ hold1/X _1029_/X _1051_/B VGND VGND VPWR VPWR _1606_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1100_ _1576_/Q _1104_/B VGND VGND VPWR VPWR _1100_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0815_ _1615_/Q _0780_/Y _1658_/Q _0817_/A _0814_/X VGND VGND VPWR VPWR _0833_/B
+ sky130_fd_sc_hd__a221o_1
X_1383__19 clkload13/A VGND VGND VPWR VPWR _1526_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1229_ _1546_/Q _1130_/D _1228_/X _1259_/C1 VGND VGND VPWR VPWR _1546_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_15_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1580_ _1580_/CLK _1580_/D VGND VGND VPWR VPWR _1580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _1609_/Q _1014_/B VGND VGND VPWR VPWR _1015_/B sky130_fd_sc_hd__or2_1
X_1428__64 clkload0/A VGND VGND VPWR VPWR _1580_/CLK sky130_fd_sc_hd__inv_2
X_1498__134 clkload10/A VGND VGND VPWR VPWR _1650_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1632_ _1632_/CLK _1632_/D VGND VGND VPWR VPWR _1632_/Q sky130_fd_sc_hd__dfxtp_1
X_1563_ _1563_/CLK _1563_/D VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
Xfanout49 _1582_/Q VGND VGND VPWR VPWR _1264_/B sky130_fd_sc_hd__buf_2
XFILLER_0_29_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout27 _0913_/Y VGND VGND VPWR VPWR _1342_/A2 sky130_fd_sc_hd__buf_2
Xfanout16 _1030_/Y VGND VGND VPWR VPWR _1060_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout38 _1587_/Q VGND VGND VPWR VPWR _1346_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ _0976_/Y _1009_/C _0994_/C VGND VGND VPWR VPWR _1616_/D sky130_fd_sc_hd__and3b_1
X_1546_ _1546_/CLK _1546_/D VGND VGND VPWR VPWR _1546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1615_ _1615_/CLK _1615_/D VGND VGND VPWR VPWR _1615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1331_ _1519_/Q _1345_/A2 _1330_/X _1331_/C1 VGND VGND VPWR VPWR _1519_/D sky130_fd_sc_hd__o211a_1
Xinput6 ui_in[4] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
X_1193_ _1547_/Q _1193_/B VGND VGND VPWR VPWR _1199_/B sky130_fd_sc_hd__or2_1
XFILLER_0_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1262_ _1538_/Q _1358_/A _1352_/A _1540_/Q VGND VGND VPWR VPWR _1262_/X sky130_fd_sc_hd__a22o_1
X_0977_ hold37/A _1616_/Q _1030_/A _0977_/D VGND VGND VPWR VPWR _0981_/D sky130_fd_sc_hd__and4_2
XFILLER_0_14_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1529_ _1529_/CLK _1529_/D VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1389__25 clkload2/A VGND VGND VPWR VPWR _1532_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ hold36/X _0984_/B _0899_/Y VGND VGND VPWR VPWR _1644_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_22_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ _0831_/A _0831_/B _0831_/C _0831_/D VGND VGND VPWR VPWR _0832_/D sky130_fd_sc_hd__or4_1
X_0762_ _1609_/Q VGND VGND VPWR VPWR _0762_/Y sky130_fd_sc_hd__inv_2
X_1314_ hold46/A _1521_/Q _1334_/S VGND VGND VPWR VPWR _1314_/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1176_ _1176_/A _1358_/A VGND VGND VPWR VPWR _1177_/S sky130_fd_sc_hd__nand2_1
X_1245_ _1654_/Q _1655_/Q _1656_/Q hold20/A VGND VGND VPWR VPWR _1246_/D sky130_fd_sc_hd__or4_1
XFILLER_0_34_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ _1030_/A _1030_/B VGND VGND VPWR VPWR _1030_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ _1621_/Q _1659_/Q VGND VGND VPWR VPWR _0814_/X sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_16_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1500__136 clkload8/A VGND VGND VPWR VPWR _1652_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1228_ _1355_/A _1203_/B _1221_/X _1227_/X VGND VGND VPWR VPWR _1228_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1159_ _1072_/A _1159_/B VGND VGND VPWR VPWR _1159_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1013_ _1010_/B _1013_/B _1019_/C VGND VGND VPWR VPWR _1610_/D sky130_fd_sc_hd__and3b_1
X_1443__79 _1454__90/A VGND VGND VPWR VPWR _1595_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload7/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1631_ _1631_/CLK _1631_/D VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
X_1562_ _1562_/CLK _1562_/D VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
X_1465__101 clkload7/A VGND VGND VPWR VPWR _1617_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 _1586_/Q VGND VGND VPWR VPWR _1076_/A sky130_fd_sc_hd__buf_2
X_1506__142 clkload8/A VGND VGND VPWR VPWR _1658_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_17_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 _1322_/B VGND VGND VPWR VPWR _1337_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ _0993_/A _0993_/B VGND VGND VPWR VPWR _0994_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_25_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1614_ _1614_/CLK _1614_/D VGND VGND VPWR VPWR _1614_/Q sky130_fd_sc_hd__dfxtp_1
X_1413__49 clkload0/A VGND VGND VPWR VPWR _1565_/CLK sky130_fd_sc_hd__inv_2
X_1545_ _1545_/CLK _1545_/D VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1261_ _1349_/A _1264_/B _1541_/Q _1080_/A _1348_/D VGND VGND VPWR VPWR _1261_/X
+ sky130_fd_sc_hd__a311o_1
X_1330_ _1340_/A1 _1329_/X _1328_/X _1344_/C1 VGND VGND VPWR VPWR _1330_/X sky130_fd_sc_hd__a211o_1
Xinput7 ui_in[5] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
X_1192_ _1192_/A _1258_/A VGND VGND VPWR VPWR _1193_/B sky130_fd_sc_hd__nor2_1
X_0976_ _0993_/A _0993_/B VGND VGND VPWR VPWR _0976_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1528_ _1528_/CLK _1528_/D VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
X_0830_ _0830_/A _0830_/B _0830_/C _0830_/D VGND VGND VPWR VPWR _0835_/B sky130_fd_sc_hd__or4_1
XFILLER_0_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0761_ _1613_/Q VGND VGND VPWR VPWR _0802_/A sky130_fd_sc_hd__inv_2
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1313_ hold46/A _1342_/A2 _1333_/B1 _1312_/X VGND VGND VPWR VPWR _1313_/X sky130_fd_sc_hd__o211a_1
X_1244_ hold16/A _1645_/Q _1244_/C VGND VGND VPWR VPWR _1248_/B sky130_fd_sc_hd__or3_1
X_1175_ _1180_/A _1175_/B VGND VGND VPWR VPWR _1555_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0959_ _0959_/A1 _0773_/Y _0945_/Y _0945_/B _1084_/A VGND VGND VPWR VPWR _0960_/B
+ sky130_fd_sc_hd__a32o_1
X_1449__85 _1454__90/A VGND VGND VPWR VPWR _1601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 uio_in[3] VGND VGND VPWR VPWR _1533_/D sky130_fd_sc_hd__clkbuf_1
X_0813_ _0829_/A _0829_/B _0829_/D VGND VGND VPWR VPWR _0818_/A sky130_fd_sc_hd__or3_1
XFILLER_0_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1227_ _1066_/X _1067_/Y _1236_/A _1226_/Y VGND VGND VPWR VPWR _1227_/X sky130_fd_sc_hd__a211o_1
X_1158_ _1148_/B _1162_/A VGND VGND VPWR VPWR _1158_/X sky130_fd_sc_hd__and2b_1
X_1089_ _1107_/A _1089_/B VGND VGND VPWR VPWR _1089_/X sky130_fd_sc_hd__or2_2
XFILLER_0_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1482__118 clkload8/A VGND VGND VPWR VPWR _1634_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1012_ _1610_/Q _1012_/B VGND VGND VPWR VPWR _1013_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1419__55 clkload5/A VGND VGND VPWR VPWR _1571_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1630_ _1630_/CLK _1630_/D VGND VGND VPWR VPWR _1630_/Q sky130_fd_sc_hd__dfxtp_1
X_1561_ _1561_/CLK _1561_/D VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout29 _0923_/A VGND VGND VPWR VPWR _0940_/A sky130_fd_sc_hd__clkbuf_2
X_1488__124 clkload1/A VGND VGND VPWR VPWR _1640_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0992_ hold37/X _0976_/Y _0978_/Y _1009_/C VGND VGND VPWR VPWR _1617_/D sky130_fd_sc_hd__o211a_1
X_1544_ _1544_/CLK _1544_/D VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfxtp_1
X_1613_ _1613_/CLK _1613_/D VGND VGND VPWR VPWR _1613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_7_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload6/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 ui_in[6] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1191_ _1188_/A _1187_/B _1189_/X VGND VGND VPWR VPWR _1258_/A sky130_fd_sc_hd__o21ai_1
X_1260_ _1260_/A _1260_/B VGND VGND VPWR VPWR _1260_/Y sky130_fd_sc_hd__nand2_1
X_0975_ _1030_/A _0977_/D VGND VGND VPWR VPWR _0993_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1527_ _1527_/CLK _1527_/D VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0760_ _1614_/Q VGND VGND VPWR VPWR _0760_/Y sky130_fd_sc_hd__inv_2
X_1174_ uo_out[5] _1173_/X _1179_/S VGND VGND VPWR VPWR _1175_/B sky130_fd_sc_hd__mux2_1
X_1312_ _1521_/Q _1337_/B VGND VGND VPWR VPWR _1312_/X sky130_fd_sc_hd__or2_1
X_1243_ _1646_/Q _1647_/Q _1648_/Q hold23/A VGND VGND VPWR VPWR _1244_/C sky130_fd_sc_hd__or4_1
X_0889_ _1616_/Q _1636_/Q VGND VGND VPWR VPWR _0889_/X sky130_fd_sc_hd__or2_1
X_0958_ _0960_/A _0958_/B VGND VGND VPWR VPWR _1628_/D sky130_fd_sc_hd__and2_1
X_1394__30 clkload4/A VGND VGND VPWR VPWR _1546_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0812_ _1607_/Q _0777_/Y _0833_/A _0830_/B _0831_/A VGND VGND VPWR VPWR _0825_/A
+ sky130_fd_sc_hd__a2111o_1
X_1226_ _1187_/B _1235_/B _1189_/X _1130_/D VGND VGND VPWR VPWR _1226_/Y sky130_fd_sc_hd__o211ai_1
X_1157_ _0903_/X _1260_/B _1148_/X _1530_/Q VGND VGND VPWR VPWR _1157_/X sky130_fd_sc_hd__a2bb2o_2
X_1088_ _1107_/A _1089_/B VGND VGND VPWR VPWR _1104_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ _1008_/B _1011_/B _1019_/C VGND VGND VPWR VPWR _1611_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ hold58/A hold53/A VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1560_ _1560_/CLK _1560_/D VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0991_ hold48/A _0981_/D _0979_/Y _1009_/C VGND VGND VPWR VPWR _1618_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1543_ _1543_/CLK _1543_/D VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfxtp_2
X_1612_ _1612_/CLK _1612_/D VGND VGND VPWR VPWR _1612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput9 ui_in[7] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
X_1190_ _1188_/A hold42/A VGND VGND VPWR VPWR _1235_/B sky130_fd_sc_hd__nand2b_1
X_0974_ _1612_/Q _1611_/Q _0998_/C _0974_/D VGND VGND VPWR VPWR _0977_/D sky130_fd_sc_hd__and4_1
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1526_ _1526_/CLK _1526_/D VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload5/A sky130_fd_sc_hd__clkbuf_8
X_1311_ hold46/X _1275_/Y _1310_/X _1336_/C1 VGND VGND VPWR VPWR _1523_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1242_ _1242_/A hold17/X VGND VGND VPWR VPWR _1542_/D sky130_fd_sc_hd__or2_1
X_1173_ _1349_/A _1172_/X _1178_/S VGND VGND VPWR VPWR _1173_/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0888_ _1613_/Q _0774_/Y _1635_/Q _0759_/Y _0887_/X VGND VGND VPWR VPWR _0888_/X
+ sky130_fd_sc_hd__a221o_1
X_0957_ _0959_/A1 _1628_/Q _0945_/Y _0945_/B hold26/A VGND VGND VPWR VPWR _0958_/B
+ sky130_fd_sc_hd__a32o_1
X_1509_ _1509_/CLK _1509_/D VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0811_ _0802_/A _1651_/Q _1654_/Q _0993_/A VGND VGND VPWR VPWR _0830_/B sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1156_ _1153_/X _1154_/X _1155_/X _1080_/A VGND VGND VPWR VPWR _1260_/B sky130_fd_sc_hd__o22ai_1
X_1225_ _1188_/A hold42/A _1066_/X _1186_/Y _1231_/B VGND VGND VPWR VPWR _1236_/A
+ sky130_fd_sc_hd__a32o_1
X_1087_ _1349_/B _1192_/A _1086_/X _1117_/C1 VGND VGND VPWR VPWR _1582_/D sky130_fd_sc_hd__o211a_1
X_1454__90 _1454__90/A VGND VGND VPWR VPWR _1606_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ _1611_/Q _1010_/B VGND VGND VPWR VPWR _1011_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1208_ hold53/A hold58/A VGND VGND VPWR VPWR _1208_/Y sky130_fd_sc_hd__nand2b_1
X_1139_ _1139_/A _1141_/A VGND VGND VPWR VPWR _1562_/D sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_26_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1424__60 clkload5/A VGND VGND VPWR VPWR _1576_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_13_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1472__108 clkload0/A VGND VGND VPWR VPWR _1624_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1611_ _1611_/CLK _1611_/D VGND VGND VPWR VPWR _1611_/Q sky130_fd_sc_hd__dfxtp_1
X_0990_ _0980_/X _1009_/C _0990_/C VGND VGND VPWR VPWR _1619_/D sky130_fd_sc_hd__and3b_1
X_1542_ _1542_/CLK _1542_/D VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1494__130 clkload10/A VGND VGND VPWR VPWR _1646_/CLK sky130_fd_sc_hd__inv_2
X_0973_ _1615_/Q _1614_/Q _1613_/Q _1610_/Q VGND VGND VPWR VPWR _0974_/D sky130_fd_sc_hd__and4_1
X_1525_ _1525_/CLK _1525_/D VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1478__114 clkload10/A VGND VGND VPWR VPWR _1630_/CLK sky130_fd_sc_hd__inv_2
X_1310_ _1178_/S _1309_/X _1308_/X _1344_/C1 VGND VGND VPWR VPWR _1310_/X sky130_fd_sc_hd__a211o_1
X_1241_ hold42/A _1130_/D _1239_/X _1240_/X _1199_/A VGND VGND VPWR VPWR _1543_/D
+ sky130_fd_sc_hd__o221a_1
X_1172_ _1157_/X uo_out[5] _1172_/S VGND VGND VPWR VPWR _1172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ _0956_/A _0956_/B VGND VGND VPWR VPWR _1629_/D sky130_fd_sc_hd__and2_1
X_0887_ _0759_/Y _1635_/Q _1637_/Q _0757_/Y VGND VGND VPWR VPWR _0887_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1385__21 clkload13/A VGND VGND VPWR VPWR _1528_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_1_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0810_ _1615_/Q _1653_/Q VGND VGND VPWR VPWR _0831_/D sky130_fd_sc_hd__and2b_1
X_1224_ _1224_/A _1224_/B VGND VGND VPWR VPWR _1231_/B sky130_fd_sc_hd__nor2_1
X_1155_ uo_out[4] uo_out[5] uo_out[6] uo_out[7] _1349_/B _1149_/A VGND VGND VPWR VPWR
+ _1155_/X sky130_fd_sc_hd__mux4_1
X_1086_ _1533_/Q _1086_/B VGND VGND VPWR VPWR _1086_/X sky130_fd_sc_hd__or2_1
X_0939_ _0937_/X _0938_/X _0855_/A VGND VGND VPWR VPWR _1636_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_5_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload4/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1207_ _1207_/A _1207_/B VGND VGND VPWR VPWR _1207_/Y sky130_fd_sc_hd__nor2_1
X_1069_ _1546_/Q hold54/A VGND VGND VPWR VPWR _1234_/A sky130_fd_sc_hd__and2b_1
X_1138_ _1138_/A hold22/X VGND VGND VPWR VPWR _1563_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1610_ _1610_/CLK _1610_/D VGND VGND VPWR VPWR _1610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ _1541_/CLK input9/X VGND VGND VPWR VPWR _1541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0972_ _1609_/Q _1608_/Q _1607_/Q VGND VGND VPWR VPWR _0998_/C sky130_fd_sc_hd__and3_1
X_1524_ _1524_/CLK _1524_/D VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1171_ _1201_/B _1355_/A VGND VGND VPWR VPWR _1172_/S sky130_fd_sc_hd__nand2_1
X_1240_ _1546_/Q _1067_/Y _1126_/Y _1127_/X _1230_/X VGND VGND VPWR VPWR _1240_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ _0882_/X _0883_/Y _0884_/Y _0885_/X _0881_/X VGND VGND VPWR VPWR _0897_/B
+ sky130_fd_sc_hd__a221o_1
X_0955_ _0955_/A1 _1629_/Q _0945_/Y _0945_/B _1176_/A VGND VGND VPWR VPWR _0956_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1154_ uo_out[0] _1358_/A _1355_/A uo_out[1] _1151_/X VGND VGND VPWR VPWR _1154_/X
+ sky130_fd_sc_hd__a221o_1
X_1223_ hold47/A hold43/A hold50/A hold49/A VGND VGND VPWR VPWR _1224_/B sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1085_ hold26/X _1084_/B _1084_/Y _0960_/A VGND VGND VPWR VPWR _1583_/D sky130_fd_sc_hd__o211a_1
X_0938_ _1149_/A _0941_/B VGND VGND VPWR VPWR _0938_/X sky130_fd_sc_hd__and2_1
X_0869_ _0959_/A1 _0778_/Y _0857_/Y wire19/X _1082_/A VGND VGND VPWR VPWR _0870_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1445__81 _1454__90/A VGND VGND VPWR VPWR _1597_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1206_ hold9/A hold27/A hold21/A hold34/A VGND VGND VPWR VPWR _1207_/B sky130_fd_sc_hd__or4_1
X_1137_ hold34/A _1141_/A hold21/X VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_35_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1068_ _1188_/A hold42/A VGND VGND VPWR VPWR _1187_/A sky130_fd_sc_hd__or2_1
XFILLER_0_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload3/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1415__51 clkload6/A VGND VGND VPWR VPWR _1567_/CLK sky130_fd_sc_hd__inv_2
X_1540_ _1541_/CLK input8/X VGND VGND VPWR VPWR _1540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1669_ hold17/A VGND VGND VPWR VPWR uio_oe[2] sky130_fd_sc_hd__buf_2
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1367__3 clkload6/A VGND VGND VPWR VPWR _1510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0971_ _0971_/A _0971_/B VGND VGND VPWR VPWR _1623_/D sky130_fd_sc_hd__and2_1
X_1503__139 clkload7/A VGND VGND VPWR VPWR _1655_/CLK sky130_fd_sc_hd__inv_2
X_1523_ _1523_/CLK _1523_/D VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ uo_out[6] _1179_/S _1168_/X _1169_/Y _1180_/A VGND VGND VPWR VPWR _1556_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ _1612_/Q _1632_/Q VGND VGND VPWR VPWR _0885_/X sky130_fd_sc_hd__or2_1
X_0954_ _0960_/A _0954_/B VGND VGND VPWR VPWR _1630_/D sky130_fd_sc_hd__and2_1
X_1299_ hold41/A hold40/A _1339_/S VGND VGND VPWR VPWR _1299_/X sky130_fd_sc_hd__mux2_1
X_1484__120 clkload1/A VGND VGND VPWR VPWR _1636_/CLK sky130_fd_sc_hd__inv_2
Xtt_um_jimktrains_vslc_64 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_64/HI uio_oe[3]
+ sky130_fd_sc_hd__conb_1
X_1376__12 _1533_/CLK VGND VGND VPWR VPWR _1519_/CLK sky130_fd_sc_hd__inv_2
X_1153_ uo_out[2] _1352_/A _1176_/A VGND VGND VPWR VPWR _1153_/X sky130_fd_sc_hd__a21o_1
X_1222_ hold51/A hold57/A hold56/A hold45/A VGND VGND VPWR VPWR _1224_/A sky130_fd_sc_hd__or4_1
X_1468__104 clkload7/A VGND VGND VPWR VPWR _1620_/CLK sky130_fd_sc_hd__inv_2
X_1084_ _1084_/A _1084_/B VGND VGND VPWR VPWR _1084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0937_ _0940_/A _1636_/Q _0940_/C VGND VGND VPWR VPWR _0937_/X sky130_fd_sc_hd__and3_1
X_0799_ _1622_/Q _1660_/Q VGND VGND VPWR VPWR _0833_/A sky130_fd_sc_hd__xor2_1
X_0868_ _0960_/A _0868_/B VGND VGND VPWR VPWR _1647_/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1460__96 clkload9/A VGND VGND VPWR VPWR _1612_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1067_ _1188_/A hold42/A VGND VGND VPWR VPWR _1067_/Y sky130_fd_sc_hd__nor2_1
X_1136_ _1136_/A _1138_/A VGND VGND VPWR VPWR _1564_/D sky130_fd_sc_hd__xnor2_1
X_1205_ hold18/A hold19/A hold58/A _1558_/Q VGND VGND VPWR VPWR _1207_/A sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ _1201_/B _1107_/X _1118_/X _1180_/A VGND VGND VPWR VPWR _1568_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1430__66 _1372__8/A VGND VGND VPWR VPWR _1582_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1668_ hold17/A VGND VGND VPWR VPWR uio_oe[1] sky130_fd_sc_hd__buf_2
X_1599_ _1599_/CLK _1599_/D VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload2/A sky130_fd_sc_hd__clkbuf_8
X_0970_ _0940_/A _1623_/Q _0963_/Y wire17/X _0941_/A VGND VGND VPWR VPWR _0971_/B
+ sky130_fd_sc_hd__a32o_1
X_1522_ _1522_/CLK _1522_/D VGND VGND VPWR VPWR _1522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1400__36 clkload3/A VGND VGND VPWR VPWR _1552_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0884_ _1612_/Q _1632_/Q VGND VGND VPWR VPWR _0884_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0953_ _0959_/A1 _1630_/Q _0945_/Y _0945_/B _1348_/D VGND VGND VPWR VPWR _0954_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1298_ hold41/A _0913_/Y _1333_/B1 _1297_/X VGND VGND VPWR VPWR _1298_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_18_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_jimktrains_vslc_65 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_65/HI uio_oe[4]
+ sky130_fd_sc_hd__conb_1
X_1391__27 clkload3/A VGND VGND VPWR VPWR _1543_/CLK sky130_fd_sc_hd__inv_2
X_1221_ _1207_/Y _1221_/B _1221_/C VGND VGND VPWR VPWR _1221_/X sky130_fd_sc_hd__and3b_1
X_1152_ _1149_/A _1349_/B VGND VGND VPWR VPWR _1355_/A sky130_fd_sc_hd__and2b_2
X_1083_ _1176_/A _1192_/A _1082_/Y _0960_/A VGND VGND VPWR VPWR _1584_/D sky130_fd_sc_hd__o211a_1
X_0936_ _0934_/X _0935_/X _0855_/A VGND VGND VPWR VPWR _1637_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0798_ _1609_/Q _1647_/Q VGND VGND VPWR VPWR _0829_/C sky130_fd_sc_hd__and2b_1
X_0867_ _0955_/A1 _1647_/Q _0857_/Y wire19/X _1176_/A VGND VGND VPWR VPWR _0868_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_38_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1436__72 clkload5/A VGND VGND VPWR VPWR _1588_/CLK sky130_fd_sc_hd__inv_2
X_1204_ _1188_/A hold42/A _1234_/A VGND VGND VPWR VPWR _1221_/C sky130_fd_sc_hd__and3b_1
XFILLER_0_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1066_ hold54/A _1546_/Q VGND VGND VPWR VPWR _1066_/X sky130_fd_sc_hd__and2b_1
X_1135_ hold9/X _1135_/B VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0919_ _0944_/A _1089_/B _0963_/A VGND VGND VPWR VPWR _0940_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1118_ hold57/X _1122_/B VGND VGND VPWR VPWR _1118_/X sky130_fd_sc_hd__or2_1
X_1049_ _1049_/A _1049_/B VGND VGND VPWR VPWR _1597_/D sky130_fd_sc_hd__nor2_1
X_1406__42 clkload3/A VGND VGND VPWR VPWR _1558_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1667_ hold17/A VGND VGND VPWR VPWR uio_oe[0] sky130_fd_sc_hd__buf_2
X_1598_ _1598_/CLK _1598_/D VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_34_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1521_ _1521_/CLK _1521_/D VGND VGND VPWR VPWR _1521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1397__33 clkload4/A VGND VGND VPWR VPWR _1549_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ hold6/X _1251_/A _0945_/Y _0945_/B _0843_/X VGND VGND VPWR VPWR _1631_/D sky130_fd_sc_hd__a32o_1
X_0883_ _1610_/Q _1630_/Q VGND VGND VPWR VPWR _0883_/Y sky130_fd_sc_hd__nand2_1
X_1366_ hold11/A _1366_/B VGND VGND VPWR VPWR _1672_/A sky130_fd_sc_hd__nor2_2
X_1297_ hold40/A _1337_/B VGND VGND VPWR VPWR _1297_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload1/A sky130_fd_sc_hd__clkbuf_8
Xtt_um_jimktrains_vslc_66 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_66/HI uio_oe[5]
+ sky130_fd_sc_hd__conb_1
X_1151_ _1349_/A _1349_/B uo_out[3] VGND VGND VPWR VPWR _1151_/X sky130_fd_sc_hd__and3_1
X_1220_ _1207_/Y _1221_/B VGND VGND VPWR VPWR _1220_/Y sky130_fd_sc_hd__nand2b_1
X_1082_ _1082_/A _1084_/B VGND VGND VPWR VPWR _1082_/Y sky130_fd_sc_hd__nand2_1
X_0935_ _1201_/B _0941_/B VGND VGND VPWR VPWR _0935_/X sky130_fd_sc_hd__and2_1
X_0866_ _0960_/A _0866_/B VGND VGND VPWR VPWR _1648_/D sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_21_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0797_ _1608_/Q _1646_/Q VGND VGND VPWR VPWR _0834_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1349_ _1349_/A _1349_/B _1358_/B VGND VGND VPWR VPWR _1350_/S sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_38_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1451__87 _1454__90/A VGND VGND VPWR VPWR _1603_/CLK sky130_fd_sc_hd__inv_2
X_1474__110 clkload0/A VGND VGND VPWR VPWR _1626_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1203_ _1355_/A _1203_/B VGND VGND VPWR VPWR _1203_/Y sky130_fd_sc_hd__nand2_1
X_1134_ hold27/A _1138_/A VGND VGND VPWR VPWR _1135_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1065_ _1351_/A _1065_/B _1065_/C VGND VGND VPWR VPWR _1590_/D sky130_fd_sc_hd__and3_1
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0849_ _0956_/A _0849_/B VGND VGND VPWR VPWR _1656_/D sky130_fd_sc_hd__and2_1
X_0918_ _1550_/Q hold55/A VGND VGND VPWR VPWR _1089_/B sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_3_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1117_ _1348_/D _1107_/X _1116_/X _1117_/C1 VGND VGND VPWR VPWR _1569_/D sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ hold7/X _1022_/X _1051_/B VGND VGND VPWR VPWR _1049_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421__57 clkload5/A VGND VGND VPWR VPWR _1573_/CLK sky130_fd_sc_hd__inv_2
X_1597_ _1597_/CLK _1597_/D VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1520_ _1520_/CLK _1520_/D VGND VGND VPWR VPWR _1520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1649_ _1649_/CLK _1649_/D VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0882_ _1610_/Q _1630_/Q VGND VGND VPWR VPWR _0882_/X sky130_fd_sc_hd__or2_1
X_0951_ _0960_/A _0951_/B VGND VGND VPWR VPWR _1632_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1365_ hold11/X _1189_/X _1236_/C _1242_/A VGND VGND VPWR VPWR _1509_/D sky130_fd_sc_hd__a211o_1
X_1296_ hold41/X _1345_/A2 _1295_/X _1336_/C1 VGND VGND VPWR VPWR _1526_/D sky130_fd_sc_hd__o211a_1
X_1457__93 clkload9/A VGND VGND VPWR VPWR _1609_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1491__127 _1372__8/A VGND VGND VPWR VPWR _1643_/CLK sky130_fd_sc_hd__inv_2
Xtt_um_jimktrains_vslc_67 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_67/HI uio_out[3]
+ sky130_fd_sc_hd__conb_1
X_1150_ _1264_/B _1349_/A VGND VGND VPWR VPWR _1352_/A sky130_fd_sc_hd__and2b_2
X_0781__1 clkload4/A VGND VGND VPWR VPWR _1509_/CLK sky130_fd_sc_hd__inv_2
X_1081_ _1348_/D _1192_/A _1080_/Y _1351_/A VGND VGND VPWR VPWR _1585_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0934_ _0940_/A _1637_/Q _0940_/C VGND VGND VPWR VPWR _0934_/X sky130_fd_sc_hd__and3_1
X_0865_ _0959_/A1 _1648_/Q _0857_/Y wire19/X _1348_/D VGND VGND VPWR VPWR _0866_/B
+ sky130_fd_sc_hd__a32o_1
X_0796_ _1654_/Q _1616_/Q VGND VGND VPWR VPWR _0829_/B sky130_fd_sc_hd__and2b_1
X_1382__18 clkload13/A VGND VGND VPWR VPWR _1525_/CLK sky130_fd_sc_hd__inv_2
X_1348_ _1201_/B _1346_/C _1348_/C _1348_/D VGND VGND VPWR VPWR _1358_/B sky130_fd_sc_hd__and4bb_2
X_1279_ _1590_/Q hold39/A _1334_/S VGND VGND VPWR VPWR _1279_/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1202_ _1202_/A VGND VGND VPWR VPWR _1203_/B sky130_fd_sc_hd__inv_2
X_1064_ _0906_/C _1061_/Y _1590_/Q VGND VGND VPWR VPWR _1065_/C sky130_fd_sc_hd__a21o_1
Xclkbuf_4_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload0/A sky130_fd_sc_hd__clkbuf_8
X_1133_ hold21/A hold34/A _1141_/A VGND VGND VPWR VPWR _1138_/A sky130_fd_sc_hd__and3_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1427__63 clkload0/A VGND VGND VPWR VPWR _1579_/CLK sky130_fd_sc_hd__inv_2
X_0779_ hold23/A VGND VGND VPWR VPWR _0807_/B sky130_fd_sc_hd__inv_2
X_0848_ _0955_/A1 _1656_/Q _0836_/Y _0836_/A _1348_/D VGND VGND VPWR VPWR _0849_/B
+ sky130_fd_sc_hd__a32o_1
X_0917_ _1550_/Q _0944_/A hold55/A VGND VGND VPWR VPWR _0941_/B sky130_fd_sc_hd__nor3b_2
XTAP_TAPCELL_ROW_3_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1497__133 clkload10/A VGND VGND VPWR VPWR _1649_/CLK sky130_fd_sc_hd__inv_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1116_ hold51/X _1122_/B VGND VGND VPWR VPWR _1116_/X sky130_fd_sc_hd__or2_1
X_1047_ _1047_/A _1047_/B VGND VGND VPWR VPWR _1598_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ _1596_/CLK _1596_/D VGND VGND VPWR VPWR _1596_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1579_ _1579_/CLK _1579_/D VGND VGND VPWR VPWR _1579_/Q sky130_fd_sc_hd__dfxtp_1
X_1648_ _1648_/CLK _1648_/D VGND VGND VPWR VPWR _1648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1388__24 clkload6/A VGND VGND VPWR VPWR _1531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0881_ _1607_/Q _1627_/Q VGND VGND VPWR VPWR _0881_/X sky130_fd_sc_hd__xor2_1
X_0950_ _0959_/A1 _1632_/Q _0945_/Y _0945_/B _1346_/A VGND VGND VPWR VPWR _0951_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1364_ _1257_/A _1361_/X _1363_/X _1180_/A VGND VGND VPWR VPWR _1510_/D sky130_fd_sc_hd__o211a_1
X_1295_ _1340_/A1 _1294_/X _1293_/X _1276_/X VGND VGND VPWR VPWR _1295_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_18_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_jimktrains_vslc_68 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_68/HI uio_out[4]
+ sky130_fd_sc_hd__conb_1
X_1080_ _1080_/A _1192_/A VGND VGND VPWR VPWR _1080_/Y sky130_fd_sc_hd__nand2_1
X_0781__2 clkload4/A VGND VGND VPWR VPWR _1366_/B sky130_fd_sc_hd__inv_2
XFILLER_0_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0795_ hold20/A _1619_/Q VGND VGND VPWR VPWR _0831_/B sky130_fd_sc_hd__and2b_1
X_0933_ _0931_/X _0932_/X _0855_/A VGND VGND VPWR VPWR _1638_/D sky130_fd_sc_hd__o21a_1
X_0864_ hold23/X _1251_/A _0857_/Y wire19/X _0843_/X VGND VGND VPWR VPWR _1649_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1347_ _0941_/A hold16/X _1347_/S VGND VGND VPWR VPWR _1515_/D sky130_fd_sc_hd__mux2_1
X_1278_ _1590_/Q _1342_/A2 _1333_/B1 _1277_/X VGND VGND VPWR VPWR _1278_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_29_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1201_ _1348_/D _1201_/B _1201_/C _1346_/D VGND VGND VPWR VPWR _1202_/A sky130_fd_sc_hd__or4_2
X_1132_ hold18/A _1143_/A VGND VGND VPWR VPWR _1141_/A sky130_fd_sc_hd__and2_1
X_1063_ _1063_/A hold32/A _0906_/C VGND VGND VPWR VPWR _1065_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0916_ _0910_/X _0915_/X _1351_/A VGND VGND VPWR VPWR _1643_/D sky130_fd_sc_hd__o21a_1
X_1442__78 clkload1/A VGND VGND VPWR VPWR _1594_/CLK sky130_fd_sc_hd__inv_2
X_0847_ hold20/X _0836_/Y _1251_/A _0843_/X _0836_/A VGND VGND VPWR VPWR _1657_/D
+ sky130_fd_sc_hd__a32o_1
X_0778_ _1646_/Q VGND VGND VPWR VPWR _0778_/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1115_ _1076_/A _1107_/X _1114_/X _1117_/C1 VGND VGND VPWR VPWR _1570_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1046_ hold28/X _1049_/A _1051_/B VGND VGND VPWR VPWR _1047_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1464__100 clkload7/A VGND VGND VPWR VPWR _1616_/CLK sky130_fd_sc_hd__inv_2
X_1372__8 _1372__8/A VGND VGND VPWR VPWR _1515_/CLK sky130_fd_sc_hd__inv_2
X_1505__141 clkload8/A VGND VGND VPWR VPWR _1657_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1454__90/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1595_ _1595_/CLK _1595_/D VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1412__48 clkload0/A VGND VGND VPWR VPWR _1564_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1029_ hold4/A _1605_/Q _1037_/A VGND VGND VPWR VPWR _1029_/X sky130_fd_sc_hd__and3_1
XFILLER_0_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1578_ _1578_/CLK _1578_/D VGND VGND VPWR VPWR _1578_/Q sky130_fd_sc_hd__dfxtp_1
X_1647_ _1647_/CLK _1647_/D VGND VGND VPWR VPWR _1647_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_38_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ _0762_/Y _1629_/Q _0873_/X _0879_/X VGND VGND VPWR VPWR _0897_/A sky130_fd_sc_hd__a211o_1
X_1363_ hold38/A _1363_/B VGND VGND VPWR VPWR _1363_/X sky130_fd_sc_hd__or2_1
X_1294_ hold44/A hold52/A _1339_/S VGND VGND VPWR VPWR _1294_/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_jimktrains_vslc_69 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_69/HI uio_out[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_5_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1448__84 _1454__90/A VGND VGND VPWR VPWR _1600_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0932_ _1260_/A _0941_/B VGND VGND VPWR VPWR _0932_/X sky130_fd_sc_hd__and2_1
XFILLER_0_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0794_ _1612_/Q _1650_/Q VGND VGND VPWR VPWR _0829_/A sky130_fd_sc_hd__and2b_1
X_0863_ _0956_/A _0863_/B VGND VGND VPWR VPWR _1650_/D sky130_fd_sc_hd__and2_1
X_1346_ _1346_/A _1346_/B _1346_/C _1346_/D VGND VGND VPWR VPWR _1347_/S sky130_fd_sc_hd__or4_1
X_1277_ hold39/A _1337_/B VGND VGND VPWR VPWR _1277_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_29_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ _1547_/Q _1193_/B _1199_/Y VGND VGND VPWR VPWR _1547_/D sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_25_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1481__117 clkload8/A VGND VGND VPWR VPWR _1633_/CLK sky130_fd_sc_hd__inv_2
X_1131_ hold19/A hold58/A _1146_/A VGND VGND VPWR VPWR _1143_/A sky130_fd_sc_hd__and3_1
X_1062_ _1148_/B _1346_/C VGND VGND VPWR VPWR _1063_/A sky130_fd_sc_hd__or2_1
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ _0910_/B _1201_/C _0915_/C VGND VGND VPWR VPWR _0915_/X sky130_fd_sc_hd__and3b_1
X_0846_ _0855_/A _0923_/A VGND VGND VPWR VPWR _1030_/B sky130_fd_sc_hd__nand2_1
X_0777_ _1645_/Q VGND VGND VPWR VPWR _0777_/Y sky130_fd_sc_hd__inv_2
X_1329_ _1520_/Q _1518_/Q _1334_/S VGND VGND VPWR VPWR _1329_/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1418__54 clkload5/A VGND VGND VPWR VPWR _1570_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
X_1114_ hold49/X _1122_/B VGND VGND VPWR VPWR _1114_/X sky130_fd_sc_hd__or2_1
X_1045_ _1045_/A _1045_/B VGND VGND VPWR VPWR _1599_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0829_ _0829_/A _0829_/B _0829_/C _0829_/D VGND VGND VPWR VPWR _0830_/D sky130_fd_sc_hd__or4_1
XFILLER_0_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1594_ _1594_/CLK _1594_/D VGND VGND VPWR VPWR _1594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1487__123 clkload2/A VGND VGND VPWR VPWR _1639_/CLK sky130_fd_sc_hd__inv_2
X_1028_ hold25/A _1028_/B VGND VGND VPWR VPWR _1037_/A sky130_fd_sc_hd__and2_1
XFILLER_0_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1646_ _1646_/CLK _1646_/D VGND VGND VPWR VPWR _1646_/Q sky130_fd_sc_hd__dfxtp_1
X_1577_ _1577_/CLK _1577_/D VGND VGND VPWR VPWR _1577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1379__15 _1541_/CLK VGND VGND VPWR VPWR _1522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_10_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1362_ _1522_/Q _1521_/Q _1520_/Q _1519_/Q _1547_/Q _1548_/Q VGND VGND VPWR VPWR
+ _1363_/B sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_2_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1293_ hold44/A _1342_/A2 _1333_/B1 _1292_/X VGND VGND VPWR VPWR _1293_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1629_ _1629_/CLK _1629_/D VGND VGND VPWR VPWR _1629_/Q sky130_fd_sc_hd__dfxtp_1
X_1463__99 clkload9/A VGND VGND VPWR VPWR _1615_/CLK sky130_fd_sc_hd__inv_2
X_0931_ _0940_/A _1638_/Q _0940_/C VGND VGND VPWR VPWR _0931_/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_15_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0862_ _0955_/A1 _1650_/Q _0857_/Y wire19/X _1346_/A VGND VGND VPWR VPWR _0863_/B
+ sky130_fd_sc_hd__a32o_1
X_0793_ _1610_/Q _1648_/Q VGND VGND VPWR VPWR _0834_/A sky130_fd_sc_hd__and2b_1
X_1345_ _1516_/Q _1345_/A2 _1344_/X _1351_/A VGND VGND VPWR VPWR _1516_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_3_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1276_ _1162_/A _1162_/C _1063_/A VGND VGND VPWR VPWR _1276_/X sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_29_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1130_ _1199_/A _1558_/Q _1192_/A _1130_/D VGND VGND VPWR VPWR _1146_/A sky130_fd_sc_hd__and4_1
XFILLER_0_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1061_ _1148_/B _1346_/C VGND VGND VPWR VPWR _1061_/Y sky130_fd_sc_hd__nor2_1
X_0845_ _0845_/A _0923_/A VGND VGND VPWR VPWR _1251_/A sky130_fd_sc_hd__and2_1
X_0914_ _1530_/Q _1337_/B VGND VGND VPWR VPWR _0915_/C sky130_fd_sc_hd__or2_1
XFILLER_0_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0776_ _1641_/Q VGND VGND VPWR VPWR _0776_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ hold8/X _1258_/A _1255_/X _1258_/Y _1259_/C1 VGND VGND VPWR VPWR _1531_/D
+ sky130_fd_sc_hd__o221a_1
X_1328_ _1520_/Q _1342_/A2 _1333_/B1 _1327_/X VGND VGND VPWR VPWR _1328_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1433__69 _1372__8/A VGND VGND VPWR VPWR _1585_/CLK sky130_fd_sc_hd__inv_2
X_1113_ _1162_/B _1107_/X _1112_/X _1117_/C1 VGND VGND VPWR VPWR _1571_/D sky130_fd_sc_hd__o211a_1
X_1044_ hold14/X _1047_/A _1060_/B VGND VGND VPWR VPWR _1045_/B sky130_fd_sc_hd__o21ai_1
X_0759_ _1615_/Q VGND VGND VPWR VPWR _0759_/Y sky130_fd_sc_hd__inv_2
X_0828_ _1607_/Q _0777_/Y _0823_/B _0823_/C _0824_/C VGND VGND VPWR VPWR _0830_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_22_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1593_ _1593_/CLK _1593_/D VGND VGND VPWR VPWR _1593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ hold5/A _1602_/Q _1043_/A VGND VGND VPWR VPWR _1028_/B sky130_fd_sc_hd__and3_1
X_1403__39 clkload6/A VGND VGND VPWR VPWR _1555_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1576_ _1576_/CLK _1576_/D VGND VGND VPWR VPWR _1576_/Q sky130_fd_sc_hd__dfxtp_1
X_1645_ _1645_/CLK _1645_/D VGND VGND VPWR VPWR _1645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1361_ _1518_/Q _1517_/Q _1516_/Q _1530_/Q _1547_/Q _1548_/Q VGND VGND VPWR VPWR
+ _1361_/X sky130_fd_sc_hd__mux4_1
X_1292_ hold52/A _1337_/B VGND VGND VPWR VPWR _1292_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1628_ _1628_/CLK _1628_/D VGND VGND VPWR VPWR _1628_/Q sky130_fd_sc_hd__dfxtp_1
X_1559_ _1559_/CLK _1559_/D VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1439__75 clkload1/A VGND VGND VPWR VPWR _1591_/CLK sky130_fd_sc_hd__inv_2
X_0792_ _0787_/Y _0788_/Y _0791_/X _1626_/Q VGND VGND VPWR VPWR _1030_/A sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_15_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0930_ _0843_/X _0941_/B _0929_/X VGND VGND VPWR VPWR _1639_/D sky130_fd_sc_hd__a21o_1
X_0861_ _0956_/A _0861_/B VGND VGND VPWR VPWR _1651_/D sky130_fd_sc_hd__and2_1
X_1344_ _1178_/S _1343_/X _1342_/X _1344_/C1 VGND VGND VPWR VPWR _1344_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1275_ _1162_/A _1162_/C _1063_/A VGND VGND VPWR VPWR _1275_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1060_ hold29/A _1060_/B VGND VGND VPWR VPWR _1591_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_34_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0775_ _1638_/Q VGND VGND VPWR VPWR _0775_/Y sky130_fd_sc_hd__inv_2
X_0844_ _0845_/A _1076_/A VGND VGND VPWR VPWR _1346_/B sky130_fd_sc_hd__nand2_1
X_0913_ _1162_/C _1346_/A VGND VGND VPWR VPWR _0913_/Y sky130_fd_sc_hd__nand2b_2
X_1258_ _1258_/A _1258_/B VGND VGND VPWR VPWR _1258_/Y sky130_fd_sc_hd__nand2_1
X_1189_ _1235_/A _1189_/B VGND VGND VPWR VPWR _1189_/X sky130_fd_sc_hd__or2_1
X_1327_ _1518_/Q _1337_/B VGND VGND VPWR VPWR _1327_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1409__45 clkload3/A VGND VGND VPWR VPWR _1561_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1043_ _1043_/A _1043_/B VGND VGND VPWR VPWR _1600_/D sky130_fd_sc_hd__nor2_1
X_1112_ hold50/X _1122_/B VGND VGND VPWR VPWR _1112_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0758_ _1616_/Q VGND VGND VPWR VPWR _0993_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ hold16/A _1030_/A wire18/X VGND VGND VPWR VPWR _0963_/A sky130_fd_sc_hd__and3_2
XFILLER_0_19_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1471__107 clkload0/A VGND VGND VPWR VPWR _1623_/CLK sky130_fd_sc_hd__inv_2
X_1592_ _1592_/CLK hold30/X VGND VGND VPWR VPWR _1592_/Q sky130_fd_sc_hd__dfxtp_1
X_1026_ hold31/A _1045_/A VGND VGND VPWR VPWR _1043_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1644_ _1644_/CLK _1644_/D VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfxtp_1
X_1575_ _1575_/CLK _1575_/D VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ _1006_/B _1009_/B _1009_/C VGND VGND VPWR VPWR _1612_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1477__113 clkload8/A VGND VGND VPWR VPWR _1629_/CLK sky130_fd_sc_hd__inv_2
X_1360_ _1157_/X _1358_/Y _1359_/X _1351_/A VGND VGND VPWR VPWR _1511_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_2_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1291_ hold44/X _1345_/A2 _1290_/X _1336_/C1 VGND VGND VPWR VPWR _1527_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1627_ _1627_/CLK _1627_/D VGND VGND VPWR VPWR _1627_/Q sky130_fd_sc_hd__dfxtp_1
X_1558_ _1558_/CLK _1558_/D VGND VGND VPWR VPWR _1558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1384__20 clkload13/A VGND VGND VPWR VPWR _1527_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ _0789_/X _0790_/X _1625_/Q VGND VGND VPWR VPWR _0791_/X sky130_fd_sc_hd__mux2_1
X_0860_ _0955_/A1 _1651_/Q _0857_/Y wire19/X _1148_/B VGND VGND VPWR VPWR _0861_/B
+ sky130_fd_sc_hd__a32o_1
X_1343_ _1530_/Q _1517_/Q _1348_/C VGND VGND VPWR VPWR _1343_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1274_ _1530_/Q _1061_/Y _1273_/X _1351_/A VGND VGND VPWR VPWR _1530_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0989_ hold48/A _0981_/D _1619_/Q VGND VGND VPWR VPWR _0990_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ _1076_/A _1346_/A VGND VGND VPWR VPWR _1322_/B sky130_fd_sc_hd__and2b_1
X_0774_ _1633_/Q VGND VGND VPWR VPWR _0774_/Y sky130_fd_sc_hd__inv_2
X_0843_ _0845_/A _1076_/A VGND VGND VPWR VPWR _0843_/X sky130_fd_sc_hd__and2_1
X_1326_ _1520_/Q _1345_/A2 _1325_/X _1331_/C1 VGND VGND VPWR VPWR _1520_/D sky130_fd_sc_hd__o211a_1
X_1257_ _1257_/A _1257_/B _1256_/X VGND VGND VPWR VPWR _1258_/B sky130_fd_sc_hd__or3b_1
X_1188_ _1188_/A hold42/A VGND VGND VPWR VPWR _1189_/B sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1111_ _1072_/A _1107_/X _1110_/X _1117_/C1 VGND VGND VPWR VPWR _1572_/D sky130_fd_sc_hd__o211a_1
X_1042_ hold31/X _1045_/A _1051_/B VGND VGND VPWR VPWR _1043_/B sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_31_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0757_ hold37/A VGND VGND VPWR VPWR _0757_/Y sky130_fd_sc_hd__inv_2
X_0826_ hold16/A wire18/X VGND VGND VPWR VPWR _0826_/X sky130_fd_sc_hd__and2_1
Xclkbuf_4_15_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1541_/CLK sky130_fd_sc_hd__clkbuf_8
X_1309_ hold40/A _1522_/Q _1334_/S VGND VGND VPWR VPWR _1309_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1591_ _1591_/CLK _1591_/D VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1660_ _1660_/CLK _1660_/D VGND VGND VPWR VPWR _1660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1025_ hold28/A hold14/A _1049_/A VGND VGND VPWR VPWR _1045_/A sky130_fd_sc_hd__and3_1
X_0809_ _1647_/Q _1609_/Q VGND VGND VPWR VPWR _0829_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1643_ _1643_/CLK _1643_/D VGND VGND VPWR VPWR _1643_/Q sky130_fd_sc_hd__dfxtp_1
X_1574_ _1574_/CLK _1574_/D VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_16_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ _1612_/Q _1008_/B VGND VGND VPWR VPWR _1009_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ _1340_/A1 _1289_/X _1288_/X _1276_/X VGND VGND VPWR VPWR _1290_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1626_ _1626_/CLK _1626_/D VGND VGND VPWR VPWR _1626_/Q sky130_fd_sc_hd__dfxtp_1
X_1557_ _1557_/CLK _1557_/D VGND VGND VPWR VPWR uo_out[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0790_ hold15/A _1596_/Q hold7/A hold28/A _1623_/Q _1624_/Q VGND VGND VPWR VPWR _0790_/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1342_ _1517_/Q _1342_/A2 _0915_/C _1342_/C1 VGND VGND VPWR VPWR _1342_/X sky130_fd_sc_hd__o211a_1
X_1273_ _1268_/X _1272_/X _1063_/A VGND VGND VPWR VPWR _1273_/X sky130_fd_sc_hd__a21o_1
X_0988_ hold24/X _0980_/X _0982_/Y _1009_/C VGND VGND VPWR VPWR _1620_/D sky130_fd_sc_hd__o211a_1
X_1609_ _1609_/CLK _1609_/D VGND VGND VPWR VPWR _1609_/Q sky130_fd_sc_hd__dfxtp_1
X_1444__80 _1454__90/A VGND VGND VPWR VPWR _1596_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0842_ _0956_/A _0842_/B VGND VGND VPWR VPWR _1658_/D sky130_fd_sc_hd__and2_1
X_0911_ _1346_/A _1076_/A VGND VGND VPWR VPWR _1201_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0773_ _1627_/Q VGND VGND VPWR VPWR _0773_/Y sky130_fd_sc_hd__inv_2
X_1325_ _1340_/A1 _1324_/X _1323_/X _1344_/C1 VGND VGND VPWR VPWR _1325_/X sky130_fd_sc_hd__a211o_1
X_1256_ hold49/A hold50/A hold43/A hold47/A _1547_/Q _1548_/Q VGND VGND VPWR VPWR
+ _1256_/X sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _1187_/A _1187_/B VGND VGND VPWR VPWR _1257_/B sky130_fd_sc_hd__or2_1
XFILLER_0_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1110_ hold43/X _1122_/B VGND VGND VPWR VPWR _1110_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1041_ hold5/X _1043_/A _1040_/Y VGND VGND VPWR VPWR _1601_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0825_ _0825_/A _0825_/B _0825_/C _0825_/D VGND VGND VPWR VPWR wire18/A sky130_fd_sc_hd__nor4_1
X_0756_ hold24/A VGND VGND VPWR VPWR _0817_/A sky130_fd_sc_hd__inv_2
XFILLER_0_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1308_ hold40/A _1342_/A2 _1333_/B1 _1307_/X VGND VGND VPWR VPWR _1308_/X sky130_fd_sc_hd__o211a_1
X_1239_ _1349_/A _1202_/A _1220_/Y _1221_/C VGND VGND VPWR VPWR _1239_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_34_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1414__50 clkload6/A VGND VGND VPWR VPWR _1566_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_30_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ _1590_/CLK _1590_/D VGND VGND VPWR VPWR _1590_/Q sky130_fd_sc_hd__dfxtp_1
X_1024_ hold28/A _1049_/A VGND VGND VPWR VPWR _1047_/A sky130_fd_sc_hd__and2_1
X_0808_ _1646_/Q _1608_/Q VGND VGND VPWR VPWR _0834_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload13/A sky130_fd_sc_hd__clkbuf_8
X_1642_ _1642_/CLK _1642_/D VGND VGND VPWR VPWR _1642_/Q sky130_fd_sc_hd__dfxtp_1
X_1573_ _1573_/CLK _1573_/D VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1007_ _1004_/B _1007_/B _1009_/C VGND VGND VPWR VPWR _1613_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1502__138 clkload2/A VGND VGND VPWR VPWR _1654_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_33_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1556_ _1556_/CLK _1556_/D VGND VGND VPWR VPWR uo_out[6] sky130_fd_sc_hd__dfxtp_4
X_1625_ _1625_/CLK _1625_/D VGND VGND VPWR VPWR _1625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1375__11 clkload13/A VGND VGND VPWR VPWR _1518_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1341_ _1517_/Q _1345_/A2 _1340_/X _1351_/A VGND VGND VPWR VPWR _1517_/D sky130_fd_sc_hd__o211a_1
X_1272_ _1516_/Q _1271_/X _1270_/X _1178_/S VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ _1621_/Q _0983_/B _0985_/B _1009_/C VGND VGND VPWR VPWR _1621_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1539_ _1541_/CLK input7/X VGND VGND VPWR VPWR _1539_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1608_ _1608_/CLK _1608_/D VGND VGND VPWR VPWR _1608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1467__103 clkload7/A VGND VGND VPWR VPWR _1619_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1508__144 clkload2/A VGND VGND VPWR VPWR _1660_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0772_ hold38/A VGND VGND VPWR VPWR _1257_/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ _0923_/A _1658_/Q _0836_/Y _0836_/A _1346_/A VGND VGND VPWR VPWR _0842_/B
+ sky130_fd_sc_hd__a32o_1
X_0910_ _0923_/A _0910_/B _0910_/C VGND VGND VPWR VPWR _0910_/X sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ _1548_/Q _1257_/B _1252_/X _1254_/X _1257_/A VGND VGND VPWR VPWR _1255_/X
+ sky130_fd_sc_hd__o311a_1
X_1324_ _1521_/Q _1519_/Q _1334_/S VGND VGND VPWR VPWR _1324_/X sky130_fd_sc_hd__mux2_1
X_1186_ _1187_/A _1187_/B VGND VGND VPWR VPWR _1186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1040_ hold5/X _1043_/A _1051_/B VGND VGND VPWR VPWR _1040_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0824_ _0830_/A _0832_/A _0824_/C _0824_/D VGND VGND VPWR VPWR _0825_/D sky130_fd_sc_hd__or4_1
X_0755_ hold36/A VGND VGND VPWR VPWR _0831_/A sky130_fd_sc_hd__inv_2
XFILLER_0_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1169_ _1080_/A _1178_/S _1179_/S VGND VGND VPWR VPWR _1169_/Y sky130_fd_sc_hd__o21ai_1
X_1238_ hold2/X _1130_/D _1237_/X _1259_/C1 VGND VGND VPWR VPWR _1544_/D sky130_fd_sc_hd__o211a_1
X_1307_ _1522_/Q _1322_/B VGND VGND VPWR VPWR _1307_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ hold15/A _1596_/Q hold7/A _1023_/D VGND VGND VPWR VPWR _1049_/A sky130_fd_sc_hd__and4_1
XFILLER_0_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0807_ _1611_/Q _0807_/B VGND VGND VPWR VPWR _0824_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
X_1572_ _1572_/CLK _1572_/D VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_1
X_1641_ _1641_/CLK _1641_/D VGND VGND VPWR VPWR _1641_/Q sky130_fd_sc_hd__dfxtp_1
X_1006_ _1613_/Q _1006_/B VGND VGND VPWR VPWR _1007_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1555_ _1555_/CLK _1555_/D VGND VGND VPWR VPWR uo_out[5] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1624_ _1624_/CLK _1624_/D VGND VGND VPWR VPWR _1624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_13_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1533_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_9_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1340_ _1340_/A1 _1339_/X _1338_/X _1344_/C1 VGND VGND VPWR VPWR _1340_/X sky130_fd_sc_hd__a211o_1
X_1390__26 clkload4/A VGND VGND VPWR VPWR _1542_/CLK sky130_fd_sc_hd__inv_2
X_1271_ _1349_/A _1349_/B _1530_/Q VGND VGND VPWR VPWR _1271_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire17 wire17/A VGND VGND VPWR VPWR wire17/X sky130_fd_sc_hd__buf_1
X_0986_ _1009_/C _0986_/B VGND VGND VPWR VPWR _1622_/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_14_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1538_ _1541_/CLK input6/X VGND VGND VPWR VPWR _1538_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1607_ _1607_/CLK _1607_/D VGND VGND VPWR VPWR _1607_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0771_ hold19/A VGND VGND VPWR VPWR _0771_/Y sky130_fd_sc_hd__inv_2
X_0840_ _0845_/A _0840_/B VGND VGND VPWR VPWR _1659_/D sky130_fd_sc_hd__and2_1
X_1435__71 clkload5/A VGND VGND VPWR VPWR _1587_/CLK sky130_fd_sc_hd__inv_2
X_1323_ _1521_/Q _0913_/Y _1333_/B1 _1322_/X VGND VGND VPWR VPWR _1323_/X sky130_fd_sc_hd__o211a_1
X_1254_ _1186_/Y _1253_/X _1548_/Q VGND VGND VPWR VPWR _1254_/X sky130_fd_sc_hd__a21bo_1
X_1185_ _1546_/Q hold54/A VGND VGND VPWR VPWR _1187_/B sky130_fd_sc_hd__nand2_1
X_0969_ _0971_/A _0969_/B VGND VGND VPWR VPWR _1624_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0754_ _1199_/A VGND VGND VPWR VPWR _1242_/A sky130_fd_sc_hd__inv_2
X_0823_ _0829_/C _0823_/B _0823_/C VGND VGND VPWR VPWR _0824_/D sky130_fd_sc_hd__or3_1
X_1306_ hold40/X _1275_/Y _1305_/X _1336_/C1 VGND VGND VPWR VPWR _1524_/D sky130_fd_sc_hd__o211a_1
X_1168_ _1157_/X _1166_/Y _1167_/X _1178_/S VGND VGND VPWR VPWR _1168_/X sky130_fd_sc_hd__o211a_1
X_1237_ _1358_/A _1203_/B _1221_/X _1236_/X VGND VGND VPWR VPWR _1237_/X sky130_fd_sc_hd__a31o_1
X_1099_ _1260_/A _1089_/X _1098_/X _0971_/A VGND VGND VPWR VPWR _1577_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1405__41 clkload6/A VGND VGND VPWR VPWR _1557_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ hold15/A _1596_/Q _1023_/D VGND VGND VPWR VPWR _1022_/X sky130_fd_sc_hd__and3_1
X_0806_ _1614_/Q _1652_/Q VGND VGND VPWR VPWR _0831_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
X_1640_ _1640_/CLK _1640_/D VGND VGND VPWR VPWR _1640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1571_ _1571_/CLK _1571_/D VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfxtp_1
X_1005_ _1002_/X _1005_/B _1009_/C VGND VGND VPWR VPWR _1614_/D sky130_fd_sc_hd__and3b_1
X_1396__32 clkload4/A VGND VGND VPWR VPWR _1548_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1554_ _1554_/CLK _1554_/D VGND VGND VPWR VPWR uo_out[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1623_ _1623_/CLK _1623_/D VGND VGND VPWR VPWR _1623_/Q sky130_fd_sc_hd__dfxtp_2
.ends

