* NGSPICE file created from tt_um_jimktrains_vslc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt tt_um_jimktrains_vslc VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_0_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1444__138 clkload0/A VGND VGND VPWR VPWR _1596_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1270_ _1459_/Q _1280_/B VGND VGND VPWR VPWR _1270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0985_ hold6/X _0987_/A _0984_/Y VGND VGND VPWR VPWR _1543_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1537_ _1537_/CLK _1537_/D VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
X_1468_ _1468_/CLK _1468_/D VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ _1550_/Q _1588_/Q VGND VGND VPWR VPWR _0770_/Y sky130_fd_sc_hd__nand2_1
X_1253_ _1283_/A1 _1252_/X _1251_/X _1287_/C1 VGND VGND VPWR VPWR _1253_/X sky130_fd_sc_hd__a211o_1
X_1184_ _1487_/Q _1131_/C _1123_/Y _1174_/X VGND VGND VPWR VPWR _1184_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0968_ hold17/A _0993_/A VGND VGND VPWR VPWR _0991_/A sky130_fd_sc_hd__and2_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload9/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0899_ _0802_/B _1571_/Q _0889_/Y _0889_/B _0734_/A VGND VGND VPWR VPWR _0900_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_25_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0822_ _0826_/A _0822_/B VGND VGND VPWR VPWR _1590_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ _1459_/Q _1458_/Q _1457_/Q _1471_/Q _1488_/Q _1489_/Q VGND VGND VPWR VPWR
+ _1306_/B sky130_fd_sc_hd__mux4_1
X_1236_ hold49/A _0864_/Y _1281_/B1 _1235_/X VGND VGND VPWR VPWR _1236_/X sky130_fd_sc_hd__o211a_1
X_1098_ _1075_/A _1096_/X _1098_/S VGND VGND VPWR VPWR _1098_/X sky130_fd_sc_hd__mux2_1
X_1167_ _1523_/Q _1109_/A _1165_/X _1166_/X VGND VGND VPWR VPWR _1182_/B sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_22_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1021_ _1289_/A _1138_/A _1020_/X _1145_/A VGND VGND VPWR VPWR _1529_/D sky130_fd_sc_hd__o211a_1
X_0805_ _0828_/A _0805_/B VGND VGND VPWR VPWR _1598_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0736_ _0736_/A VGND VGND VPWR VPWR _1069_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1219_ _0859_/B _1528_/Q _1007_/A VGND VGND VPWR VPWR _1219_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
X_1570_ _1570_/CLK _1570_/D VGND VGND VPWR VPWR _1570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1004_ hold29/A _1004_/B VGND VGND VPWR VPWR _1533_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1553_ _1553_/CLK _1553_/D VGND VGND VPWR VPWR _1553_/Q sky130_fd_sc_hd__dfxtp_1
X_1484_ _1484_/CLK _1484_/D VGND VGND VPWR VPWR _1484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_37_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1375__69 _1475_/CLK VGND VGND VPWR VPWR _1527_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ hold6/X _0987_/A _0983_/B VGND VGND VPWR VPWR _0984_/Y sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1536_ _1536_/CLK _1536_/D VGND VGND VPWR VPWR _1536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1467_ _1467_/CLK _1467_/D VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1411__105 clkload0/A VGND VGND VPWR VPWR _1563_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1252_ hold37/A _1463_/Q _1277_/S VGND VGND VPWR VPWR _1252_/X sky130_fd_sc_hd__mux2_1
X_1183_ _1072_/A _1182_/X _1168_/A VGND VGND VPWR VPWR _1183_/Y sky130_fd_sc_hd__a21boi_1
X_0967_ hold11/A _1538_/Q hold9/A _0967_/D VGND VGND VPWR VPWR _0993_/A sky130_fd_sc_hd__and4_1
X_0898_ _0915_/A _0898_/B VGND VGND VPWR VPWR _1572_/D sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1519_ _1519_/CLK _1519_/D VGND VGND VPWR VPWR _1519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1345__39 clkload8/A VGND VGND VPWR VPWR _1497_/CLK sky130_fd_sc_hd__inv_2
X_0752_ _1600_/Q VGND VGND VPWR VPWR _0752_/Y sky130_fd_sc_hd__inv_2
X_0821_ _0823_/A1 _1590_/Q _0813_/Y _0813_/B _1169_/A VGND VGND VPWR VPWR _0822_/B
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_24_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1304_ _1463_/Q _1462_/Q _1461_/Q hold54/A _1488_/Q _1489_/Q VGND VGND VPWR VPWR
+ _1304_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1166_ hold13/A hold24/A hold32/A hold22/A VGND VGND VPWR VPWR _1166_/X sky130_fd_sc_hd__or4_1
X_1235_ hold41/A _1275_/B VGND VGND VPWR VPWR _1235_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1097_ uo_out[5] _1097_/B VGND VGND VPWR VPWR _1097_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1417__111 clkload9/A VGND VGND VPWR VPWR _1569_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload8/A sky130_fd_sc_hd__clkbuf_8
X_1020_ _1020_/A _1030_/B VGND VGND VPWR VPWR _1020_/X sky130_fd_sc_hd__or2_1
X_0804_ _0823_/A1 _1598_/Q _0792_/Y _0792_/A _1169_/A VGND VGND VPWR VPWR _0805_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0735_ _1075_/A VGND VGND VPWR VPWR _1072_/A sky130_fd_sc_hd__inv_2
X_1149_ _1149_/A _1149_/B VGND VGND VPWR VPWR _1149_/Y sky130_fd_sc_hd__nor2_1
X_1218_ _0859_/B _1528_/Q _1007_/A VGND VGND VPWR VPWR _1218_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1003_ hold29/X _1534_/Q _1002_/Y VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1552_ _1552_/CLK _1552_/D VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfxtp_2
X_1483_ _1483_/CLK input9/X VGND VGND VPWR VPWR _1483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ _0972_/B _0983_/B _0983_/C VGND VGND VPWR VPWR _1544_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1535_ _1535_/CLK _1535_/D VGND VGND VPWR VPWR _1535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1466_ _1466_/CLK _1466_/D VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1450__144 _1450__144/A VGND VGND VPWR VPWR _1602_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1251_ hold37/A _1285_/A2 _1285_/C1 _1250_/X VGND VGND VPWR VPWR _1251_/X sky130_fd_sc_hd__o211a_1
X_1182_ _1182_/A _1182_/B _1182_/C VGND VGND VPWR VPWR _1182_/X sky130_fd_sc_hd__and3_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0966_ hold11/A _1538_/Q _0967_/D VGND VGND VPWR VPWR _0966_/X sky130_fd_sc_hd__and3_1
X_0897_ _0802_/B _1572_/Q _0889_/Y _0889_/B _1291_/D VGND VGND VPWR VPWR _0898_/B
+ sky130_fd_sc_hd__a32o_1
X_1434__128 clkload2/A VGND VGND VPWR VPWR _1586_/CLK sky130_fd_sc_hd__inv_2
X_1518_ _1518_/CLK _1518_/D VGND VGND VPWR VPWR _1518_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0751_ _1597_/Q VGND VGND VPWR VPWR _0751_/Y sky130_fd_sc_hd__inv_2
X_0820_ hold31/X _0801_/X _0813_/Y _0813_/B _0800_/A VGND VGND VPWR VPWR _1591_/D
+ sky130_fd_sc_hd__a32o_1
X_1303_ _1292_/B _1301_/Y _1302_/X _1303_/C1 VGND VGND VPWR VPWR _1452_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1096_ _1292_/B uo_out[5] _1096_/S VGND VGND VPWR VPWR _1096_/X sky130_fd_sc_hd__mux2_1
X_1165_ hold19/A hold33/A _1496_/Q hold36/A VGND VGND VPWR VPWR _1165_/X sky130_fd_sc_hd__or4_1
XFILLER_0_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1234_ hold49/X _1288_/A2 _1233_/X _1284_/C1 VGND VGND VPWR VPWR _1468_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_22_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0949_ _0946_/X _0949_/B _0963_/B VGND VGND VPWR VPWR _1556_/D sky130_fd_sc_hd__and3b_1
X_1405__99 clkload1/A VGND VGND VPWR VPWR _1557_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0734_ _0734_/A VGND VGND VPWR VPWR _1024_/A sky130_fd_sc_hd__inv_2
X_0803_ hold18/X _0792_/Y _0801_/X _0800_/A _0792_/A VGND VGND VPWR VPWR _1599_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1079_ _1074_/X _1076_/X _1078_/X _1169_/B VGND VGND VPWR VPWR _1207_/B sky130_fd_sc_hd__o22ai_1
X_1217_ _1471_/Q _1005_/Y _1214_/X _1216_/X _1294_/A VGND VGND VPWR VPWR _1471_/D
+ sky130_fd_sc_hd__o221a_1
X_1148_ hold47/A hold50/A hold52/A hold46/A VGND VGND VPWR VPWR _1149_/B sky130_fd_sc_hd__or4_1
XFILLER_0_30_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ hold29/A _1534_/Q _1004_/B VGND VGND VPWR VPWR _1002_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload7/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1482_ _1483_/CLK input8/X VGND VGND VPWR VPWR _1482_/Q sky130_fd_sc_hd__dfxtp_1
X_1551_ _1551_/CLK _1551_/D VGND VGND VPWR VPWR _1551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0982_ hold23/A hold6/A _0989_/A _1544_/Q VGND VGND VPWR VPWR _0983_/C sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_14_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1465_ _1465_/CLK _1465_/D VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1534_ _1534_/CLK hold30/X VGND VGND VPWR VPWR _1534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1380__74 clkload9/A VGND VGND VPWR VPWR _1532_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1250_ _1463_/Q _1280_/B VGND VGND VPWR VPWR _1250_/X sky130_fd_sc_hd__or2_1
X_1181_ hold38/X _1126_/B _1180_/X _1196_/A VGND VGND VPWR VPWR _1485_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0965_ hold29/A _1534_/Q _1535_/Q _1536_/Q VGND VGND VPWR VPWR _0967_/D sky130_fd_sc_hd__and4_1
X_0896_ hold15/X _0801_/X _0889_/Y _0889_/B _0800_/A VGND VGND VPWR VPWR _1573_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1517_ _1517_/CLK _1517_/D VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0750_ _1593_/Q VGND VGND VPWR VPWR _0750_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1302_ _1301_/A _1301_/B uo_out[0] VGND VGND VPWR VPWR _1302_/X sky130_fd_sc_hd__a21o_1
X_1233_ _1283_/A1 _1232_/X _1231_/X _1287_/C1 VGND VGND VPWR VPWR _1233_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1095_ _1169_/B _1298_/A VGND VGND VPWR VPWR _1096_/S sky130_fd_sc_hd__nand2_1
X_1164_ _1523_/Q _1109_/A _1153_/Y _1162_/X _1163_/X VGND VGND VPWR VPWR _1182_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0948_ _1556_/Q _0951_/A VGND VGND VPWR VPWR _0949_/B sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0879_ _0903_/A1 _1580_/Q _0871_/Y _0871_/B _1291_/D VGND VGND VPWR VPWR _0880_/B
+ sky130_fd_sc_hd__a32o_1
X_1350__44 clkload11/A VGND VGND VPWR VPWR _1502_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0802_ _0915_/A _0802_/B VGND VGND VPWR VPWR _0974_/B sky130_fd_sc_hd__nand2_1
X_0733_ _1553_/Q VGND VGND VPWR VPWR _0733_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1216_ _1285_/C1 _1215_/X _1007_/A VGND VGND VPWR VPWR _1216_/X sky130_fd_sc_hd__a21o_1
X_1078_ uo_out[3] _1069_/Y _1295_/A uo_out[2] _1077_/X VGND VGND VPWR VPWR _1078_/X
+ sky130_fd_sc_hd__a221o_1
X_1147_ _1511_/Q hold45/A hold53/A hold44/A VGND VGND VPWR VPWR _1149_/A sky130_fd_sc_hd__or4_1
XFILLER_0_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1001_ _1001_/A _1004_/B _1001_/C VGND VGND VPWR VPWR _1535_/D sky130_fd_sc_hd__and3_1
XFILLER_0_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320__14 _1483_/CLK VGND VGND VPWR VPWR _1463_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1407__101 clkload0/A VGND VGND VPWR VPWR _1559_/CLK sky130_fd_sc_hd__inv_2
X_1481_ _1483_/CLK input7/X VGND VGND VPWR VPWR _1481_/Q sky130_fd_sc_hd__dfxtp_1
X_1550_ _1550_/CLK _1550_/D VGND VGND VPWR VPWR _1550_/Q sky130_fd_sc_hd__dfxtp_1
X_1386__80 clkload7/A VGND VGND VPWR VPWR _1538_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ _0981_/A _0981_/B VGND VGND VPWR VPWR _1545_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1602_ _1602_/CLK _1602_/D VGND VGND VPWR VPWR _1602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1464_ _1464_/CLK _1464_/D VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1533_ _1533_/CLK _1533_/D VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1356__50 _1359__53/A VGND VGND VPWR VPWR _1508_/CLK sky130_fd_sc_hd__inv_2
X_1180_ _1301_/A _1168_/X _1182_/C _1179_/X VGND VGND VPWR VPWR _1180_/X sky130_fd_sc_hd__a31o_1
X_0964_ hold29/A _1534_/Q _1535_/Q VGND VGND VPWR VPWR _1001_/A sky130_fd_sc_hd__nand3_1
X_0895_ _1022_/A _0895_/B VGND VGND VPWR VPWR _1574_/D sky130_fd_sc_hd__and2_1
X_1516_ _1516_/CLK _1516_/D VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1301_ _1301_/A _1301_/B VGND VGND VPWR VPWR _1301_/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1232_ hold39/A hold42/A _1277_/S VGND VGND VPWR VPWR _1232_/X sky130_fd_sc_hd__mux2_1
X_1094_ uo_out[6] _1097_/B _1092_/X _1093_/X _1145_/A VGND VGND VPWR VPWR _1505_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ hold24/A hold51/A VGND VGND VPWR VPWR _1163_/X sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_30_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ _1557_/Q _0946_/X _0963_/B _0920_/Y VGND VGND VPWR VPWR _1557_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1440__134 _1450__144/A VGND VGND VPWR VPWR _1592_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ hold16/X _0801_/X _0871_/Y _0871_/B _0800_/A VGND VGND VPWR VPWR _1581_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload0 clkload0/A VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_2
X_1326__20 clkload11/A VGND VGND VPWR VPWR _1469_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_28_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1424__118 clkload6/A VGND VGND VPWR VPWR _1576_/CLK sky130_fd_sc_hd__inv_2
X_0801_ _0904_/A _1196_/B VGND VGND VPWR VPWR _0801_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0732_ _1556_/Q VGND VGND VPWR VPWR _0732_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1146_ _1488_/Q _1139_/B _1145_/Y VGND VGND VPWR VPWR _1488_/D sky130_fd_sc_hd__a21o_1
X_1215_ _1291_/D _0734_/A _1075_/A _1075_/B _1471_/Q _1457_/Q VGND VGND VPWR VPWR
+ _1215_/X sky130_fd_sc_hd__mux4_1
X_1077_ uo_out[1] _1298_/A _1301_/A uo_out[0] VGND VGND VPWR VPWR _1077_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1000_ hold29/A _1534_/Q _1535_/Q VGND VGND VPWR VPWR _1001_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1446__140 clkload0/A VGND VGND VPWR VPWR _1598_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1129_ hold38/X _1492_/Q _1130_/S VGND VGND VPWR VPWR _1492_/D sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ _1483_/CLK input6/X VGND VGND VPWR VPWR _1480_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ hold26/X _0972_/B _0983_/B VGND VGND VPWR VPWR _0981_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1601_ _1601_/CLK _1601_/D VGND VGND VPWR VPWR _1601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1532_ _1532_/CLK _1532_/D VGND VGND VPWR VPWR _1532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1463_ _1463_/CLK _1463_/D VGND VGND VPWR VPWR _1463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1371__65 clkload9/A VGND VGND VPWR VPWR _1523_/CLK sky130_fd_sc_hd__inv_2
X_0963_ _0960_/B _0963_/B _0963_/C VGND VGND VPWR VPWR _1549_/D sky130_fd_sc_hd__and3b_1
X_0894_ _0903_/A1 _1574_/Q _0889_/Y _0889_/B _1289_/A VGND VGND VPWR VPWR _0895_/B
+ sky130_fd_sc_hd__a32o_1
X_1515_ _1515_/CLK _1515_/D VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1300_ _1292_/B _1298_/Y _1299_/X _1303_/C1 VGND VGND VPWR VPWR _1453_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1162_ _1521_/Q _1112_/A _1160_/X _1161_/X VGND VGND VPWR VPWR _1162_/X sky130_fd_sc_hd__a22o_1
X_1231_ hold39/A _0864_/Y _1281_/B1 _1230_/X VGND VGND VPWR VPWR _1231_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1093_ _1169_/B _1285_/C1 _1087_/Y VGND VGND VPWR VPWR _1093_/X sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_22_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0946_ _1556_/Q _1555_/Q _0946_/C VGND VGND VPWR VPWR _0946_/X sky130_fd_sc_hd__and3_1
X_0877_ _0904_/A _0877_/B VGND VGND VPWR VPWR _1582_/D sky130_fd_sc_hd__and2_1
Xclkload1 clkload1/A VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_4
XFILLER_0_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1341__35 clkload3/A VGND VGND VPWR VPWR _1493_/CLK sky130_fd_sc_hd__inv_2
X_0731_ _1557_/Q VGND VGND VPWR VPWR _0731_/Y sky130_fd_sc_hd__inv_2
X_0800_ _0800_/A VGND VGND VPWR VPWR _1289_/B sky130_fd_sc_hd__inv_2
X_1145_ _1145_/A _1145_/B VGND VGND VPWR VPWR _1145_/Y sky130_fd_sc_hd__nand2_1
X_1214_ _1457_/Q _1282_/S _1098_/S _1213_/X VGND VGND VPWR VPWR _1214_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1076_ uo_out[6] _1295_/A _1301_/A uo_out[4] _1024_/A VGND VGND VPWR VPWR _1076_/X
+ sky130_fd_sc_hd__a221o_1
X_0929_ _1564_/Q _0931_/B VGND VGND VPWR VPWR _0932_/A sky130_fd_sc_hd__or2_1
XFILLER_0_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1128_ _1486_/Q hold3/X _1130_/S VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1059_ _1020_/A _1051_/X _1058_/X _1126_/A VGND VGND VPWR VPWR _1512_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1377__71 clkload4/A VGND VGND VPWR VPWR _1529_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1462_ _1462_/CLK _1462_/D VGND VGND VPWR VPWR _1462_/Q sky130_fd_sc_hd__dfxtp_1
X_1531_ _1531_/CLK _1531_/D VGND VGND VPWR VPWR _1531_/Q sky130_fd_sc_hd__dfxtp_1
X_1600_ _1600_/CLK _1600_/D VGND VGND VPWR VPWR _1600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0962_ _1549_/Q _0974_/A VGND VGND VPWR VPWR _0963_/C sky130_fd_sc_hd__or2_1
X_0893_ _0915_/A _0893_/B VGND VGND VPWR VPWR _1575_/D sky130_fd_sc_hd__and2_1
X_1514_ _1514_/CLK _1514_/D VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfxtp_1
X_1347__41 clkload11/A VGND VGND VPWR VPWR _1499_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1309__3 _1475_/CLK VGND VGND VPWR VPWR _1452_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout60 input1/X VGND VGND VPWR VPWR _1303_/C1 sky130_fd_sc_hd__clkbuf_2
X_1092_ _1292_/B _1090_/Y _1091_/X _1098_/S VGND VGND VPWR VPWR _1092_/X sky130_fd_sc_hd__o211a_1
X_1230_ hold42/A _1280_/B VGND VGND VPWR VPWR _1230_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1161_ _1521_/Q _1112_/A _0739_/Y _1520_/Q VGND VGND VPWR VPWR _1161_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_35_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0945_ _1555_/Q _0946_/C VGND VGND VPWR VPWR _0951_/A sky130_fd_sc_hd__and2_1
X_0876_ _0903_/A1 _1582_/Q _0871_/Y _0871_/B _1289_/A VGND VGND VPWR VPWR _0877_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload2 clkload2/A VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_6
X_0730_ _1558_/Q VGND VGND VPWR VPWR _0730_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1317__11 _1483_/CLK VGND VGND VPWR VPWR _1460_/CLK sky130_fd_sc_hd__inv_2
X_1213_ _1207_/Y _1210_/X _1212_/X _1291_/C VGND VGND VPWR VPWR _1213_/X sky130_fd_sc_hd__a31o_1
X_1144_ _1144_/A _1144_/B VGND VGND VPWR VPWR _1489_/D sky130_fd_sc_hd__nand2_1
X_1075_ _1075_/A _1075_/B VGND VGND VPWR VPWR _1301_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ _1563_/Q _1562_/Q _0928_/C VGND VGND VPWR VPWR _0931_/B sky130_fd_sc_hd__and3_1
X_0859_ _1071_/A _0859_/B _0906_/C VGND VGND VPWR VPWR _0859_/X sky130_fd_sc_hd__or3_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
X_1401__95 clkload1/A VGND VGND VPWR VPWR _1553_/CLK sky130_fd_sc_hd__inv_2
X_1430__124 clkload2/A VGND VGND VPWR VPWR _1582_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_32_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1127_ _1178_/A hold7/X _1130_/S VGND VGND VPWR VPWR _1494_/D sky130_fd_sc_hd__mux2_1
X_1058_ hold46/X _1066_/B VGND VGND VPWR VPWR _1058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1414__108 clkload7/A VGND VGND VPWR VPWR _1566_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1392__86 clkload7/A VGND VGND VPWR VPWR _1544_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1461_ _1461_/CLK _1461_/D VGND VGND VPWR VPWR _1461_/Q sky130_fd_sc_hd__dfxtp_1
X_1436__130 _1450__144/A VGND VGND VPWR VPWR _1588_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1530_ _1530_/CLK _1530_/D VGND VGND VPWR VPWR _1530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0961_ _0958_/B _0961_/B _0963_/B VGND VGND VPWR VPWR _1550_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0892_ _0802_/B _1575_/Q _0889_/Y _0889_/B _1071_/A VGND VGND VPWR VPWR _0893_/B
+ sky130_fd_sc_hd__a32o_1
X_1513_ _1513_/CLK _1513_/D VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfxtp_1
X_1362__56 clkload3/A VGND VGND VPWR VPWR _1514_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_10_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout50 _0904_/A VGND VGND VPWR VPWR _0828_/A sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1091_ _1169_/B _1295_/A uo_out[6] VGND VGND VPWR VPWR _1091_/X sky130_fd_sc_hd__a21o_1
X_1160_ _1157_/X _1158_/X _1159_/X VGND VGND VPWR VPWR _1160_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_27_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0944_ _1554_/Q _0960_/B _0944_/C VGND VGND VPWR VPWR _0946_/C sky130_fd_sc_hd__and3_1
XFILLER_0_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0875_ _0904_/A _0875_/B VGND VGND VPWR VPWR _1583_/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1311__5 clkload5/A VGND VGND VPWR VPWR _1454_/CLK sky130_fd_sc_hd__inv_2
X_1289_ _1289_/A _1289_/B _1289_/C _1289_/D VGND VGND VPWR VPWR _1290_/S sky130_fd_sc_hd__or4_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload3 clkload3/A VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_21_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1212_ _1477_/Q _1298_/A _1206_/X _1211_/X VGND VGND VPWR VPWR _1212_/X sky130_fd_sc_hd__a211o_1
X_1332__26 clkload4/A VGND VGND VPWR VPWR _1484_/CLK sky130_fd_sc_hd__inv_2
X_1143_ _1489_/Q _1145_/B _1068_/A VGND VGND VPWR VPWR _1144_/B sky130_fd_sc_hd__a21oi_1
X_1074_ uo_out[7] _1069_/Y _1298_/A uo_out[5] VGND VGND VPWR VPWR _1074_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ _1562_/Q _0928_/C VGND VGND VPWR VPWR _0927_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0789_ hold21/A _0789_/B _0789_/C _0789_/D VGND VGND VPWR VPWR _0789_/X sky130_fd_sc_hd__and4_1
X_0858_ _1071_/A _1082_/B _0906_/C VGND VGND VPWR VPWR _1291_/C sky130_fd_sc_hd__nor3_2
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_1398__92 _1400__94/A VGND VGND VPWR VPWR _1550_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1126_ _1126_/A _1126_/B VGND VGND VPWR VPWR _1130_/S sky130_fd_sc_hd__nand2_1
X_1057_ _0864_/B _1051_/X _1056_/X _1126_/A VGND VGND VPWR VPWR _1513_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _1109_/A _1111_/A VGND VGND VPWR VPWR _1502_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1368__62 clkload9/A VGND VGND VPWR VPWR _1520_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ _1460_/CLK _1460_/D VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1589_ _1589_/CLK _1589_/D VGND VGND VPWR VPWR _1589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ _1550_/Q _0960_/B VGND VGND VPWR VPWR _0961_/B sky130_fd_sc_hd__or2_1
X_0891_ _0915_/A _0891_/B VGND VGND VPWR VPWR _1576_/D sky130_fd_sc_hd__and2_1
X_1512_ _1512_/CLK _1512_/D VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1338__32 _1359__53/A VGND VGND VPWR VPWR _1490_/CLK sky130_fd_sc_hd__inv_2
Xfanout40 _1169_/A VGND VGND VPWR VPWR _1207_/A sky130_fd_sc_hd__clkbuf_2
Xfanout51 _1196_/A VGND VGND VPWR VPWR _0904_/A sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ _1169_/B _1295_/A VGND VGND VPWR VPWR _1090_/Y sky130_fd_sc_hd__nand2_1
Xclkload10 _1475_/CLK VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0943_ _0960_/B _0944_/C VGND VGND VPWR VPWR _0952_/B sky130_fd_sc_hd__and2_1
X_0874_ _0903_/A1 _1583_/Q _0871_/Y _0871_/B _1016_/A VGND VGND VPWR VPWR _0875_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_38_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1288_ _1457_/Q _1288_/A2 _1287_/X _1294_/A VGND VGND VPWR VPWR _1457_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_21_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload4 clkload4/A VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_6
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ _1478_/Q _1295_/A _1207_/A _1169_/B VGND VGND VPWR VPWR _1211_/X sky130_fd_sc_hd__a211o_1
X_1142_ _1490_/Q _1144_/A _1141_/Y VGND VGND VPWR VPWR _1490_/D sky130_fd_sc_hd__a21o_1
X_1073_ _1075_/A _1075_/B VGND VGND VPWR VPWR _1298_/A sky130_fd_sc_hd__and2b_2
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ _0928_/C VGND VGND VPWR VPWR _0926_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ _1289_/A _1020_/A VGND VGND VPWR VPWR _0906_/C sky130_fd_sc_hd__nor2_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ _1553_/Q _0749_/Y _0751_/Y _1559_/Q _0773_/X VGND VGND VPWR VPWR _0790_/C
+ sky130_fd_sc_hd__a221o_1
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1125_ _1126_/B VGND VGND VPWR VPWR _1125_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ hold52/X _1066_/B VGND VGND VPWR VPWR _1056_/X sky130_fd_sc_hd__or2_1
X_0909_ _0915_/A _0909_/B VGND VGND VPWR VPWR _1568_/D sky130_fd_sc_hd__and2_1
XFILLER_0_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1039_ _1289_/A _1033_/X _1038_/X _1022_/A VGND VGND VPWR VPWR _1521_/D sky130_fd_sc_hd__o211a_1
X_1108_ hold24/A hold32/A _1114_/A VGND VGND VPWR VPWR _1111_/A sky130_fd_sc_hd__and3_1
X_1420__114 _1400__94/A VGND VGND VPWR VPWR _1572_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1383__77 clkload8/A VGND VGND VPWR VPWR _1535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1588_ _1588_/CLK _1588_/D VGND VGND VPWR VPWR _1588_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0802_/B _1576_/Q _0889_/Y _0889_/B _0859_/B VGND VGND VPWR VPWR _0891_/B
+ sky130_fd_sc_hd__a32o_1
X_1511_ _1511_/CLK _1511_/D VGND VGND VPWR VPWR _1511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1353__47 clkload5/A VGND VGND VPWR VPWR _1505_/CLK sky130_fd_sc_hd__inv_2
Xfanout52 _1145_/A VGND VGND VPWR VPWR _1126_/A sky130_fd_sc_hd__buf_2
Xfanout41 _1527_/Q VGND VGND VPWR VPWR _1169_/A sky130_fd_sc_hd__clkbuf_4
X_1426__120 _1400__94/A VGND VGND VPWR VPWR _1578_/CLK sky130_fd_sc_hd__inv_2
Xfanout30 _1585_/Q VGND VGND VPWR VPWR _0903_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload11 clkload11/A VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_4
X_0942_ _1551_/Q _1550_/Q _0960_/B VGND VGND VPWR VPWR _0942_/X sky130_fd_sc_hd__and3_1
X_0873_ _0904_/A _0873_/B VGND VGND VPWR VPWR _1584_/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ _1098_/S _1286_/X _1285_/X _1287_/C1 VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__a211o_1
Xclkload5 clkload5/A VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1141_ _1490_/Q _1144_/A _1145_/A VGND VGND VPWR VPWR _1141_/Y sky130_fd_sc_hd__o21ai_1
X_1210_ _1483_/Q _1069_/Y _1208_/X _1209_/X VGND VGND VPWR VPWR _1210_/X sky130_fd_sc_hd__a211o_1
X_1072_ _1072_/A _1075_/B VGND VGND VPWR VPWR _1295_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0856_ _1071_/A _1082_/B _1471_/Q _1289_/A VGND VGND VPWR VPWR _0856_/X sky130_fd_sc_hd__or4b_1
X_0925_ hold40/A _1560_/Q _1559_/Q _0925_/D VGND VGND VPWR VPWR _0928_/C sky130_fd_sc_hd__and4_1
X_0787_ _0769_/X _0770_/Y _0771_/X _0772_/Y _0768_/X VGND VGND VPWR VPWR _0790_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_1323__17 clkload11/A VGND VGND VPWR VPWR _1466_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1389__83 clkload7/A VGND VGND VPWR VPWR _1541_/CLK sky130_fd_sc_hd__inv_2
X_1124_ _1490_/Q _1489_/Q _1488_/Q _1123_/A VGND VGND VPWR VPWR _1126_/B sky130_fd_sc_hd__o31ai_4
X_1055_ _1530_/Q _1051_/X _1054_/X _1126_/A VGND VGND VPWR VPWR _1514_/D sky130_fd_sc_hd__o211a_1
X_0908_ _0802_/B _1568_/Q _0907_/Y _0907_/B _1291_/D VGND VGND VPWR VPWR _0909_/B
+ sky130_fd_sc_hd__a32o_1
X_0839_ _0732_/Y _1576_/Q _1550_/Q _0744_/Y VGND VGND VPWR VPWR _0841_/C sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_17_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ hold22/A _1116_/A VGND VGND VPWR VPWR _1114_/A sky130_fd_sc_hd__and2_1
X_1038_ _1521_/Q _1048_/B VGND VGND VPWR VPWR _1038_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1359__53 _1359__53/A VGND VGND VPWR VPWR _1511_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1443__137 clkload0/A VGND VGND VPWR VPWR _1595_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1587_ _1587_/CLK _1587_/D VGND VGND VPWR VPWR _1587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1510_ _1510_/CLK _1510_/D VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout53 _1196_/A VGND VGND VPWR VPWR _1145_/A sky130_fd_sc_hd__buf_2
Xfanout31 _1053_/A1 VGND VGND VPWR VPWR _1082_/B sky130_fd_sc_hd__buf_2
Xfanout42 _0734_/A VGND VGND VPWR VPWR _1169_/B sky130_fd_sc_hd__clkbuf_4
Xfanout20 _0859_/X VGND VGND VPWR VPWR _1282_/S sky130_fd_sc_hd__clkbuf_2
X_1329__23 _1359__53/A VGND VGND VPWR VPWR _1472_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0941_ _1550_/Q _0960_/B VGND VGND VPWR VPWR _0958_/B sky130_fd_sc_hd__and2_1
Xclkload12 _1483_/CLK VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_6
XFILLER_0_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0872_ _1196_/B _1584_/Q _0871_/Y _0871_/B _1053_/A1 VGND VGND VPWR VPWR _0873_/B
+ sky130_fd_sc_hd__a32o_1
X_1286_ _1471_/Q _1458_/Q _1291_/C VGND VGND VPWR VPWR _1286_/X sky130_fd_sc_hd__mux2_1
X_1449__143 _1450__144/A VGND VGND VPWR VPWR _1601_/CLK sky130_fd_sc_hd__inv_2
Xclkload6 clkload6/A VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_4
XFILLER_0_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ _1489_/Q _1145_/B VGND VGND VPWR VPWR _1144_/A sky130_fd_sc_hd__or2_1
X_1071_ _1071_/A _1082_/B _0864_/B _1020_/A VGND VGND VPWR VPWR _1071_/X sky130_fd_sc_hd__or4bb_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ _0937_/A _0937_/B VGND VGND VPWR VPWR _0924_/Y sky130_fd_sc_hd__nor2_1
X_0786_ _1555_/Q _0750_/Y _0778_/X _0784_/X _0785_/Y VGND VGND VPWR VPWR _0790_/A
+ sky130_fd_sc_hd__a2111o_1
X_0855_ _0888_/A _1492_/Q hold48/A VGND VGND VPWR VPWR _1289_/C sky130_fd_sc_hd__or3b_4
XFILLER_0_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ _1461_/Q _1288_/A2 _1268_/X _1303_/C1 VGND VGND VPWR VPWR _1461_/D sky130_fd_sc_hd__o211a_1
X_1123_ _1123_/A VGND VGND VPWR VPWR _1123_/Y sky130_fd_sc_hd__inv_2
X_1054_ hold50/X _1066_/B VGND VGND VPWR VPWR _1054_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0907_ _0907_/A _0907_/B VGND VGND VPWR VPWR _0907_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0769_ _1550_/Q _1588_/Q VGND VGND VPWR VPWR _0769_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0838_ _1549_/Q _0743_/Y _0745_/Y _1551_/Q VGND VGND VPWR VPWR _0841_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1106_ hold19/A hold33/A _1117_/B VGND VGND VPWR VPWR _1116_/A sky130_fd_sc_hd__and3_1
XFILLER_0_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1037_ _1071_/A _1033_/X _1036_/X _1022_/A VGND VGND VPWR VPWR _1522_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1374__68 clkload4/A VGND VGND VPWR VPWR _1526_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1586_ _1586_/CLK _1586_/D VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
X_1314__8 _1475_/CLK VGND VGND VPWR VPWR _1457_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410__104 clkload0/A VGND VGND VPWR VPWR _1562_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1569_ _1569_/CLK _1569_/D VGND VGND VPWR VPWR _1569_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout21 _1098_/S VGND VGND VPWR VPWR _1283_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout54 input1/X VGND VGND VPWR VPWR _1196_/A sky130_fd_sc_hd__clkbuf_2
Xfanout32 _1053_/A1 VGND VGND VPWR VPWR _0859_/B sky130_fd_sc_hd__clkbuf_2
Xfanout43 _1063_/A1 VGND VGND VPWR VPWR _0734_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1344__38 clkload8/A VGND VGND VPWR VPWR _1496_/CLK sky130_fd_sc_hd__inv_2
X_0940_ _1558_/Q _0920_/A _0922_/Y _0959_/C VGND VGND VPWR VPWR _1558_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0871_ _0907_/A _0871_/B VGND VGND VPWR VPWR _0871_/Y sky130_fd_sc_hd__nor2_2
X_1285_ _1458_/Q _1285_/A2 _0867_/C _1285_/C1 VGND VGND VPWR VPWR _1285_/X sky130_fd_sc_hd__o211a_1
Xclkload7 clkload7/A VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _1075_/A _1075_/B VGND VGND VPWR VPWR _1292_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0923_ _1559_/Q _0925_/D VGND VGND VPWR VPWR _0937_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0854_ _0854_/A hold7/A hold3/A VGND VGND VPWR VPWR _0888_/A sky130_fd_sc_hd__or3b_4
X_1416__110 _1400__94/A VGND VGND VPWR VPWR _1568_/CLK sky130_fd_sc_hd__inv_2
X_0785_ _0730_/Y _1596_/Q _0767_/Y _0776_/Y _0777_/Y VGND VGND VPWR VPWR _0785_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1268_ _1098_/S _1267_/X _1266_/X _1219_/X VGND VGND VPWR VPWR _1268_/X sky130_fd_sc_hd__a211o_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_1199_ _1490_/Q _1201_/A _1199_/C VGND VGND VPWR VPWR _1199_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_14_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ _1178_/A _1486_/Q _1122_/C VGND VGND VPWR VPWR _1123_/A sky130_fd_sc_hd__or3_2
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1053_ _1053_/A1 _1051_/X _1052_/X _1126_/A VGND VGND VPWR VPWR _1515_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_3_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0837_ _0729_/Y _1579_/Q _1580_/Q _0937_/A _0831_/X VGND VGND VPWR VPWR _0841_/A
+ sky130_fd_sc_hd__a221o_1
X_0906_ _1082_/B _1289_/C _0906_/C _1071_/A VGND VGND VPWR VPWR _0907_/B sky130_fd_sc_hd__and4bb_2
X_0768_ hold10/A _1590_/Q VGND VGND VPWR VPWR _0768_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ _1105_/A _1496_/Q hold36/A _1105_/D VGND VGND VPWR VPWR _1117_/B sky130_fd_sc_hd__and4_1
XFILLER_0_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1036_ hold51/X _1048_/B VGND VGND VPWR VPWR _1036_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1585_ _1585_/CLK _1585_/D VGND VGND VPWR VPWR _1585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _1016_/A _1138_/A _1018_/X _1294_/A VGND VGND VPWR VPWR _1530_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1568_ _1568_/CLK _1568_/D VGND VGND VPWR VPWR _1568_/Q sky130_fd_sc_hd__dfxtp_1
X_1499_ _1499_/CLK _1499_/D VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dfxtp_1
Xfanout22 _1082_/Y VGND VGND VPWR VPWR _1098_/S sky130_fd_sc_hd__clkbuf_4
Xfanout33 _1531_/Q VGND VGND VPWR VPWR _1053_/A1 sky130_fd_sc_hd__buf_2
Xfanout11 _0930_/Y VGND VGND VPWR VPWR _0959_/C sky130_fd_sc_hd__buf_2
Xfanout55 _1105_/A VGND VGND VPWR VPWR _0915_/A sky130_fd_sc_hd__clkbuf_2
Xfanout44 _1526_/Q VGND VGND VPWR VPWR _1063_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1433__127 clkload9/A VGND VGND VPWR VPWR _1585_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ _0888_/A _1033_/B VGND VGND VPWR VPWR _0871_/B sky130_fd_sc_hd__nor2_4
X_1284_ _1458_/Q _1288_/A2 _1283_/X _1284_/C1 VGND VGND VPWR VPWR _1458_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0999_ _0967_/D _1004_/B _0999_/C VGND VGND VPWR VPWR _1536_/D sky130_fd_sc_hd__and3b_1
Xclkload8 clkload8/A VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1404__98 clkload1/A VGND VGND VPWR VPWR _1556_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0753__1 clkload5/A VGND VGND VPWR VPWR _1451_/CLK sky130_fd_sc_hd__inv_2
X_0922_ _0925_/D VGND VGND VPWR VPWR _0922_/Y sky130_fd_sc_hd__inv_2
X_0853_ hold21/X _0930_/B _0852_/Y VGND VGND VPWR VPWR _1586_/D sky130_fd_sc_hd__o21a_1
X_0784_ _1549_/Q _0747_/Y _0765_/X _0774_/X _0775_/X VGND VGND VPWR VPWR _0784_/X
+ sky130_fd_sc_hd__a2111o_1
Xinput1 rst_n VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1267_ _1462_/Q hold54/A _1277_/S VGND VGND VPWR VPWR _1267_/X sky130_fd_sc_hd__mux2_1
X_1198_ hold46/A hold52/A hold50/A hold47/A _1488_/Q _1489_/Q VGND VGND VPWR VPWR
+ _1199_/C sky130_fd_sc_hd__mux4_1
XFILLER_0_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1439__133 _1450__144/A VGND VGND VPWR VPWR _1591_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_27_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ _1484_/Q hold38/A VGND VGND VPWR VPWR _1122_/C sky130_fd_sc_hd__and2b_1
X_1052_ hold47/X _1066_/B VGND VGND VPWR VPWR _1052_/X sky130_fd_sc_hd__or2_1
X_0767_ _1554_/Q _1592_/Q VGND VGND VPWR VPWR _0767_/Y sky130_fd_sc_hd__nand2b_1
X_0836_ _0733_/Y hold15/A _0829_/Y _0835_/X hold21/A VGND VGND VPWR VPWR _0850_/A
+ sky130_fd_sc_hd__a2111o_1
X_0905_ _1082_/B _1016_/A VGND VGND VPWR VPWR _1289_/D sky130_fd_sc_hd__nand2b_1
X_1395__89 _1400__94/A VGND VGND VPWR VPWR _1547_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1104_ uo_out[4] _1097_/B _1103_/X _1145_/A VGND VGND VPWR VPWR _1503_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1035_ _0859_/B _1033_/X _1034_/X _1105_/A VGND VGND VPWR VPWR _1523_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ _0826_/A _0819_/B VGND VGND VPWR VPWR _1592_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1584_ _1584_/CLK _1584_/D VGND VGND VPWR VPWR _1584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1365__59 clkload8/A VGND VGND VPWR VPWR _1517_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ _1289_/A _1030_/B VGND VGND VPWR VPWR _1018_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1567_ _1567_/CLK _1567_/D VGND VGND VPWR VPWR _1567_/Q sky130_fd_sc_hd__dfxtp_1
X_1498_ _1498_/CLK _1498_/D VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
Xfanout34 _1016_/A VGND VGND VPWR VPWR _1071_/A sky130_fd_sc_hd__buf_2
Xfanout12 _0930_/Y VGND VGND VPWR VPWR _0963_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout56 _1105_/A VGND VGND VPWR VPWR _1022_/A sky130_fd_sc_hd__clkbuf_2
Xfanout45 _1525_/Q VGND VGND VPWR VPWR _1075_/A sky130_fd_sc_hd__clkbuf_4
Xfanout23 _1285_/C1 VGND VGND VPWR VPWR _1281_/B1 sky130_fd_sc_hd__buf_2
XFILLER_0_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1335__29 clkload5/A VGND VGND VPWR VPWR _1487_/CLK sky130_fd_sc_hd__inv_2
X_1283_ _1283_/A1 _1282_/X _1281_/X _1287_/C1 VGND VGND VPWR VPWR _1283_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload9 clkload9/A VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_8
X_0998_ hold29/A _1534_/Q _1535_/Q _1536_/Q VGND VGND VPWR VPWR _0999_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0753__2 clkload5/A VGND VGND VPWR VPWR _1308_/B sky130_fd_sc_hd__inv_2
X_0921_ _1558_/Q _0960_/B _0944_/C _0921_/D VGND VGND VPWR VPWR _0925_/D sky130_fd_sc_hd__and4_1
X_0783_ _0732_/Y _1594_/Q _1595_/Q _0731_/Y _0766_/X VGND VGND VPWR VPWR _0789_/D
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0852_ hold21/A _0930_/B _0974_/B VGND VGND VPWR VPWR _0852_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 ui_in[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
X_1197_ hold45/A _1511_/Q _1488_/Q VGND VGND VPWR VPWR _1201_/B sky130_fd_sc_hd__mux2_1
X_1266_ _1462_/Q _1285_/A2 _1285_/C1 _1265_/X VGND VGND VPWR VPWR _1266_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1120_ hold36/X _1120_/B VGND VGND VPWR VPWR _1495_/D sky130_fd_sc_hd__xnor2_1
X_1051_ _1051_/A _1051_/B VGND VGND VPWR VPWR _1051_/X sky130_fd_sc_hd__or2_2
XFILLER_0_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0904_ _0904_/A _0904_/B VGND VGND VPWR VPWR _1569_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0766_ hold18/A hold40/A VGND VGND VPWR VPWR _0766_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0835_ _0727_/Y hold16/A _1582_/Q _0726_/Y _0834_/X VGND VGND VPWR VPWR _0835_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1249_ hold37/X _1288_/A2 _1248_/X _1284_/C1 VGND VGND VPWR VPWR _1465_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1406__100 clkload1/A VGND VGND VPWR VPWR _1558_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1103_ _1075_/B _1285_/C1 _1087_/Y _1102_/X VGND VGND VPWR VPWR _1103_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1034_ _1523_/Q _1048_/B VGND VGND VPWR VPWR _1034_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0749_ hold31/A VGND VGND VPWR VPWR _0749_/Y sky130_fd_sc_hd__inv_2
X_0818_ _0823_/A1 _1592_/Q _0813_/Y _0813_/B _0864_/B VGND VGND VPWR VPWR _0819_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1583_ _1583_/CLK _1583_/D VGND VGND VPWR VPWR _1583_/Q sky130_fd_sc_hd__dfxtp_1
X_1017_ _1082_/B _1138_/A _1016_/X _1145_/A VGND VGND VPWR VPWR _1531_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1566_ _1566_/CLK _1566_/D VGND VGND VPWR VPWR _1566_/Q sky130_fd_sc_hd__dfxtp_1
X_1497_ _1497_/CLK _1497_/D VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout46 _0736_/A VGND VGND VPWR VPWR _1075_/B sky130_fd_sc_hd__clkbuf_4
Xfanout13 _1219_/X VGND VGND VPWR VPWR _1287_/C1 sky130_fd_sc_hd__buf_2
Xfanout24 _1081_/X VGND VGND VPWR VPWR _1285_/C1 sky130_fd_sc_hd__buf_2
Xfanout35 _1530_/Q VGND VGND VPWR VPWR _1016_/A sky130_fd_sc_hd__clkbuf_2
Xfanout57 input1/X VGND VGND VPWR VPWR _1105_/A sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1282_ _1459_/Q _1457_/Q _1282_/S VGND VGND VPWR VPWR _1282_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1618_ _1618_/A VGND VGND VPWR VPWR uio_out[7] sky130_fd_sc_hd__buf_2
X_0997_ hold11/X _0967_/D _0996_/Y VGND VGND VPWR VPWR _1537_/D sky130_fd_sc_hd__a21oi_1
X_1549_ _1549_/CLK _1549_/D VGND VGND VPWR VPWR _1549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0920_ _0920_/A VGND VGND VPWR VPWR _0920_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0782_ _1549_/Q _0747_/Y _1594_/Q _0732_/Y _0781_/Y VGND VGND VPWR VPWR _0789_/C
+ sky130_fd_sc_hd__o221a_1
X_0851_ _0791_/C _0850_/Y _0974_/A VGND VGND VPWR VPWR _0930_/B sky130_fd_sc_hd__o21a_1
X_1265_ hold54/A _1280_/B VGND VGND VPWR VPWR _1265_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 ui_in[1] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1196_ _1196_/A _1196_/B _1196_/C VGND VGND VPWR VPWR _1473_/D sky130_fd_sc_hd__and3_1
X_1423__117 clkload6/A VGND VGND VPWR VPWR _1575_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _1051_/A _1051_/B VGND VGND VPWR VPWR _1066_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0834_ _1564_/Q _1584_/Q VGND VGND VPWR VPWR _0834_/X sky130_fd_sc_hd__xor2_1
X_0903_ _0903_/A1 _0743_/Y _0889_/Y _0889_/B _1069_/B VGND VGND VPWR VPWR _0904_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0765_ _1592_/Q _1554_/Q VGND VGND VPWR VPWR _0765_/X sky130_fd_sc_hd__and2b_1
X_1248_ _1283_/A1 _1247_/X _1246_/X _1287_/C1 VGND VGND VPWR VPWR _1248_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ _1152_/A _1122_/C _1125_/Y _1150_/X _1178_/Y VGND VGND VPWR VPWR _1179_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1102_ _1292_/B _1100_/Y _1101_/X _1098_/S VGND VGND VPWR VPWR _1102_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1033_ _1051_/A _1033_/B VGND VGND VPWR VPWR _1033_/X sky130_fd_sc_hd__or2_2
XFILLER_0_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0817_ _0826_/A _0817_/B VGND VGND VPWR VPWR _1593_/D sky130_fd_sc_hd__and2_1
X_0748_ _1588_/Q VGND VGND VPWR VPWR _0748_/Y sky130_fd_sc_hd__inv_2
X_1429__123 clkload2/A VGND VGND VPWR VPWR _1581_/CLK sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1582_ _1582_/CLK _1582_/D VGND VGND VPWR VPWR _1582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1016_ _1016_/A _1030_/B VGND VGND VPWR VPWR _1016_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1370__64 clkload9/A VGND VGND VPWR VPWR _1522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1565_ _1565_/CLK _1565_/D VGND VGND VPWR VPWR _1565_/Q sky130_fd_sc_hd__dfxtp_2
X_1496_ _1496_/CLK _1496_/D VGND VGND VPWR VPWR _1496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout58 _1303_/C1 VGND VGND VPWR VPWR _1294_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_32_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout14 _1218_/Y VGND VGND VPWR VPWR _1288_/A2 sky130_fd_sc_hd__buf_2
XFILLER_0_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout25 _0864_/Y VGND VGND VPWR VPWR _1285_/A2 sky130_fd_sc_hd__buf_2
Xfanout47 _1524_/Q VGND VGND VPWR VPWR _0736_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout36 _0864_/B VGND VGND VPWR VPWR _1289_/A sky130_fd_sc_hd__buf_2
X_1281_ _1459_/Q _1285_/A2 _1281_/B1 _1280_/X VGND VGND VPWR VPWR _1281_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0996_ hold11/X _0967_/D _1004_/B VGND VGND VPWR VPWR _0996_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1617_ _1617_/A VGND VGND VPWR VPWR uio_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1479_ _1483_/CLK input5/X VGND VGND VPWR VPWR _1479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1548_ _1548_/CLK _1548_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1340__34 clkload3/A VGND VGND VPWR VPWR _1492_/CLK sky130_fd_sc_hd__inv_2
X_0850_ _0850_/A _0850_/B _0850_/C VGND VGND VPWR VPWR _0850_/Y sky130_fd_sc_hd__nor3_1
X_0781_ _1564_/Q _1602_/Q VGND VGND VPWR VPWR _0781_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 ui_in[2] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
X_1264_ _1462_/Q _1218_/Y _1263_/X _1303_/C1 VGND VGND VPWR VPWR _1462_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1195_ _1618_/A _1194_/Y _1195_/S VGND VGND VPWR VPWR _1196_/C sky130_fd_sc_hd__mux2_1
X_0979_ hold5/X _0981_/A _0978_/Y VGND VGND VPWR VPWR _1546_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0902_ _0915_/A _0902_/B VGND VGND VPWR VPWR _1570_/D sky130_fd_sc_hd__and2_1
X_0833_ _1551_/Q _1571_/Q VGND VGND VPWR VPWR _0833_/X sky130_fd_sc_hd__and2b_1
X_0764_ _0758_/X _0760_/X _0763_/X _1568_/Q VGND VGND VPWR VPWR _0974_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1247_ hold41/A hold35/A _1277_/S VGND VGND VPWR VPWR _1247_/X sky130_fd_sc_hd__mux2_1
X_1178_ _1178_/A _1486_/Q _1152_/B VGND VGND VPWR VPWR _1178_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ _1169_/B _1301_/A uo_out[4] VGND VGND VPWR VPWR _1101_/X sky130_fd_sc_hd__a21o_1
X_1032_ _1051_/A _1033_/B VGND VGND VPWR VPWR _1048_/B sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0747_ _1587_/Q VGND VGND VPWR VPWR _0747_/Y sky130_fd_sc_hd__inv_2
X_0816_ _1196_/B _1593_/Q _0813_/Y _0813_/B _1530_/Q VGND VGND VPWR VPWR _0817_/B
+ sky130_fd_sc_hd__a32o_1
X_1376__70 clkload4/A VGND VGND VPWR VPWR _1528_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1581_ _1581_/CLK _1581_/D VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
X_1015_ _1173_/B _1152_/A _1173_/A VGND VGND VPWR VPWR _1105_/D sky130_fd_sc_hd__a21o_2
XFILLER_0_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1564_ _1564_/CLK _1564_/D VGND VGND VPWR VPWR _1564_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_18_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1346__40 clkload8/A VGND VGND VPWR VPWR _1498_/CLK sky130_fd_sc_hd__inv_2
X_1495_ _1495_/CLK _1495_/D VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfxtp_1
Xfanout26 _1275_/B VGND VGND VPWR VPWR _1280_/B sky130_fd_sc_hd__clkbuf_2
Xfanout15 _0974_/Y VGND VGND VPWR VPWR _0983_/B sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout37 _1529_/Q VGND VGND VPWR VPWR _0864_/B sky130_fd_sc_hd__buf_2
Xfanout59 _1303_/C1 VGND VGND VPWR VPWR _1284_/C1 sky130_fd_sc_hd__buf_2
Xfanout48 _1487_/Q VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_32_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _1457_/Q _1280_/B VGND VGND VPWR VPWR _1280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ _0966_/X _1004_/B _0995_/C VGND VGND VPWR VPWR _1538_/D sky130_fd_sc_hd__and3b_1
X_1616_ hold2/A VGND VGND VPWR VPWR uio_out[2] sky130_fd_sc_hd__clkbuf_4
X_1547_ _1547_/CLK _1547_/D VGND VGND VPWR VPWR _1547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1478_ _1483_/CLK input4/X VGND VGND VPWR VPWR _1478_/Q sky130_fd_sc_hd__dfxtp_1
X_0780_ _0731_/Y _1595_/Q _0752_/Y _1562_/Q _0779_/Y VGND VGND VPWR VPWR _0789_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_1_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 ui_in[3] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
X_1263_ _1098_/S _1262_/X _1261_/X _1219_/X VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__a211o_1
X_1316__10 _1475_/CLK VGND VGND VPWR VPWR _1459_/CLK sky130_fd_sc_hd__inv_2
X_1194_ hold34/A _1192_/A _1618_/A VGND VGND VPWR VPWR _1194_/Y sky130_fd_sc_hd__a21oi_1
X_0978_ hold5/X _0981_/A _0983_/B VGND VGND VPWR VPWR _0978_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400__94 _1400__94/A VGND VGND VPWR VPWR _1552_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_36_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0763_ _0761_/X _0762_/X _1567_/Q VGND VGND VPWR VPWR _0763_/X sky130_fd_sc_hd__mux2_1
X_0832_ _1556_/Q _1576_/Q VGND VGND VPWR VPWR _0832_/Y sky130_fd_sc_hd__nand2b_1
X_0901_ _0802_/B _1570_/Q _0889_/Y _0889_/B _1525_/Q VGND VGND VPWR VPWR _0902_/B
+ sky130_fd_sc_hd__a32o_1
X_1177_ _1486_/Q _1126_/B _1176_/X _1145_/A VGND VGND VPWR VPWR _1486_/D sky130_fd_sc_hd__o211a_1
X_1246_ hold41/A _0864_/Y _1281_/B1 _1245_/X VGND VGND VPWR VPWR _1246_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_9_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload6/A sky130_fd_sc_hd__clkbuf_8
X_1413__107 clkload8/A VGND VGND VPWR VPWR _1565_/CLK sky130_fd_sc_hd__inv_2
X_1100_ _1169_/B _1301_/A VGND VGND VPWR VPWR _1100_/Y sky130_fd_sc_hd__nand2_1
X_1031_ _1075_/B _1138_/A _1030_/X _1294_/A VGND VGND VPWR VPWR _1524_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0746_ _1583_/Q VGND VGND VPWR VPWR _0829_/B sky130_fd_sc_hd__inv_2
X_0815_ _0826_/A _0815_/B VGND VGND VPWR VPWR _1594_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1391__85 clkload7/A VGND VGND VPWR VPWR _1543_/CLK sky130_fd_sc_hd__inv_2
X_1229_ hold39/X _1288_/A2 _1228_/X _1284_/C1 VGND VGND VPWR VPWR _1469_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1580_/CLK _1580_/D VGND VGND VPWR VPWR _1580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _1173_/B _1152_/A _1173_/A VGND VGND VPWR VPWR _1030_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ _1559_/Q VGND VGND VPWR VPWR _0729_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1563_ _1563_/CLK _1563_/D VGND VGND VPWR VPWR _1563_/Q sky130_fd_sc_hd__dfxtp_1
X_1419__113 clkload6/A VGND VGND VPWR VPWR _1571_/CLK sky130_fd_sc_hd__inv_2
X_1494_ _1494_/CLK _1494_/D VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
X_1361__55 clkload3/A VGND VGND VPWR VPWR _1513_/CLK sky130_fd_sc_hd__inv_2
Xfanout16 _0974_/Y VGND VGND VPWR VPWR _1004_/B sky130_fd_sc_hd__buf_1
Xfanout27 _1196_/B VGND VGND VPWR VPWR _0823_/A1 sky130_fd_sc_hd__buf_2
Xfanout49 _0828_/A VGND VGND VPWR VPWR _0826_/A sky130_fd_sc_hd__clkbuf_2
Xfanout38 _1528_/Q VGND VGND VPWR VPWR _1020_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ hold11/A _0967_/D _1538_/Q VGND VGND VPWR VPWR _0995_/C sky130_fd_sc_hd__a21o_1
X_1477_ _1483_/CLK input3/X VGND VGND VPWR VPWR _1477_/Q sky130_fd_sc_hd__dfxtp_1
X_1615_ hold12/A VGND VGND VPWR VPWR uio_out[1] sky130_fd_sc_hd__clkbuf_4
X_1546_ _1546_/CLK _1546_/D VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 ui_in[4] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
X_1331__25 _1359__53/A VGND VGND VPWR VPWR _1474_/CLK sky130_fd_sc_hd__inv_2
X_1262_ _1463_/Q _1461_/Q _1277_/S VGND VGND VPWR VPWR _1262_/X sky130_fd_sc_hd__mux2_1
X_1193_ hold34/A _1587_/Q _1187_/X _1192_/Y _0930_/B VGND VGND VPWR VPWR _1195_/S
+ sky130_fd_sc_hd__o41a_1
X_0977_ _0973_/X _0983_/B _0977_/C VGND VGND VPWR VPWR _1547_/D sky130_fd_sc_hd__and3b_1
X_1529_ _1529_/CLK _1529_/D VGND VGND VPWR VPWR _1529_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1397__91 _1400__94/A VGND VGND VPWR VPWR _1549_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0915_/A _0900_/B VGND VGND VPWR VPWR _1571_/D sky130_fd_sc_hd__and2_1
X_0762_ hold11/A _1538_/Q hold9/A hold17/A _1565_/Q _1566_/Q VGND VGND VPWR VPWR _0762_/X
+ sky130_fd_sc_hd__mux4_1
X_0831_ _1555_/Q _1575_/Q VGND VGND VPWR VPWR _0831_/X sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_22_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1176_ _1168_/X _1170_/Y _1174_/X _1175_/X _1137_/B VGND VGND VPWR VPWR _1176_/X
+ sky130_fd_sc_hd__a2111o_1
X_1245_ hold35/A _1275_/B VGND VGND VPWR VPWR _1245_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1030_ _1475_/Q _1030_/B VGND VGND VPWR VPWR _1030_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0814_ _0823_/A1 _1594_/Q _0813_/Y _0813_/B _1053_/A1 VGND VGND VPWR VPWR _0815_/B
+ sky130_fd_sc_hd__a32o_1
X_0745_ _1571_/Q VGND VGND VPWR VPWR _0745_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1228_ _1283_/A1 _1227_/X _1226_/X _1287_/C1 VGND VGND VPWR VPWR _1228_/X sky130_fd_sc_hd__a211o_1
X_1159_ _1520_/Q _0739_/Y _0740_/Y _1519_/Q VGND VGND VPWR VPWR _1159_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1367__61 clkload6/A VGND VGND VPWR VPWR _1519_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1013_ _1178_/A _1486_/Q VGND VGND VPWR VPWR _1152_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_8_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0728_ _1560_/Q VGND VGND VPWR VPWR _0937_/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1400__94/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1562_ _1562_/CLK _1562_/D VGND VGND VPWR VPWR _1562_/Q sky130_fd_sc_hd__dfxtp_1
X_1493_ _1493_/CLK hold4/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfxtp_1
Xfanout39 _1169_/A VGND VGND VPWR VPWR _1291_/D sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout28 _1585_/Q VGND VGND VPWR VPWR _1196_/B sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1337__31 _1359__53/A VGND VGND VPWR VPWR _1489_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0993_ _0993_/A _0993_/B VGND VGND VPWR VPWR _1539_/D sky130_fd_sc_hd__nor2_1
X_1614_ _1614_/A VGND VGND VPWR VPWR uio_out[0] sky130_fd_sc_hd__buf_2
X_1476_ _1483_/CLK input2/X VGND VGND VPWR VPWR _1476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1545_ _1545_/CLK _1545_/D VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1261_ _1463_/Q _1285_/A2 _1285_/C1 _1260_/X VGND VGND VPWR VPWR _1261_/X sky130_fd_sc_hd__o211a_1
Xinput7 ui_in[5] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
X_1192_ _1192_/A _1192_/B VGND VGND VPWR VPWR _1192_/Y sky130_fd_sc_hd__nand2_1
X_0976_ hold26/A hold5/A _0972_/B _1547_/Q VGND VGND VPWR VPWR _0977_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_14_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1459_ _1459_/CLK _1459_/D VGND VGND VPWR VPWR _1459_/Q sky130_fd_sc_hd__dfxtp_1
X_1528_ _1528_/CLK _1528_/D VGND VGND VPWR VPWR _1528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0830_ _1557_/Q _1577_/Q VGND VGND VPWR VPWR _0830_/Y sky130_fd_sc_hd__xnor2_1
X_0761_ hold29/A _1534_/Q _1535_/Q _1536_/Q _1565_/Q _1566_/Q VGND VGND VPWR VPWR
+ _0761_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1244_ hold41/X _1218_/Y _1243_/X _1284_/C1 VGND VGND VPWR VPWR _1466_/D sky130_fd_sc_hd__o211a_1
X_1175_ _1149_/Y _1201_/A VGND VGND VPWR VPWR _1175_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0959_ _0942_/X _0959_/B _0959_/C VGND VGND VPWR VPWR _1551_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_33_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 uio_in[3] VGND VGND VPWR VPWR _1475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0813_ _0907_/A _0813_/B VGND VGND VPWR VPWR _0813_/Y sky130_fd_sc_hd__nor2_2
X_0744_ _1570_/Q VGND VGND VPWR VPWR _0744_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1158_ _1519_/Q _0740_/Y _1117_/A _1518_/Q VGND VGND VPWR VPWR _1158_/X sky130_fd_sc_hd__o22a_1
X_1227_ hold27/A hold49/A _1277_/S VGND VGND VPWR VPWR _1227_/X sky130_fd_sc_hd__mux2_1
X_1089_ uo_out[7] _1097_/B _1088_/X _1145_/A VGND VGND VPWR VPWR _1506_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1382__76 clkload8/A VGND VGND VPWR VPWR _1534_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1012_ hold38/A _1484_/Q VGND VGND VPWR VPWR _1173_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0727_ hold40/A VGND VGND VPWR VPWR _0727_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1561_ _1561_/CLK _1561_/D VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfxtp_1
X_1492_ _1492_/CLK _1492_/D VGND VGND VPWR VPWR _1492_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_32_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout29 _0903_/A1 VGND VGND VPWR VPWR _0802_/B sky130_fd_sc_hd__buf_2
Xfanout18 _1105_/D VGND VGND VPWR VPWR _1138_/A sky130_fd_sc_hd__buf_2
X_1352__46 clkload5/A VGND VGND VPWR VPWR _1504_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0992_ hold9/X _0966_/X _0983_/B VGND VGND VPWR VPWR _0993_/B sky130_fd_sc_hd__o21ai_1
X_1613_ hold14/A VGND VGND VPWR VPWR uio_oe[7] sky130_fd_sc_hd__buf_2
X_1544_ _1544_/CLK _1544_/D VGND VGND VPWR VPWR _1544_/Q sky130_fd_sc_hd__dfxtp_1
X_1475_ _1475_/CLK _1475_/D VGND VGND VPWR VPWR _1475_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_7_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload5/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1409__103 clkload0/A VGND VGND VPWR VPWR _1561_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 ui_in[6] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
X_1260_ _1461_/Q _1280_/B VGND VGND VPWR VPWR _1260_/X sky130_fd_sc_hd__or2_1
X_1191_ _1191_/A _1191_/B _1191_/C VGND VGND VPWR VPWR _1192_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0975_ hold1/X _0973_/X _0983_/B VGND VGND VPWR VPWR _1548_/D sky130_fd_sc_hd__o21a_1
X_1527_ _1527_/CLK _1527_/D VGND VGND VPWR VPWR _1527_/Q sky130_fd_sc_hd__dfxtp_1
X_1322__16 clkload11/A VGND VGND VPWR VPWR _1465_/CLK sky130_fd_sc_hd__inv_2
X_1458_ _1458_/CLK _1458_/D VGND VGND VPWR VPWR _1458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0760_ _1567_/Q _0759_/X _1568_/Q VGND VGND VPWR VPWR _0760_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1388__82 clkload7/A VGND VGND VPWR VPWR _1540_/CLK sky130_fd_sc_hd__inv_2
X_1174_ hold38/A _1152_/A _1125_/Y _1173_/X VGND VGND VPWR VPWR _1174_/X sky130_fd_sc_hd__a211o_1
X_1243_ _1283_/A1 _1242_/X _1241_/X _1287_/C1 VGND VGND VPWR VPWR _1243_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_19_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0958_ _1551_/Q _0958_/B VGND VGND VPWR VPWR _0959_/B sky130_fd_sc_hd__or2_1
X_0889_ _0907_/A _0889_/B VGND VGND VPWR VPWR _0889_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_18_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0743_ _1569_/Q VGND VGND VPWR VPWR _0743_/Y sky130_fd_sc_hd__inv_2
X_0812_ _1051_/A _1492_/Q hold48/A VGND VGND VPWR VPWR _0813_/B sky130_fd_sc_hd__nor3b_4
X_1157_ _1518_/Q _1117_/A _1154_/Y _1156_/Y _1155_/X VGND VGND VPWR VPWR _1157_/X
+ sky130_fd_sc_hd__a221o_1
X_1226_ hold27/A _1285_/A2 _1281_/B1 _1225_/X VGND VGND VPWR VPWR _1226_/X sky130_fd_sc_hd__o211a_1
X_1088_ _1207_/A _1285_/C1 _1084_/X _1087_/Y VGND VGND VPWR VPWR _1088_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_7_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1358__52 _1359__53/A VGND VGND VPWR VPWR _1510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1011_ hold38/A _1484_/Q VGND VGND VPWR VPWR _1131_/C sky130_fd_sc_hd__nor2_1
X_0726_ _1562_/Q VGND VGND VPWR VPWR _0726_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ _1482_/Q _1295_/A _1298_/A _1481_/Q VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__a22o_1
X_1442__136 _1450__144/A VGND VGND VPWR VPWR _1594_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1560_ _1560_/CLK _1560_/D VGND VGND VPWR VPWR _1560_/Q sky130_fd_sc_hd__dfxtp_1
X_1491_ _1491_/CLK _1491_/D VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_2
Xfanout19 _1282_/S VGND VGND VPWR VPWR _1277_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1328__22 _1475_/CLK VGND VGND VPWR VPWR _1471_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0991_ _0991_/A _0991_/B VGND VGND VPWR VPWR _1540_/D sky130_fd_sc_hd__nor2_1
X_1612_ hold14/A VGND VGND VPWR VPWR uio_oe[6] sky130_fd_sc_hd__buf_2
X_1474_ _1474_/CLK _1474_/D VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1543_ _1543_/CLK _1543_/D VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1448__142 _1450__144/A VGND VGND VPWR VPWR _1600_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 ui_in[7] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
X_1190_ _1592_/Q _1593_/Q _1594_/Q _1595_/Q VGND VGND VPWR VPWR _1191_/C sky130_fd_sc_hd__or4_1
X_0974_ _0974_/A _0974_/B VGND VGND VPWR VPWR _0974_/Y sky130_fd_sc_hd__nor2_1
X_1457_ _1457_/CLK _1457_/D VGND VGND VPWR VPWR _1457_/Q sky130_fd_sc_hd__dfxtp_1
X_1526_ _1526_/CLK _1526_/D VGND VGND VPWR VPWR _1526_/Q sky130_fd_sc_hd__dfxtp_1
X_1312__6 clkload5/A VGND VGND VPWR VPWR _1455_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_6_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload4/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1173_ _1173_/A _1173_/B _1173_/C VGND VGND VPWR VPWR _1173_/X sky130_fd_sc_hd__and3_1
X_1242_ hold42/A hold37/A _1277_/S VGND VGND VPWR VPWR _1242_/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0957_ hold10/X _0942_/X _0956_/Y VGND VGND VPWR VPWR _1552_/D sky130_fd_sc_hd__a21oi_1
X_0888_ _0888_/A _1051_/B VGND VGND VPWR VPWR _0889_/B sky130_fd_sc_hd__nor2_4
X_1509_ _1509_/CLK _1509_/D VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_jimktrains_vslc_61 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_61/HI uio_oe[3]
+ sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_26_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0742_ _1490_/Q VGND VGND VPWR VPWR _1306_/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_10_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0811_ _0828_/A _0811_/B VGND VGND VPWR VPWR _1595_/D sky130_fd_sc_hd__and2_1
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1087_ _1082_/B _1085_/X _1005_/Y VGND VGND VPWR VPWR _1087_/Y sky130_fd_sc_hd__o21ai_2
X_1156_ hold28/A hold36/A VGND VGND VPWR VPWR _1156_/Y sky130_fd_sc_hd__nand2b_1
X_1225_ hold49/A _1280_/B VGND VGND VPWR VPWR _1225_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_7_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1373__67 clkload4/A VGND VGND VPWR VPWR _1525_/CLK sky130_fd_sc_hd__inv_2
X_1010_ _1486_/Q _1178_/A VGND VGND VPWR VPWR _1173_/A sky130_fd_sc_hd__and2b_1
X_0725_ _1126_/A VGND VGND VPWR VPWR _1068_/A sky130_fd_sc_hd__inv_2
X_1208_ _1480_/Q _1301_/A _1207_/A _1024_/A VGND VGND VPWR VPWR _1208_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_4_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1139_ _1488_/Q _1139_/B VGND VGND VPWR VPWR _1145_/B sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1490_ _1490_/CLK _1490_/D VGND VGND VPWR VPWR _1490_/Q sky130_fd_sc_hd__dfxtp_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1343__37 clkload6/A VGND VGND VPWR VPWR _1495_/CLK sky130_fd_sc_hd__inv_2
X_1611_ hold14/A VGND VGND VPWR VPWR uio_oe[2] sky130_fd_sc_hd__buf_2
X_0990_ hold17/X _0993_/A _0983_/B VGND VGND VPWR VPWR _0991_/B sky130_fd_sc_hd__o21ai_1
X_1542_ _1542_/CLK _1542_/D VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1473_ _1473_/CLK _1473_/D VGND VGND VPWR VPWR _1618_/A sky130_fd_sc_hd__dfxtp_1
X_0973_ hold5/A _1547_/Q _0981_/A VGND VGND VPWR VPWR _0973_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1456_ _1456_/CLK _1456_/D VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
X_1525_ _1525_/CLK _1525_/D VGND VGND VPWR VPWR _1525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1241_ hold42/A _0864_/Y _1281_/B1 _1240_/X VGND VGND VPWR VPWR _1241_/X sky130_fd_sc_hd__o211a_1
X_1172_ _1178_/A _1126_/B _1171_/X _1196_/A VGND VGND VPWR VPWR _1487_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ hold10/X _0942_/X _0963_/B VGND VGND VPWR VPWR _0956_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1379__73 clkload4/A VGND VGND VPWR VPWR _1531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0887_ _1492_/Q hold48/A VGND VGND VPWR VPWR _1051_/B sky130_fd_sc_hd__nand2_2
X_1508_ _1508_/CLK _1508_/D VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfxtp_1
Xmax_cap17 _0791_/C VGND VGND VPWR VPWR _1192_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtt_um_jimktrains_vslc_62 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_62/HI uio_oe[4]
+ sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_1_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0810_ _0823_/A1 _1595_/Q _0792_/Y _0792_/A _0736_/A VGND VGND VPWR VPWR _0811_/B
+ sky130_fd_sc_hd__a32o_1
X_0741_ hold33/X VGND VGND VPWR VPWR _1117_/A sky130_fd_sc_hd__inv_2
X_1224_ hold27/X _1288_/A2 _1223_/X _1284_/C1 VGND VGND VPWR VPWR _1470_/D sky130_fd_sc_hd__o211a_1
X_1086_ _1082_/B _1085_/X _1005_/Y VGND VGND VPWR VPWR _1097_/B sky130_fd_sc_hd__o21a_1
X_1155_ _1496_/Q hold43/A VGND VGND VPWR VPWR _1155_/X sky130_fd_sc_hd__and2b_1
X_0939_ _1559_/Q _0925_/D _0937_/B _0959_/C VGND VGND VPWR VPWR _1559_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_5_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1359__53/A sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_38_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1349__43 clkload11/A VGND VGND VPWR VPWR _1501_/CLK sky130_fd_sc_hd__inv_2
X_1207_ _1207_/A _1207_/B VGND VGND VPWR VPWR _1207_/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1138_ _1138_/A _1138_/B VGND VGND VPWR VPWR _1139_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1069_ _1072_/A _1069_/B VGND VGND VPWR VPWR _1069_/Y sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_26_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1610_ hold14/A VGND VGND VPWR VPWR uio_oe[1] sky130_fd_sc_hd__buf_2
XFILLER_0_26_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1319__13 _1483_/CLK VGND VGND VPWR VPWR _1462_/CLK sky130_fd_sc_hd__inv_2
X_1472_ _1472_/CLK _1472_/D VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ _1541_/CLK _1541_/D VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
X_1432__126 clkload2/A VGND VGND VPWR VPWR _1584_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1403__97 clkload1/A VGND VGND VPWR VPWR _1555_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0972_ hold26/A _0972_/B VGND VGND VPWR VPWR _0981_/A sky130_fd_sc_hd__and2_1
X_1524_ _1524_/CLK _1524_/D VGND VGND VPWR VPWR _1524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1455_ _1455_/CLK _1455_/D VGND VGND VPWR VPWR uo_out[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1171_ _1298_/A _1168_/X _1182_/C _1151_/X VGND VGND VPWR VPWR _1171_/X sky130_fd_sc_hd__a31o_1
X_1240_ hold37/A _1275_/B VGND VGND VPWR VPWR _1240_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0955_ _0952_/B _0955_/B _0959_/C VGND VGND VPWR VPWR _1553_/D sky130_fd_sc_hd__and3b_1
X_0886_ _0904_/A _0886_/B VGND VGND VPWR VPWR _1577_/D sky130_fd_sc_hd__and2_1
X_1507_ _1507_/CLK _1507_/D VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
X_1394__88 _1400__94/A VGND VGND VPWR VPWR _1546_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1438__132 _1450__144/A VGND VGND VPWR VPWR _1590_/CLK sky130_fd_sc_hd__inv_2
Xtt_um_jimktrains_vslc_63 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_63/HI uio_oe[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ hold19/A VGND VGND VPWR VPWR _0740_/Y sky130_fd_sc_hd__inv_2
X_1154_ hold43/A _1496_/Q VGND VGND VPWR VPWR _1154_/Y sky130_fd_sc_hd__nand2b_1
X_1223_ _1283_/A1 _1222_/X _1221_/X _1287_/C1 VGND VGND VPWR VPWR _1223_/X sky130_fd_sc_hd__a211o_1
X_1085_ _1289_/A _1020_/A _1291_/D VGND VGND VPWR VPWR _1085_/X sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_15_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0938_ _0924_/Y _0959_/C _0938_/C VGND VGND VPWR VPWR _1560_/D sky130_fd_sc_hd__and3b_1
X_0869_ hold48/A _1492_/Q VGND VGND VPWR VPWR _1033_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1364__58 clkload6/A VGND VGND VPWR VPWR _1516_/CLK sky130_fd_sc_hd__inv_2
X_1206_ _1479_/Q _1069_/Y _1301_/A _1476_/Q VGND VGND VPWR VPWR _1206_/X sky130_fd_sc_hd__a22o_1
X_1137_ _1201_/A _1137_/B VGND VGND VPWR VPWR _1138_/B sky130_fd_sc_hd__or2_1
X_1068_ _1068_/A hold14/X VGND VGND VPWR VPWR _1507_/D sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload3/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1540_ _1540_/CLK _1540_/D VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1334__28 _1359__53/A VGND VGND VPWR VPWR _1486_/CLK sky130_fd_sc_hd__inv_2
X_1471_ _1471_/CLK _1471_/D VGND VGND VPWR VPWR _1471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0971_ hold6/A _1544_/Q _0987_/A VGND VGND VPWR VPWR _0972_/B sky130_fd_sc_hd__and3_1
X_1454_ _1454_/CLK _1454_/D VGND VGND VPWR VPWR uo_out[2] sky130_fd_sc_hd__dfxtp_4
X_1523_ _1523_/CLK _1523_/D VGND VGND VPWR VPWR _1523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _1298_/A _1182_/C VGND VGND VPWR VPWR _1170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0954_ hold10/A _0942_/X _1553_/Q VGND VGND VPWR VPWR _0955_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ _1196_/B _1577_/Q _0871_/Y _0871_/B _0736_/A VGND VGND VPWR VPWR _0886_/B
+ sky130_fd_sc_hd__a32o_1
X_1506_ _1506_/CLK _1506_/D VGND VGND VPWR VPWR uo_out[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1299_ _1298_/A _1301_/B uo_out[1] VGND VGND VPWR VPWR _1299_/X sky130_fd_sc_hd__a21o_1
Xtt_um_jimktrains_vslc_64 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_64/HI uio_out[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1084_ _1024_/A _1292_/A _1292_/B _1098_/S _1083_/X VGND VGND VPWR VPWR _1084_/X
+ sky130_fd_sc_hd__o311a_1
X_1153_ hold51/A hold24/A VGND VGND VPWR VPWR _1153_/Y sky130_fd_sc_hd__nand2b_1
X_1222_ _1532_/Q hold39/A _1282_/S VGND VGND VPWR VPWR _1222_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0937_ _0937_/A _0937_/B VGND VGND VPWR VPWR _0938_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0799_ _0826_/A _1020_/A VGND VGND VPWR VPWR _0800_/A sky130_fd_sc_hd__and2_2
X_0868_ _0860_/X _0867_/Y _0862_/X VGND VGND VPWR VPWR _1585_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1205_ hold2/X _1138_/B _1204_/X VGND VGND VPWR VPWR _1472_/D sky130_fd_sc_hd__o21ba_1
X_1067_ _0736_/A _1051_/X _1066_/X _1126_/A VGND VGND VPWR VPWR _1508_/D sky130_fd_sc_hd__o211a_1
X_1136_ _1178_/A _1486_/Q _1152_/B _1135_/X VGND VGND VPWR VPWR _1137_/B sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1315__9 _1475_/CLK VGND VGND VPWR VPWR _1458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1119_ _1117_/B _1119_/B VGND VGND VPWR VPWR _1496_/D sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_23_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1470_ _1470_/CLK _1470_/D VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1599_ _1599_/CLK _1599_/D VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload2/A sky130_fd_sc_hd__clkbuf_8
X_0970_ hold23/A _0989_/A VGND VGND VPWR VPWR _0987_/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ _1453_/CLK _1453_/D VGND VGND VPWR VPWR uo_out[1] sky130_fd_sc_hd__dfxtp_4
X_1522_ _1522_/CLK _1522_/D VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1422__116 clkload6/A VGND VGND VPWR VPWR _1574_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0884_ _0904_/A _0884_/B VGND VGND VPWR VPWR _1578_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0953_ _0946_/C _0953_/B _0963_/B VGND VGND VPWR VPWR _1554_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1505_ _1505_/CLK _1505_/D VGND VGND VPWR VPWR uo_out[6] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ _1298_/A _1301_/B VGND VGND VPWR VPWR _1298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtt_um_jimktrains_vslc_65 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_65/HI uio_out[4]
+ sky130_fd_sc_hd__conb_1
X_1385__79 clkload7/A VGND VGND VPWR VPWR _1537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1221_ _1532_/Q _1285_/A2 _1281_/B1 _1220_/X VGND VGND VPWR VPWR _1221_/X sky130_fd_sc_hd__o211a_1
X_1083_ _1169_/B _1075_/A _1075_/B uo_out[7] VGND VGND VPWR VPWR _1083_/X sky130_fd_sc_hd__a31o_1
X_1152_ _1152_/A _1152_/B VGND VGND VPWR VPWR _1168_/A sky130_fd_sc_hd__and2_1
X_0936_ hold40/X _0924_/Y _0926_/Y _0959_/C VGND VGND VPWR VPWR _1561_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0798_ _0826_/A _0798_/B VGND VGND VPWR VPWR _1600_/D sky130_fd_sc_hd__and2_1
X_0867_ _1294_/A _1291_/C _0867_/C _1169_/C VGND VGND VPWR VPWR _0867_/Y sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_38_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1428__122 clkload1/A VGND VGND VPWR VPWR _1580_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1204_ _1138_/B _1199_/Y _1203_/X _1068_/A VGND VGND VPWR VPWR _1204_/X sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1066_ hold44/X _1066_/B VGND VGND VPWR VPWR _1066_/X sky130_fd_sc_hd__or2_1
X_1135_ _1178_/A _1486_/Q hold38/A _1484_/Q VGND VGND VPWR VPWR _1135_/X sky130_fd_sc_hd__and4bb_1
X_0919_ _0960_/B _0944_/C _0921_/D VGND VGND VPWR VPWR _0920_/A sky130_fd_sc_hd__and3_1
X_1355__49 _1359__53/A VGND VGND VPWR VPWR _1507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1049_ _1075_/B _1033_/X _1048_/X _1022_/A VGND VGND VPWR VPWR _1516_/D sky130_fd_sc_hd__o211a_1
X_1118_ _1105_/A hold36/A _1105_/D _1496_/Q VGND VGND VPWR VPWR _1119_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1598_ _1598_/CLK _1598_/D VGND VGND VPWR VPWR _1598_/Q sky130_fd_sc_hd__dfxtp_1
X_1325__19 clkload11/A VGND VGND VPWR VPWR _1468_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_34_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1452_ _1452_/CLK _1452_/D VGND VGND VPWR VPWR uo_out[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1521_ _1521_/CLK _1521_/D VGND VGND VPWR VPWR _1521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ _1554_/Q _0952_/B VGND VGND VPWR VPWR _0953_/B sky130_fd_sc_hd__or2_1
X_1504_ _1504_/CLK _1504_/D VGND VGND VPWR VPWR uo_out[5] sky130_fd_sc_hd__dfxtp_4
X_0883_ _0903_/A1 _1578_/Q _0871_/Y _0871_/B _1525_/Q VGND VGND VPWR VPWR _0884_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1297_ _1292_/B _1295_/Y _1296_/X _1294_/A VGND VGND VPWR VPWR _1454_/D sky130_fd_sc_hd__o211a_1
X_1445__139 clkload0/A VGND VGND VPWR VPWR _1597_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload1/A sky130_fd_sc_hd__clkbuf_8
Xtt_um_jimktrains_vslc_66 VGND VGND VPWR VPWR tt_um_jimktrains_vslc_66/HI uio_out[5]
+ sky130_fd_sc_hd__conb_1
X_1151_ _1173_/A _1131_/C _1125_/Y _1137_/B _1150_/X VGND VGND VPWR VPWR _1151_/X
+ sky130_fd_sc_hd__a2111o_1
X_1220_ hold39/A _1280_/B VGND VGND VPWR VPWR _1220_/X sky130_fd_sc_hd__or2_1
X_1082_ _1016_/A _1082_/B VGND VGND VPWR VPWR _1082_/Y sky130_fd_sc_hd__nand2b_1
X_0935_ _1562_/Q _0928_/C _0927_/Y _0959_/C VGND VGND VPWR VPWR _1562_/D sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_21_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0866_ _1289_/A _1020_/A VGND VGND VPWR VPWR _1169_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0797_ _0823_/A1 _1600_/Q _0792_/Y _0792_/A _0864_/B VGND VGND VPWR VPWR _0798_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1203_ _1489_/Q _1201_/Y _1202_/Y _1201_/A _1490_/Q VGND VGND VPWR VPWR _1203_/X
+ sky130_fd_sc_hd__a221o_1
X_1134_ hold38/A _1484_/Q VGND VGND VPWR VPWR _1152_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1065_ _1075_/A _1051_/X _1064_/X _1126_/A VGND VGND VPWR VPWR _1509_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_7_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0918_ _1557_/Q _1556_/Q _1555_/Q _1554_/Q VGND VGND VPWR VPWR _0921_/D sky130_fd_sc_hd__and4_1
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0849_ _0849_/A _0849_/B _0849_/C _0849_/D VGND VGND VPWR VPWR _0850_/C sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_3_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_1117_ _1117_/A _1117_/B VGND VGND VPWR VPWR _1497_/D sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ hold28/X _1048_/B VGND VGND VPWR VPWR _1048_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1597_ _1597_/CLK _1597_/D VGND VGND VPWR VPWR _1597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1520_ _1520_/CLK _1520_/D VGND VGND VPWR VPWR _1520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1451_ _1451_/CLK _1451_/D VGND VGND VPWR VPWR _1617_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0882_ _0904_/A _0882_/B VGND VGND VPWR VPWR _1579_/D sky130_fd_sc_hd__and2_1
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0951_ _0951_/A _0951_/B VGND VGND VPWR VPWR _1555_/D sky130_fd_sc_hd__nor2_1
X_1503_ _1503_/CLK _1503_/D VGND VGND VPWR VPWR uo_out[4] sky130_fd_sc_hd__dfxtp_4
X_1296_ _1295_/A _1301_/B uo_out[2] VGND VGND VPWR VPWR _1296_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1150_ _1178_/A _1133_/Y _1149_/Y _1201_/A VGND VGND VPWR VPWR _1150_/X sky130_fd_sc_hd__a22o_1
X_1081_ _1071_/A _1082_/B VGND VGND VPWR VPWR _1081_/X sky130_fd_sc_hd__and2b_1
X_0865_ _1471_/Q _1280_/B VGND VGND VPWR VPWR _0867_/C sky130_fd_sc_hd__or2_1
X_0934_ _0931_/B _0959_/C _0934_/C VGND VGND VPWR VPWR _1563_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1412__106 clkload0/A VGND VGND VPWR VPWR _1564_/CLK sky130_fd_sc_hd__inv_2
X_0796_ _0826_/A _0796_/B VGND VGND VPWR VPWR _1601_/D sky130_fd_sc_hd__and2_1
X_1279_ _1459_/Q _1288_/A2 _1278_/X _1284_/C1 VGND VGND VPWR VPWR _1459_/D sky130_fd_sc_hd__o211a_1
X_1390__84 clkload7/A VGND VGND VPWR VPWR _1542_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1202_ _1489_/Q _1202_/B VGND VGND VPWR VPWR _1202_/Y sky130_fd_sc_hd__nor2_1
X_1064_ hold53/X _1066_/B VGND VGND VPWR VPWR _1064_/X sky130_fd_sc_hd__or2_1
X_1133_ _1486_/Q _1173_/C VGND VGND VPWR VPWR _1133_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_4_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1450__144/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0917_ _1553_/Q hold10/A _1551_/Q _1550_/Q VGND VGND VPWR VPWR _0944_/C sky130_fd_sc_hd__and4_1
XFILLER_0_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0848_ _0729_/Y _1579_/Q _1580_/Q _0937_/A _0832_/Y VGND VGND VPWR VPWR _0849_/D
+ sky130_fd_sc_hd__o221a_1
X_0779_ _1563_/Q _1601_/Q VGND VGND VPWR VPWR _0779_/Y sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_3_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1047_ _1525_/Q _1033_/X _1046_/X _1105_/A VGND VGND VPWR VPWR _1517_/D sky130_fd_sc_hd__o211a_1
X_1116_ _1116_/A hold20/X VGND VGND VPWR VPWR _1498_/D sky130_fd_sc_hd__nor2_1
X_1360__54 clkload3/A VGND VGND VPWR VPWR _1512_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1418__112 clkload6/A VGND VGND VPWR VPWR _1570_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ _1596_/CLK _1596_/D VGND VGND VPWR VPWR _1596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1330__24 clkload2/A VGND VGND VPWR VPWR _1473_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1579_ _1579_/CLK _1579_/D VGND VGND VPWR VPWR _1579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1396__90 _1400__94/A VGND VGND VPWR VPWR _1548_/CLK sky130_fd_sc_hd__inv_2
X_0950_ _1555_/Q _0946_/C _0959_/C VGND VGND VPWR VPWR _0951_/B sky130_fd_sc_hd__o21ai_1
X_0881_ _0903_/A1 _1579_/Q _0871_/Y _0871_/B _0734_/A VGND VGND VPWR VPWR _0882_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1502_ _1502_/CLK _1502_/D VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfxtp_1
X_1295_ _1295_/A _1301_/B VGND VGND VPWR VPWR _1295_/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1080_ _0856_/X _1207_/B _1071_/X _1471_/Q VGND VGND VPWR VPWR _1292_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_23_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0933_ _1562_/Q _0928_/C _1563_/Q VGND VGND VPWR VPWR _0934_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0795_ _0823_/A1 _1601_/Q _0792_/Y _0792_/A _1530_/Q VGND VGND VPWR VPWR _0796_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0864_ _1020_/A _0864_/B VGND VGND VPWR VPWR _0864_/Y sky130_fd_sc_hd__nand2b_2
X_1278_ _1283_/A1 _1277_/X _1276_/X _1287_/C1 VGND VGND VPWR VPWR _1278_/X sky130_fd_sc_hd__a211o_1
X_1366__60 clkload8/A VGND VGND VPWR VPWR _1518_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1201_ _1201_/A _1201_/B VGND VGND VPWR VPWR _1201_/Y sky130_fd_sc_hd__nand2_1
X_1435__129 clkload2/A VGND VGND VPWR VPWR _1587_/CLK sky130_fd_sc_hd__inv_2
X_1063_ _1063_/A1 _1051_/X _1062_/X _1126_/A VGND VGND VPWR VPWR _1510_/D sky130_fd_sc_hd__o211a_1
X_1132_ hold38/A _1484_/Q VGND VGND VPWR VPWR _1173_/C sky130_fd_sc_hd__nand2_1
X_0916_ _0758_/X _0760_/X _0763_/X _1568_/Q _1549_/Q VGND VGND VPWR VPWR _0960_/B
+ sky130_fd_sc_hd__o221a_2
X_0778_ _1555_/Q _0750_/Y _1596_/Q _0730_/Y VGND VGND VPWR VPWR _0778_/X sky130_fd_sc_hd__a2bb2o_1
X_0847_ _0733_/Y hold15/A hold16/A _0727_/Y _0830_/Y VGND VGND VPWR VPWR _0849_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_1046_ hold43/X _1048_/B VGND VGND VPWR VPWR _1046_/X sky130_fd_sc_hd__or2_1
X_1115_ hold33/A _1117_/B hold19/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1336__30 _1359__53/A VGND VGND VPWR VPWR _1488_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload0/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1595_ _1595_/CLK _1595_/D VGND VGND VPWR VPWR _1595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1029_ _1075_/A _1138_/A _1028_/Y _1022_/A VGND VGND VPWR VPWR _1525_/D sky130_fd_sc_hd__o211a_1
X_1578_ _1578_/CLK _1578_/D VGND VGND VPWR VPWR _1578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_38_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0880_ _0904_/A _0880_/B VGND VGND VPWR VPWR _1580_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1501_ _1501_/CLK _1501_/D VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
X_1294_ _1294_/A _1294_/B _1294_/C VGND VGND VPWR VPWR _1455_/D sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_18_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0932_ _0932_/A _0959_/C _0932_/C VGND VGND VPWR VPWR _1564_/D sky130_fd_sc_hd__and3_1
XFILLER_0_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0794_ _0826_/A _0794_/B VGND VGND VPWR VPWR _1602_/D sky130_fd_sc_hd__and2_1
X_0863_ _1020_/A _0864_/B VGND VGND VPWR VPWR _1275_/B sky130_fd_sc_hd__and2b_1
X_1277_ hold54/A _1458_/Q _1277_/S VGND VGND VPWR VPWR _1277_/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1381__75 clkload8/A VGND VGND VPWR VPWR _1533_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ hold44/A hold53/A _1488_/Q VGND VGND VPWR VPWR _1202_/B sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1062_ hold45/X _1066_/B VGND VGND VPWR VPWR _1062_/X sky130_fd_sc_hd__or2_1
X_1131_ _1178_/A _1486_/Q _1131_/C VGND VGND VPWR VPWR _1201_/A sky130_fd_sc_hd__and3_1
X_0915_ _0915_/A _0915_/B VGND VGND VPWR VPWR _1565_/D sky130_fd_sc_hd__and2_1
X_0846_ _0846_/A _0846_/B VGND VGND VPWR VPWR _0849_/B sky130_fd_sc_hd__nor2_1
X_0777_ _1589_/Q _1551_/Q VGND VGND VPWR VPWR _0777_/Y sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_3_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1114_ _1114_/A _1114_/B VGND VGND VPWR VPWR _1499_/D sky130_fd_sc_hd__nor2_1
X_1045_ _0734_/A _1033_/X _1044_/X _1105_/A VGND VGND VPWR VPWR _1518_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0829_ _1563_/Q _0829_/B VGND VGND VPWR VPWR _0829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1351__45 clkload5/A VGND VGND VPWR VPWR _1503_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1594_ _1594_/CLK _1594_/D VGND VGND VPWR VPWR _1594_/Q sky130_fd_sc_hd__dfxtp_1
X_1028_ _1069_/B _1138_/A VGND VGND VPWR VPWR _1028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1408__102 clkload0/A VGND VGND VPWR VPWR _1560_/CLK sky130_fd_sc_hd__inv_2
X_1577_ _1577_/CLK _1577_/D VGND VGND VPWR VPWR _1577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1321__15 _1483_/CLK VGND VGND VPWR VPWR _1464_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_27_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1500_ _1500_/CLK _1500_/D VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
X_1293_ _1069_/Y _1301_/B uo_out[3] VGND VGND VPWR VPWR _1294_/C sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1387__81 clkload7/A VGND VGND VPWR VPWR _1539_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0931_ _1564_/Q _0931_/B VGND VGND VPWR VPWR _0932_/C sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0862_ _0862_/A _0974_/B _0860_/X VGND VGND VPWR VPWR _0862_/X sky130_fd_sc_hd__or3b_1
X_0793_ _1196_/B _1602_/Q _0792_/Y _0792_/A _1053_/A1 VGND VGND VPWR VPWR _0794_/B
+ sky130_fd_sc_hd__a32o_1
X_1276_ hold54/A _1285_/A2 _1281_/B1 _1275_/X VGND VGND VPWR VPWR _1276_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1357__51 _1359__53/A VGND VGND VPWR VPWR _1509_/CLK sky130_fd_sc_hd__inv_2
X_1130_ _1484_/Q hold48/X _1130_/S VGND VGND VPWR VPWR _1491_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_34_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ _1169_/A _1051_/X _1060_/X _1126_/A VGND VGND VPWR VPWR _1511_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0845_ _1558_/Q _1578_/Q VGND VGND VPWR VPWR _0846_/B sky130_fd_sc_hd__xor2_1
X_0914_ _0802_/B _1565_/Q _0907_/Y _0907_/B _1075_/B VGND VGND VPWR VPWR _0915_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0776_ _1551_/Q _1589_/Q VGND VGND VPWR VPWR _0776_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ _1463_/Q _1218_/Y _1258_/X _1284_/C1 VGND VGND VPWR VPWR _1463_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1310__4 _1475_/CLK VGND VGND VPWR VPWR _1453_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1441__135 _1450__144/A VGND VGND VPWR VPWR _1593_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1044_ _1518_/Q _1048_/B VGND VGND VPWR VPWR _1044_/X sky130_fd_sc_hd__or2_1
X_1113_ hold22/X _1116_/A VGND VGND VPWR VPWR _1114_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0759_ hold26/A hold5/A _1547_/Q hold1/A _1565_/Q _1566_/Q VGND VGND VPWR VPWR _0759_/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0828_ _0828_/A _0828_/B VGND VGND VPWR VPWR _1587_/D sky130_fd_sc_hd__and2_1
X_1425__119 clkload1/A VGND VGND VPWR VPWR _1577_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1327__21 clkload9/A VGND VGND VPWR VPWR _1470_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1593_ _1593_/CLK _1593_/D VGND VGND VPWR VPWR _1593_/Q sky130_fd_sc_hd__dfxtp_1
X_1027_ _1063_/A1 _1138_/A _1026_/Y _1145_/A VGND VGND VPWR VPWR _1526_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1447__141 _1450__144/A VGND VGND VPWR VPWR _1599_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1576_ _1576_/CLK _1576_/D VGND VGND VPWR VPWR _1576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ _1292_/A _1292_/B _1301_/B VGND VGND VPWR VPWR _1294_/B sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_18_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1559_ _1559_/CLK _1559_/D VGND VGND VPWR VPWR _1559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0930_ _0974_/B _0930_/B VGND VGND VPWR VPWR _0930_/Y sky130_fd_sc_hd__nor2_1
X_0792_ _0792_/A _0907_/A VGND VGND VPWR VPWR _0792_/Y sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_15_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0861_ _1207_/A _1289_/C _0856_/X _0907_/A VGND VGND VPWR VPWR _0862_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1275_ _1458_/Q _1275_/B VGND VGND VPWR VPWR _1275_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ _1511_/Q _1066_/B VGND VGND VPWR VPWR _1060_/X sky130_fd_sc_hd__or2_1
X_1372__66 _1475_/CLK VGND VGND VPWR VPWR _1524_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0844_ hold10/A _1572_/Q VGND VGND VPWR VPWR _0846_/A sky130_fd_sc_hd__xor2_1
X_0913_ _0915_/A _0913_/B VGND VGND VPWR VPWR _1566_/D sky130_fd_sc_hd__and2_1
X_0775_ _1559_/Q _1597_/Q VGND VGND VPWR VPWR _0775_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1258_ _1098_/S _1257_/X _1256_/X _1219_/X VGND VGND VPWR VPWR _1258_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1189_ _1596_/Q _1597_/Q _1598_/Q hold18/A VGND VGND VPWR VPWR _1191_/B sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1043_ _1291_/D _1033_/X _1042_/X _1022_/A VGND VGND VPWR VPWR _1519_/D sky130_fd_sc_hd__o211a_1
X_1112_ _1112_/A _1114_/A VGND VGND VPWR VPWR _1500_/D sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0758_ _1567_/Q _0758_/B VGND VGND VPWR VPWR _0758_/X sky130_fd_sc_hd__and2b_1
X_0827_ _1196_/B _1587_/Q _0813_/Y _0813_/B _0736_/A VGND VGND VPWR VPWR _0828_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1342__36 clkload3/A VGND VGND VPWR VPWR _1494_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1592_ _1592_/CLK _1592_/D VGND VGND VPWR VPWR _1592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1026_ _1072_/A _1138_/A VGND VGND VPWR VPWR _1026_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1575_ _1575_/CLK _1575_/D VGND VGND VPWR VPWR _1575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1009_ _1294_/A _1009_/B _1009_/C VGND VGND VPWR VPWR _1532_/D sky130_fd_sc_hd__and3_1
XFILLER_0_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1291_ _0734_/A _1289_/C _1291_/C _1291_/D VGND VGND VPWR VPWR _1301_/B sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_18_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1489_ _1489_/CLK _1489_/D VGND VGND VPWR VPWR _1489_/Q sky130_fd_sc_hd__dfxtp_4
X_1558_ _1558_/CLK _1558_/D VGND VGND VPWR VPWR _1558_/Q sky130_fd_sc_hd__dfxtp_1
X_1378__72 clkload4/A VGND VGND VPWR VPWR _1530_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ hold34/A _0974_/A _0791_/C VGND VGND VPWR VPWR _0907_/A sky130_fd_sc_hd__and3_2
X_0860_ _1291_/D _1289_/C _1282_/S _0856_/X VGND VGND VPWR VPWR _0860_/X sky130_fd_sc_hd__or4b_1
X_1274_ hold54/X _1288_/A2 _1273_/X _1303_/C1 VGND VGND VPWR VPWR _1460_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0989_/A _0989_/B VGND VGND VPWR VPWR _1541_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ _0802_/B _1566_/Q _0907_/Y _0907_/B _1525_/Q VGND VGND VPWR VPWR _0913_/B
+ sky130_fd_sc_hd__a32o_1
X_0843_ _1550_/Q _0744_/Y _1582_/Q _0726_/Y _0842_/Y VGND VGND VPWR VPWR _0849_/A
+ sky130_fd_sc_hd__o221a_1
X_0774_ _1553_/Q hold31/A VGND VGND VPWR VPWR _0774_/X sky130_fd_sc_hd__and2b_1
X_1348__42 clkload11/A VGND VGND VPWR VPWR _1500_/CLK sky130_fd_sc_hd__inv_2
X_1257_ hold35/A _1462_/Q _1277_/S VGND VGND VPWR VPWR _1257_/X sky130_fd_sc_hd__mux2_1
X_1188_ _1600_/Q _1601_/Q _1602_/Q VGND VGND VPWR VPWR _1191_/A sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_34_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1042_ _1519_/Q _1048_/B VGND VGND VPWR VPWR _1042_/X sky130_fd_sc_hd__or2_1
X_1111_ _1111_/A hold25/X VGND VGND VPWR VPWR _1501_/D sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0757_ hold8/A hold23/A hold6/A _1544_/Q _1565_/Q _1566_/Q VGND VGND VPWR VPWR _0758_/B
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0826_ _0826_/A _0826_/B VGND VGND VPWR VPWR _1588_/D sky130_fd_sc_hd__nand2_1
Xclkbuf_4_15_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1483_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1318__12 _1483_/CLK VGND VGND VPWR VPWR _1461_/CLK sky130_fd_sc_hd__inv_2
X_1591_ _1591_/CLK _1591_/D VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfxtp_1
X_1025_ _1291_/D _1105_/D _1024_/Y _1294_/A VGND VGND VPWR VPWR _1527_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0809_ _0828_/A _0809_/B VGND VGND VPWR VPWR _1596_/D sky130_fd_sc_hd__and2_1
X_1431__125 clkload2/A VGND VGND VPWR VPWR _1583_/CLK sky130_fd_sc_hd__inv_2
X_1402__96 clkload1/A VGND VGND VPWR VPWR _1554_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1415__109 clkload7/A VGND VGND VPWR VPWR _1567_/CLK sky130_fd_sc_hd__inv_2
X_1574_ _1574_/CLK _1574_/D VGND VGND VPWR VPWR _1574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1008_ _0906_/C _1005_/Y _1532_/Q VGND VGND VPWR VPWR _1009_/C sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1290_ _0736_/A hold34/X _1290_/S VGND VGND VPWR VPWR _1456_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1488_ _1488_/CLK _1488_/D VGND VGND VPWR VPWR _1488_/Q sky130_fd_sc_hd__dfxtp_4
X_1393__87 _1400__94/A VGND VGND VPWR VPWR _1545_/CLK sky130_fd_sc_hd__inv_2
X_1557_ _1557_/CLK _1557_/D VGND VGND VPWR VPWR _1557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1437__131 _1450__144/A VGND VGND VPWR VPWR _1589_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0790_ _0790_/A _0790_/B _0790_/C _0789_/X VGND VGND VPWR VPWR _0791_/C sky130_fd_sc_hd__nor4b_1
XFILLER_0_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1273_ _1283_/A1 _1272_/X _1271_/X _1287_/C1 VGND VGND VPWR VPWR _1273_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ hold8/X _0991_/A _0983_/B VGND VGND VPWR VPWR _0989_/B sky130_fd_sc_hd__o21ai_1
X_1609_ hold14/A VGND VGND VPWR VPWR uio_oe[0] sky130_fd_sc_hd__buf_2
XFILLER_0_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0911_ _0915_/A _0911_/B VGND VGND VPWR VPWR _1567_/D sky130_fd_sc_hd__and2_1
X_0842_ _1554_/Q _1574_/Q VGND VGND VPWR VPWR _0842_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0773_ _0727_/Y hold18/A _0752_/Y _1562_/Q VGND VGND VPWR VPWR _0773_/X sky130_fd_sc_hd__a22o_1
X_1256_ hold35/A _1285_/A2 _1281_/B1 _1255_/X VGND VGND VPWR VPWR _1256_/X sky130_fd_sc_hd__o211a_1
X_1363__57 clkload3/A VGND VGND VPWR VPWR _1515_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _1588_/Q _1589_/Q _1590_/Q hold31/A VGND VGND VPWR VPWR _1187_/X sky130_fd_sc_hd__or4_1
XFILLER_0_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1110_ hold32/A _1114_/A hold24/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _1020_/A _1033_/X _1040_/X _1105_/A VGND VGND VPWR VPWR _1520_/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_31_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ _1196_/B _0748_/Y _0813_/Y _0813_/B _1072_/A VGND VGND VPWR VPWR _0826_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0756_ _1492_/Q hold48/A _1051_/A VGND VGND VPWR VPWR _0792_/A sky130_fd_sc_hd__nor3_4
X_1308_ hold12/A _1308_/B VGND VGND VPWR VPWR _1614_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1239_ hold42/X _1218_/Y _1238_/X _1284_/C1 VGND VGND VPWR VPWR _1467_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_19_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ _1590_/CLK _1590_/D VGND VGND VPWR VPWR _1590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1024_ _1024_/A _1105_/D VGND VGND VPWR VPWR _1024_/Y sky130_fd_sc_hd__nand2_1
X_1333__27 clkload5/A VGND VGND VPWR VPWR _1485_/CLK sky130_fd_sc_hd__inv_2
X_0808_ _0823_/A1 _1596_/Q _0792_/Y _0792_/A _1075_/A VGND VGND VPWR VPWR _0809_/B
+ sky130_fd_sc_hd__a32o_1
X_0739_ hold22/A VGND VGND VPWR VPWR _0739_/Y sky130_fd_sc_hd__inv_2
X_1399__93 _1400__94/A VGND VGND VPWR VPWR _1551_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload11/A sky130_fd_sc_hd__clkbuf_8
X_1573_ _1573_/CLK _1573_/D VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1007_ _1007_/A hold27/A _0906_/C VGND VGND VPWR VPWR _1009_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1556_ _1556_/CLK _1556_/D VGND VGND VPWR VPWR _1556_/Q sky130_fd_sc_hd__dfxtp_1
X_1487_ _1487_/CLK _1487_/D VGND VGND VPWR VPWR _1487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1313__7 clkload4/A VGND VGND VPWR VPWR _1456_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1369__63 clkload6/A VGND VGND VPWR VPWR _1521_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1272_ _1461_/Q _1459_/Q _1282_/S VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ _0987_/A _0987_/B VGND VGND VPWR VPWR _1542_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1539_ _1539_/CLK _1539_/D VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0772_ _1560_/Q _1598_/Q VGND VGND VPWR VPWR _0772_/Y sky130_fd_sc_hd__nand2_1
X_0910_ _0802_/B _1567_/Q _0907_/Y _0907_/B _0734_/A VGND VGND VPWR VPWR _0911_/B
+ sky130_fd_sc_hd__a32o_1
X_0841_ _0841_/A _0841_/B _0841_/C _0841_/D VGND VGND VPWR VPWR _0850_/B sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ hold12/X _1139_/B _1178_/Y _1068_/A VGND VGND VPWR VPWR _1474_/D sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ _1462_/Q _1280_/B VGND VGND VPWR VPWR _1255_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1339__33 clkload3/A VGND VGND VPWR VPWR _1491_/CLK sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1040_ _1520_/Q _1048_/B VGND VGND VPWR VPWR _1040_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0824_ _0826_/A _0824_/B VGND VGND VPWR VPWR _1589_/D sky130_fd_sc_hd__and2_1
X_0755_ hold3/A _0854_/A hold7/A VGND VGND VPWR VPWR _1051_/A sky130_fd_sc_hd__or3b_4
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1307_ _1490_/Q _1304_/X _1306_/X _1196_/A VGND VGND VPWR VPWR _1451_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1238_ _1283_/A1 _1237_/X _1236_/X _1219_/X VGND VGND VPWR VPWR _1238_/X sky130_fd_sc_hd__a211o_1
X_1169_ _1169_/A _1169_/B _1169_/C _1289_/D VGND VGND VPWR VPWR _1182_/C sky130_fd_sc_hd__nor4_2
XFILLER_0_19_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ _1291_/D _1030_/B _1120_/B _1289_/B VGND VGND VPWR VPWR _1528_/D sky130_fd_sc_hd__a2bb2oi_1
X_0807_ _0828_/A _0807_/B VGND VGND VPWR VPWR _1597_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0738_ hold32/X VGND VGND VPWR VPWR _1112_/A sky130_fd_sc_hd__inv_2
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1572_ _1572_/CLK _1572_/D VGND VGND VPWR VPWR _1572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1006_ _1071_/A _1289_/C VGND VGND VPWR VPWR _1007_/A sky130_fd_sc_hd__or2_1
XFILLER_0_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421__115 clkload2/A VGND VGND VPWR VPWR _1573_/CLK sky130_fd_sc_hd__inv_2
X_1555_ _1555_/CLK _1555_/D VGND VGND VPWR VPWR _1555_/Q sky130_fd_sc_hd__dfxtp_1
X_1486_ _1486_/CLK _1486_/D VGND VGND VPWR VPWR _1486_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_13_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1475_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_9_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1384__78 clkload8/A VGND VGND VPWR VPWR _1536_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1271_ _1461_/Q _1285_/A2 _1281_/B1 _1270_/X VGND VGND VPWR VPWR _1271_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ hold23/X _0989_/A _0983_/B VGND VGND VPWR VPWR _0987_/B sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1538_ _1538_/CLK _1538_/D VGND VGND VPWR VPWR _1538_/Q sky130_fd_sc_hd__dfxtp_1
X_1469_ _1469_/CLK _1469_/D VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0771_ _1560_/Q _1598_/Q VGND VGND VPWR VPWR _0771_/X sky130_fd_sc_hd__or2_1
X_0840_ _1549_/Q _0743_/Y _0829_/B _1563_/Q _0833_/X VGND VGND VPWR VPWR _0841_/D
+ sky130_fd_sc_hd__a221o_1
X_1254_ hold35/X _1288_/A2 _1253_/X _1284_/C1 VGND VGND VPWR VPWR _1464_/D sky130_fd_sc_hd__o211a_1
X_1185_ _1484_/Q _1126_/B _1183_/Y _1184_/X _1196_/A VGND VGND VPWR VPWR _1484_/D
+ sky130_fd_sc_hd__o221a_1
X_1427__121 clkload1/A VGND VGND VPWR VPWR _1579_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0969_ hold17/A hold8/A _0993_/A VGND VGND VPWR VPWR _0989_/A sky130_fd_sc_hd__and3_1
X_1354__48 clkload5/A VGND VGND VPWR VPWR _1506_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0754_ _1490_/Q _1489_/Q _1488_/Q VGND VGND VPWR VPWR _0854_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0823_ _0823_/A1 _1589_/Q _0813_/Y _0813_/B _1063_/A1 VGND VGND VPWR VPWR _0824_/B
+ sky130_fd_sc_hd__a32o_1
X_1306_ _1306_/A _1306_/B VGND VGND VPWR VPWR _1306_/X sky130_fd_sc_hd__or2_1
X_1099_ _1087_/Y _1098_/X _1097_/X _1294_/A VGND VGND VPWR VPWR _1504_/D sky130_fd_sc_hd__o211a_1
X_1168_ _1168_/A _1182_/A _1182_/B VGND VGND VPWR VPWR _1168_/X sky130_fd_sc_hd__and3_1
X_1237_ hold49/A hold41/A _1277_/S VGND VGND VPWR VPWR _1237_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _1022_/A _1138_/A VGND VGND VPWR VPWR _1120_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0806_ _0823_/A1 _1597_/Q _0792_/Y _0792_/A _1063_/A1 VGND VGND VPWR VPWR _0807_/B
+ sky130_fd_sc_hd__a32o_1
X_0737_ hold13/X VGND VGND VPWR VPWR _1109_/A sky130_fd_sc_hd__inv_2
X_1324__18 clkload11/A VGND VGND VPWR VPWR _1467_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
X_1571_ _1571_/CLK _1571_/D VGND VGND VPWR VPWR _1571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1005_ _1071_/A _1289_/C VGND VGND VPWR VPWR _1005_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1485_ _1485_/CLK _1485_/D VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_2
X_1554_ _1554_/CLK _1554_/D VGND VGND VPWR VPWR _1554_/Q sky130_fd_sc_hd__dfxtp_1
.ends

