VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 35.840 ;
  OBS
      LAYER met1 ;
        RECT 0.000 35.000 35.840 35.840 ;
        RECT 0.000 34.720 4.760 35.000 ;
      LAYER met1 ;
        RECT 4.760 34.720 7.840 35.000 ;
      LAYER met1 ;
        RECT 7.840 34.720 12.040 35.000 ;
      LAYER met1 ;
        RECT 12.040 34.720 13.720 35.000 ;
      LAYER met1 ;
        RECT 13.720 34.720 17.920 35.000 ;
      LAYER met1 ;
        RECT 17.920 34.720 21.000 35.000 ;
      LAYER met1 ;
        RECT 21.000 34.720 23.800 35.000 ;
      LAYER met1 ;
        RECT 23.800 34.720 28.280 35.000 ;
      LAYER met1 ;
        RECT 0.000 33.600 4.480 34.720 ;
      LAYER met1 ;
        RECT 4.480 33.880 7.840 34.720 ;
      LAYER met1 ;
        RECT 7.840 33.880 11.760 34.720 ;
      LAYER met1 ;
        RECT 4.480 33.600 8.120 33.880 ;
      LAYER met1 ;
        RECT 8.120 33.600 11.760 33.880 ;
      LAYER met1 ;
        RECT 11.760 33.600 13.720 34.720 ;
      LAYER met1 ;
        RECT 13.720 33.600 17.640 34.720 ;
      LAYER met1 ;
        RECT 17.640 33.880 21.000 34.720 ;
      LAYER met1 ;
        RECT 21.000 33.880 23.520 34.720 ;
      LAYER met1 ;
        RECT 17.640 33.600 21.280 33.880 ;
      LAYER met1 ;
        RECT 21.280 33.600 23.520 33.880 ;
        RECT 0.000 32.480 3.920 33.600 ;
      LAYER met1 ;
        RECT 3.920 33.320 8.400 33.600 ;
      LAYER met1 ;
        RECT 8.400 33.320 11.480 33.600 ;
      LAYER met1 ;
        RECT 11.480 33.320 14.280 33.600 ;
      LAYER met1 ;
        RECT 14.280 33.320 17.080 33.600 ;
      LAYER met1 ;
        RECT 17.080 33.320 21.560 33.600 ;
      LAYER met1 ;
        RECT 21.560 33.320 23.520 33.600 ;
      LAYER met1 ;
        RECT 3.920 33.040 8.680 33.320 ;
        RECT 3.920 32.480 5.040 33.040 ;
      LAYER met1 ;
        RECT 5.040 32.480 6.720 33.040 ;
        RECT 0.000 32.200 4.200 32.480 ;
      LAYER met1 ;
        RECT 4.200 32.200 4.480 32.480 ;
      LAYER met1 ;
        RECT 4.480 32.200 6.720 32.480 ;
        RECT 0.000 30.800 6.720 32.200 ;
      LAYER met1 ;
        RECT 6.720 31.080 8.680 33.040 ;
      LAYER met1 ;
        RECT 8.680 32.200 11.200 33.320 ;
      LAYER met1 ;
        RECT 11.200 33.040 14.560 33.320 ;
        RECT 11.200 32.200 12.320 33.040 ;
      LAYER met1 ;
        RECT 12.320 32.760 13.160 33.040 ;
      LAYER met1 ;
        RECT 13.160 32.760 14.560 33.040 ;
      LAYER met1 ;
        RECT 14.560 32.760 17.080 33.320 ;
      LAYER met1 ;
        RECT 17.080 33.040 21.840 33.320 ;
      LAYER met1 ;
        RECT 8.680 31.920 10.640 32.200 ;
      LAYER met1 ;
        RECT 10.640 31.920 12.320 32.200 ;
      LAYER met1 ;
        RECT 8.680 31.080 10.360 31.920 ;
      LAYER met1 ;
        RECT 6.720 30.800 8.400 31.080 ;
      LAYER met1 ;
        RECT 8.400 30.800 10.360 31.080 ;
        RECT 0.000 30.520 6.440 30.800 ;
      LAYER met1 ;
        RECT 6.440 30.520 8.120 30.800 ;
      LAYER met1 ;
        RECT 8.120 30.520 10.360 30.800 ;
        RECT 0.000 30.240 6.160 30.520 ;
      LAYER met1 ;
        RECT 6.160 30.240 7.840 30.520 ;
      LAYER met1 ;
        RECT 0.000 29.960 5.880 30.240 ;
      LAYER met1 ;
        RECT 5.880 29.960 7.840 30.240 ;
      LAYER met1 ;
        RECT 0.000 29.680 5.600 29.960 ;
      LAYER met1 ;
        RECT 5.600 29.680 7.840 29.960 ;
      LAYER met1 ;
        RECT 0.000 28.560 5.320 29.680 ;
      LAYER met1 ;
        RECT 5.320 29.400 7.840 29.680 ;
      LAYER met1 ;
        RECT 7.840 29.400 10.360 30.520 ;
      LAYER met1 ;
        RECT 5.320 28.840 7.280 29.400 ;
      LAYER met1 ;
        RECT 7.280 28.840 10.360 29.400 ;
      LAYER met1 ;
        RECT 10.360 28.840 12.320 31.920 ;
        RECT 5.320 28.560 7.000 28.840 ;
      LAYER met1 ;
        RECT 7.000 28.560 10.640 28.840 ;
      LAYER met1 ;
        RECT 10.640 28.560 12.320 28.840 ;
      LAYER met1 ;
        RECT 0.000 28.280 5.040 28.560 ;
      LAYER met1 ;
        RECT 5.040 28.280 6.440 28.560 ;
      LAYER met1 ;
        RECT 6.440 28.280 10.920 28.560 ;
      LAYER met1 ;
        RECT 10.920 28.280 12.320 28.560 ;
      LAYER met1 ;
        RECT 0.000 27.160 4.480 28.280 ;
      LAYER met1 ;
        RECT 4.480 27.160 6.440 28.280 ;
      LAYER met1 ;
        RECT 6.440 27.720 11.200 28.280 ;
      LAYER met1 ;
        RECT 11.200 27.720 12.320 28.280 ;
      LAYER met1 ;
        RECT 12.320 28.000 13.440 32.760 ;
      LAYER met1 ;
        RECT 13.440 28.000 15.120 32.760 ;
      LAYER met1 ;
        RECT 15.120 32.480 17.080 32.760 ;
      LAYER met1 ;
        RECT 17.080 32.480 18.200 33.040 ;
      LAYER met1 ;
        RECT 18.200 32.480 19.880 33.040 ;
        RECT 15.120 32.200 17.360 32.480 ;
      LAYER met1 ;
        RECT 17.360 32.200 17.640 32.480 ;
      LAYER met1 ;
        RECT 17.640 32.200 19.880 32.480 ;
        RECT 15.120 30.800 19.880 32.200 ;
      LAYER met1 ;
        RECT 19.880 31.080 21.840 33.040 ;
      LAYER met1 ;
        RECT 21.840 31.080 23.520 33.320 ;
      LAYER met1 ;
        RECT 23.520 33.040 28.280 34.720 ;
      LAYER met1 ;
        RECT 28.280 33.040 35.840 35.000 ;
      LAYER met1 ;
        RECT 23.520 32.200 25.480 33.040 ;
      LAYER met1 ;
        RECT 25.480 32.200 35.840 33.040 ;
      LAYER met1 ;
        RECT 23.520 31.920 25.760 32.200 ;
      LAYER met1 ;
        RECT 25.760 31.920 35.840 32.200 ;
      LAYER met1 ;
        RECT 23.520 31.360 27.720 31.920 ;
      LAYER met1 ;
        RECT 27.720 31.360 35.840 31.920 ;
      LAYER met1 ;
        RECT 19.880 30.800 21.560 31.080 ;
      LAYER met1 ;
        RECT 21.560 30.800 23.520 31.080 ;
        RECT 15.120 30.520 19.600 30.800 ;
      LAYER met1 ;
        RECT 19.600 30.520 21.280 30.800 ;
      LAYER met1 ;
        RECT 21.280 30.520 23.520 30.800 ;
        RECT 15.120 30.240 19.320 30.520 ;
      LAYER met1 ;
        RECT 19.320 30.240 21.000 30.520 ;
      LAYER met1 ;
        RECT 15.120 29.960 19.040 30.240 ;
      LAYER met1 ;
        RECT 19.040 29.960 21.000 30.240 ;
      LAYER met1 ;
        RECT 15.120 29.680 18.760 29.960 ;
      LAYER met1 ;
        RECT 18.760 29.680 21.000 29.960 ;
      LAYER met1 ;
        RECT 21.000 29.680 23.520 30.520 ;
      LAYER met1 ;
        RECT 23.520 30.240 28.280 31.360 ;
        RECT 23.520 29.960 25.760 30.240 ;
      LAYER met1 ;
        RECT 25.760 29.960 26.040 30.240 ;
      LAYER met1 ;
        RECT 26.040 29.960 28.280 30.240 ;
        RECT 23.520 29.680 25.480 29.960 ;
      LAYER met1 ;
        RECT 25.480 29.680 26.320 29.960 ;
      LAYER met1 ;
        RECT 26.320 29.680 28.280 29.960 ;
      LAYER met1 ;
        RECT 15.120 28.560 18.480 29.680 ;
      LAYER met1 ;
        RECT 18.480 29.400 21.000 29.680 ;
      LAYER met1 ;
        RECT 21.000 29.400 23.800 29.680 ;
      LAYER met1 ;
        RECT 23.800 29.400 25.200 29.680 ;
      LAYER met1 ;
        RECT 25.200 29.400 26.600 29.680 ;
      LAYER met1 ;
        RECT 26.600 29.400 28.280 29.680 ;
        RECT 18.480 28.840 20.440 29.400 ;
      LAYER met1 ;
        RECT 20.440 28.840 27.160 29.400 ;
      LAYER met1 ;
        RECT 18.480 28.560 20.160 28.840 ;
      LAYER met1 ;
        RECT 20.160 28.560 27.160 28.840 ;
      LAYER met1 ;
        RECT 27.160 28.560 28.280 29.400 ;
      LAYER met1 ;
        RECT 15.120 28.280 18.200 28.560 ;
      LAYER met1 ;
        RECT 18.200 28.280 19.600 28.560 ;
      LAYER met1 ;
        RECT 19.600 28.280 26.880 28.560 ;
      LAYER met1 ;
        RECT 26.880 28.280 28.280 28.560 ;
      LAYER met1 ;
        RECT 15.120 28.000 17.640 28.280 ;
        RECT 12.320 27.720 13.160 28.000 ;
      LAYER met1 ;
        RECT 13.160 27.720 14.840 28.000 ;
      LAYER met1 ;
        RECT 14.840 27.720 17.640 28.000 ;
        RECT 6.440 27.160 7.560 27.720 ;
      LAYER met1 ;
        RECT 7.560 27.440 8.400 27.720 ;
      LAYER met1 ;
        RECT 8.400 27.440 11.200 27.720 ;
      LAYER met1 ;
        RECT 7.560 27.160 8.680 27.440 ;
      LAYER met1 ;
        RECT 8.680 27.160 11.200 27.440 ;
      LAYER met1 ;
        RECT 11.200 27.160 14.560 27.720 ;
      LAYER met1 ;
        RECT 14.560 27.160 17.640 27.720 ;
      LAYER met1 ;
        RECT 17.640 27.160 19.600 28.280 ;
      LAYER met1 ;
        RECT 19.600 27.720 23.520 28.280 ;
      LAYER met1 ;
        RECT 23.520 28.000 24.640 28.280 ;
      LAYER met1 ;
        RECT 24.640 28.000 26.600 28.280 ;
      LAYER met1 ;
        RECT 23.520 27.720 24.920 28.000 ;
      LAYER met1 ;
        RECT 24.920 27.720 26.600 28.000 ;
        RECT 19.600 27.160 20.720 27.720 ;
      LAYER met1 ;
        RECT 20.720 27.440 21.560 27.720 ;
      LAYER met1 ;
        RECT 21.560 27.440 23.520 27.720 ;
      LAYER met1 ;
        RECT 23.520 27.440 25.200 27.720 ;
      LAYER met1 ;
        RECT 25.200 27.440 26.600 27.720 ;
      LAYER met1 ;
        RECT 20.720 27.160 21.840 27.440 ;
      LAYER met1 ;
        RECT 21.840 27.160 23.800 27.440 ;
      LAYER met1 ;
        RECT 23.800 27.160 25.480 27.440 ;
      LAYER met1 ;
        RECT 25.480 27.160 26.600 27.440 ;
      LAYER met1 ;
        RECT 26.600 27.160 28.280 28.280 ;
      LAYER met1 ;
        RECT 28.280 27.160 35.840 31.360 ;
        RECT 0.000 26.880 4.200 27.160 ;
      LAYER met1 ;
        RECT 4.200 26.880 6.720 27.160 ;
      LAYER met1 ;
        RECT 6.720 26.880 7.280 27.160 ;
      LAYER met1 ;
        RECT 7.280 26.880 8.680 27.160 ;
      LAYER met1 ;
        RECT 0.000 25.760 3.920 26.880 ;
      LAYER met1 ;
        RECT 3.920 26.040 8.680 26.880 ;
      LAYER met1 ;
        RECT 8.680 26.040 11.760 27.160 ;
      LAYER met1 ;
        RECT 11.760 26.600 14.560 27.160 ;
      LAYER met1 ;
        RECT 14.560 26.880 17.360 27.160 ;
      LAYER met1 ;
        RECT 17.360 26.880 19.880 27.160 ;
      LAYER met1 ;
        RECT 19.880 26.880 20.440 27.160 ;
      LAYER met1 ;
        RECT 20.440 26.880 21.840 27.160 ;
      LAYER met1 ;
        RECT 21.840 26.880 24.080 27.160 ;
      LAYER met1 ;
        RECT 24.080 26.880 25.760 27.160 ;
      LAYER met1 ;
        RECT 25.760 26.880 26.320 27.160 ;
      LAYER met1 ;
        RECT 26.320 26.880 27.720 27.160 ;
      LAYER met1 ;
        RECT 14.560 26.600 17.080 26.880 ;
      LAYER met1 ;
        RECT 11.760 26.320 14.280 26.600 ;
      LAYER met1 ;
        RECT 14.280 26.320 17.080 26.600 ;
      LAYER met1 ;
        RECT 11.760 26.040 13.720 26.320 ;
        RECT 3.920 25.760 8.400 26.040 ;
      LAYER met1 ;
        RECT 8.400 25.760 12.040 26.040 ;
      LAYER met1 ;
        RECT 12.040 25.760 13.720 26.040 ;
      LAYER met1 ;
        RECT 13.720 25.760 17.080 26.320 ;
      LAYER met1 ;
        RECT 17.080 26.040 21.840 26.880 ;
      LAYER met1 ;
        RECT 21.840 26.040 24.360 26.880 ;
      LAYER met1 ;
        RECT 24.360 26.040 27.720 26.880 ;
      LAYER met1 ;
        RECT 27.720 26.040 35.840 27.160 ;
      LAYER met1 ;
        RECT 17.080 25.760 21.560 26.040 ;
      LAYER met1 ;
        RECT 21.560 25.760 24.360 26.040 ;
      LAYER met1 ;
        RECT 24.360 25.760 27.440 26.040 ;
      LAYER met1 ;
        RECT 27.440 25.760 35.840 26.040 ;
        RECT 0.000 24.640 35.840 25.760 ;
        RECT 0.000 22.960 3.080 24.640 ;
      LAYER met1 ;
        RECT 3.080 22.960 8.680 24.640 ;
      LAYER met1 ;
        RECT 8.680 24.080 11.760 24.640 ;
      LAYER met1 ;
        RECT 11.760 24.080 18.200 24.640 ;
      LAYER met1 ;
        RECT 0.000 22.680 3.360 22.960 ;
      LAYER met1 ;
        RECT 3.360 22.680 8.680 22.960 ;
      LAYER met1 ;
        RECT 8.680 22.680 11.200 24.080 ;
      LAYER met1 ;
        RECT 11.200 22.960 18.200 24.080 ;
        RECT 11.200 22.680 14.280 22.960 ;
      LAYER met1 ;
        RECT 14.280 22.680 15.680 22.960 ;
      LAYER met1 ;
        RECT 15.680 22.680 18.200 22.960 ;
      LAYER met1 ;
        RECT 18.200 22.680 19.880 24.640 ;
        RECT 0.000 22.400 3.640 22.680 ;
      LAYER met1 ;
        RECT 3.640 22.400 8.680 22.680 ;
      LAYER met1 ;
        RECT 8.680 22.400 10.640 22.680 ;
      LAYER met1 ;
        RECT 10.640 22.400 13.720 22.680 ;
      LAYER met1 ;
        RECT 0.000 22.120 3.920 22.400 ;
      LAYER met1 ;
        RECT 3.920 22.120 8.680 22.400 ;
      LAYER met1 ;
        RECT 8.680 22.120 10.360 22.400 ;
      LAYER met1 ;
        RECT 10.360 22.120 13.720 22.400 ;
      LAYER met1 ;
        RECT 13.720 22.120 16.240 22.680 ;
      LAYER met1 ;
        RECT 16.240 22.400 18.480 22.680 ;
      LAYER met1 ;
        RECT 18.480 22.400 19.880 22.680 ;
        RECT 0.000 21.840 4.200 22.120 ;
      LAYER met1 ;
        RECT 4.200 21.840 7.280 22.120 ;
      LAYER met1 ;
        RECT 0.000 15.120 4.480 21.840 ;
        RECT 0.000 13.440 0.840 15.120 ;
      LAYER met1 ;
        RECT 0.840 14.280 3.360 15.120 ;
      LAYER met1 ;
        RECT 3.360 14.280 4.480 15.120 ;
      LAYER met1 ;
        RECT 0.840 13.720 3.640 14.280 ;
      LAYER met1 ;
        RECT 3.640 13.720 4.480 14.280 ;
      LAYER met1 ;
        RECT 4.480 13.720 7.280 21.840 ;
      LAYER met1 ;
        RECT 7.280 19.320 10.360 22.120 ;
      LAYER met1 ;
        RECT 10.360 21.560 13.160 22.120 ;
      LAYER met1 ;
        RECT 13.160 21.560 16.240 22.120 ;
      LAYER met1 ;
        RECT 10.360 20.160 12.880 21.560 ;
      LAYER met1 ;
        RECT 12.880 20.720 16.240 21.560 ;
      LAYER met1 ;
        RECT 16.240 20.720 18.760 22.400 ;
      LAYER met1 ;
        RECT 18.760 20.720 19.880 22.400 ;
        RECT 12.880 20.160 19.880 20.720 ;
      LAYER met1 ;
        RECT 10.360 19.600 13.160 20.160 ;
      LAYER met1 ;
        RECT 13.160 19.600 19.880 20.160 ;
      LAYER met1 ;
        RECT 10.360 19.320 13.720 19.600 ;
      LAYER met1 ;
        RECT 7.280 19.040 10.640 19.320 ;
      LAYER met1 ;
        RECT 10.640 19.040 13.720 19.320 ;
      LAYER met1 ;
        RECT 13.720 19.040 16.240 19.600 ;
      LAYER met1 ;
        RECT 16.240 19.040 17.360 19.600 ;
      LAYER met1 ;
        RECT 17.360 19.040 19.880 19.600 ;
      LAYER met1 ;
        RECT 19.880 19.320 22.400 24.640 ;
      LAYER met1 ;
        RECT 22.400 23.520 25.760 24.640 ;
      LAYER met1 ;
        RECT 25.760 23.520 28.280 24.640 ;
      LAYER met1 ;
        RECT 22.400 23.240 25.480 23.520 ;
      LAYER met1 ;
        RECT 25.480 23.240 28.280 23.520 ;
      LAYER met1 ;
        RECT 22.400 22.960 25.200 23.240 ;
      LAYER met1 ;
        RECT 25.200 22.960 28.280 23.240 ;
      LAYER met1 ;
        RECT 28.280 22.960 35.840 24.640 ;
        RECT 22.400 21.280 24.920 22.960 ;
      LAYER met1 ;
        RECT 24.920 22.680 28.000 22.960 ;
      LAYER met1 ;
        RECT 28.000 22.680 35.840 22.960 ;
      LAYER met1 ;
        RECT 24.920 21.280 27.720 22.680 ;
      LAYER met1 ;
        RECT 22.400 21.000 24.640 21.280 ;
      LAYER met1 ;
        RECT 24.640 21.000 27.720 21.280 ;
      LAYER met1 ;
        RECT 22.400 19.320 23.520 21.000 ;
      LAYER met1 ;
        RECT 23.520 20.720 27.720 21.000 ;
      LAYER met1 ;
        RECT 27.720 20.720 35.840 22.680 ;
      LAYER met1 ;
        RECT 23.520 20.440 26.600 20.720 ;
      LAYER met1 ;
        RECT 26.600 20.440 35.840 20.720 ;
      LAYER met1 ;
        RECT 23.520 20.160 26.320 20.440 ;
      LAYER met1 ;
        RECT 26.320 20.160 35.840 20.440 ;
      LAYER met1 ;
        RECT 19.880 19.040 22.680 19.320 ;
      LAYER met1 ;
        RECT 22.680 19.040 23.520 19.320 ;
      LAYER met1 ;
        RECT 23.520 19.040 26.040 20.160 ;
      LAYER met1 ;
        RECT 7.280 18.760 10.920 19.040 ;
      LAYER met1 ;
        RECT 10.920 18.760 14.000 19.040 ;
      LAYER met1 ;
        RECT 14.000 18.760 15.960 19.040 ;
      LAYER met1 ;
        RECT 15.960 18.760 17.640 19.040 ;
      LAYER met1 ;
        RECT 17.640 18.760 19.880 19.040 ;
      LAYER met1 ;
        RECT 19.880 18.760 22.960 19.040 ;
      LAYER met1 ;
        RECT 22.960 18.760 23.240 19.040 ;
      LAYER met1 ;
        RECT 23.240 18.760 26.040 19.040 ;
      LAYER met1 ;
        RECT 7.280 17.640 11.200 18.760 ;
      LAYER met1 ;
        RECT 11.200 17.640 18.200 18.760 ;
      LAYER met1 ;
        RECT 18.200 17.640 19.880 18.760 ;
      LAYER met1 ;
        RECT 19.880 18.480 26.040 18.760 ;
      LAYER met1 ;
        RECT 26.040 18.480 35.840 20.160 ;
      LAYER met1 ;
        RECT 19.880 18.200 24.920 18.480 ;
      LAYER met1 ;
        RECT 24.920 18.200 35.840 18.480 ;
      LAYER met1 ;
        RECT 19.880 17.640 24.640 18.200 ;
      LAYER met1 ;
        RECT 24.640 17.640 35.840 18.200 ;
        RECT 7.280 17.080 11.760 17.640 ;
      LAYER met1 ;
        RECT 11.760 17.360 18.480 17.640 ;
      LAYER met1 ;
        RECT 18.480 17.360 19.880 17.640 ;
      LAYER met1 ;
        RECT 19.880 17.360 24.920 17.640 ;
      LAYER met1 ;
        RECT 24.920 17.360 35.840 17.640 ;
      LAYER met1 ;
        RECT 11.760 17.080 18.760 17.360 ;
      LAYER met1 ;
        RECT 7.280 16.800 15.960 17.080 ;
      LAYER met1 ;
        RECT 15.960 16.800 18.760 17.080 ;
      LAYER met1 ;
        RECT 7.280 15.120 16.240 16.800 ;
        RECT 7.280 13.720 10.360 15.120 ;
      LAYER met1 ;
        RECT 10.360 14.280 12.880 15.120 ;
      LAYER met1 ;
        RECT 12.880 14.280 16.240 15.120 ;
      LAYER met1 ;
        RECT 10.360 13.720 13.160 14.280 ;
      LAYER met1 ;
        RECT 13.160 14.000 16.240 14.280 ;
      LAYER met1 ;
        RECT 16.240 14.000 18.760 16.800 ;
      LAYER met1 ;
        RECT 13.160 13.720 15.960 14.000 ;
      LAYER met1 ;
        RECT 15.960 13.720 18.760 14.000 ;
        RECT 0.840 13.440 7.000 13.720 ;
      LAYER met1 ;
        RECT 7.000 13.440 10.360 13.720 ;
      LAYER met1 ;
        RECT 10.360 13.440 18.760 13.720 ;
      LAYER met1 ;
        RECT 18.760 13.440 19.880 17.360 ;
      LAYER met1 ;
        RECT 19.880 17.080 26.040 17.360 ;
        RECT 19.880 16.800 22.960 17.080 ;
      LAYER met1 ;
        RECT 22.960 16.800 23.240 17.080 ;
      LAYER met1 ;
        RECT 23.240 16.800 26.040 17.080 ;
        RECT 19.880 16.520 22.680 16.800 ;
      LAYER met1 ;
        RECT 22.680 16.520 23.520 16.800 ;
        RECT 0.000 13.160 1.120 13.440 ;
      LAYER met1 ;
        RECT 1.120 13.160 6.720 13.440 ;
      LAYER met1 ;
        RECT 6.720 13.160 10.640 13.440 ;
      LAYER met1 ;
        RECT 10.640 13.160 18.480 13.440 ;
      LAYER met1 ;
        RECT 18.480 13.160 19.880 13.440 ;
        RECT 0.000 12.040 1.680 13.160 ;
      LAYER met1 ;
        RECT 1.680 12.040 6.440 13.160 ;
      LAYER met1 ;
        RECT 0.000 11.760 1.960 12.040 ;
      LAYER met1 ;
        RECT 1.960 11.760 6.440 12.040 ;
      LAYER met1 ;
        RECT 6.440 11.760 11.200 13.160 ;
      LAYER met1 ;
        RECT 11.200 11.760 18.200 13.160 ;
      LAYER met1 ;
        RECT 0.000 11.480 2.240 11.760 ;
      LAYER met1 ;
        RECT 2.240 11.480 6.440 11.760 ;
      LAYER met1 ;
        RECT 0.000 11.200 2.520 11.480 ;
      LAYER met1 ;
        RECT 2.520 11.200 6.440 11.480 ;
      LAYER met1 ;
        RECT 6.440 11.200 11.760 11.760 ;
      LAYER met1 ;
        RECT 11.760 11.200 18.200 11.760 ;
      LAYER met1 ;
        RECT 18.200 11.200 19.880 13.160 ;
      LAYER met1 ;
        RECT 19.880 11.200 22.400 16.520 ;
      LAYER met1 ;
        RECT 22.400 14.840 23.520 16.520 ;
      LAYER met1 ;
        RECT 23.520 15.680 26.040 16.800 ;
      LAYER met1 ;
        RECT 26.040 15.680 35.840 17.360 ;
      LAYER met1 ;
        RECT 23.520 15.400 26.320 15.680 ;
      LAYER met1 ;
        RECT 26.320 15.400 35.840 15.680 ;
      LAYER met1 ;
        RECT 23.520 15.120 26.600 15.400 ;
      LAYER met1 ;
        RECT 26.600 15.120 35.840 15.400 ;
      LAYER met1 ;
        RECT 23.520 14.840 27.720 15.120 ;
      LAYER met1 ;
        RECT 22.400 14.560 24.640 14.840 ;
      LAYER met1 ;
        RECT 24.640 14.560 27.720 14.840 ;
      LAYER met1 ;
        RECT 22.400 13.440 24.920 14.560 ;
      LAYER met1 ;
        RECT 24.920 14.000 27.720 14.560 ;
      LAYER met1 ;
        RECT 27.720 14.000 35.840 15.120 ;
      LAYER met1 ;
        RECT 24.920 13.720 28.000 14.000 ;
      LAYER met1 ;
        RECT 28.000 13.720 35.840 14.000 ;
      LAYER met1 ;
        RECT 24.920 13.440 28.280 13.720 ;
      LAYER met1 ;
        RECT 22.400 13.160 25.480 13.440 ;
      LAYER met1 ;
        RECT 25.480 13.160 28.280 13.440 ;
      LAYER met1 ;
        RECT 22.400 11.200 25.760 13.160 ;
      LAYER met1 ;
        RECT 25.760 11.200 28.280 13.160 ;
      LAYER met1 ;
        RECT 28.280 11.200 35.840 13.720 ;
        RECT 0.000 10.080 35.840 11.200 ;
        RECT 0.000 8.400 3.080 10.080 ;
      LAYER met1 ;
        RECT 3.080 9.520 7.840 10.080 ;
      LAYER met1 ;
        RECT 7.840 9.520 9.800 10.080 ;
      LAYER met1 ;
        RECT 9.800 9.800 14.280 10.080 ;
      LAYER met1 ;
        RECT 14.280 9.800 18.480 10.080 ;
      LAYER met1 ;
        RECT 9.800 9.520 14.560 9.800 ;
      LAYER met1 ;
        RECT 14.560 9.520 18.480 9.800 ;
      LAYER met1 ;
        RECT 18.480 9.520 19.600 10.080 ;
        RECT 3.080 8.960 8.400 9.520 ;
      LAYER met1 ;
        RECT 8.400 8.960 9.800 9.520 ;
      LAYER met1 ;
        RECT 9.800 9.240 14.840 9.520 ;
      LAYER met1 ;
        RECT 14.840 9.240 17.920 9.520 ;
      LAYER met1 ;
        RECT 17.920 9.240 19.600 9.520 ;
        RECT 9.800 8.960 15.120 9.240 ;
      LAYER met1 ;
        RECT 15.120 8.960 17.640 9.240 ;
      LAYER met1 ;
        RECT 3.080 8.680 8.120 8.960 ;
      LAYER met1 ;
        RECT 8.120 8.680 9.800 8.960 ;
      LAYER met1 ;
        RECT 9.800 8.680 14.840 8.960 ;
      LAYER met1 ;
        RECT 14.840 8.680 17.640 8.960 ;
      LAYER met1 ;
        RECT 17.640 8.680 19.600 9.240 ;
      LAYER met1 ;
        RECT 19.600 8.960 24.360 10.080 ;
      LAYER met1 ;
        RECT 24.360 8.960 26.040 10.080 ;
      LAYER met1 ;
        RECT 26.040 8.960 35.840 10.080 ;
        RECT 19.600 8.680 24.080 8.960 ;
      LAYER met1 ;
        RECT 24.080 8.680 26.320 8.960 ;
      LAYER met1 ;
        RECT 26.320 8.680 35.840 8.960 ;
      LAYER met1 ;
        RECT 3.080 8.400 7.840 8.680 ;
      LAYER met1 ;
        RECT 7.840 8.400 9.800 8.680 ;
      LAYER met1 ;
        RECT 9.800 8.400 14.560 8.680 ;
      LAYER met1 ;
        RECT 14.560 8.400 17.080 8.680 ;
        RECT 0.000 8.120 3.360 8.400 ;
      LAYER met1 ;
        RECT 3.360 8.120 7.560 8.400 ;
      LAYER met1 ;
        RECT 7.560 8.120 9.800 8.400 ;
      LAYER met1 ;
        RECT 9.800 8.120 14.280 8.400 ;
      LAYER met1 ;
        RECT 14.280 8.120 17.080 8.400 ;
        RECT 0.000 1.120 4.480 8.120 ;
      LAYER met1 ;
        RECT 4.480 1.120 6.440 8.120 ;
      LAYER met1 ;
        RECT 6.440 7.840 10.920 8.120 ;
      LAYER met1 ;
        RECT 10.920 7.840 13.160 8.120 ;
      LAYER met1 ;
        RECT 13.160 7.840 17.080 8.120 ;
        RECT 6.440 1.120 11.200 7.840 ;
        RECT 0.000 0.840 4.760 1.120 ;
      LAYER met1 ;
        RECT 4.760 0.840 6.160 1.120 ;
      LAYER met1 ;
        RECT 6.160 0.840 11.200 1.120 ;
      LAYER met1 ;
        RECT 11.200 0.840 12.880 7.840 ;
      LAYER met1 ;
        RECT 12.880 7.560 17.080 7.840 ;
      LAYER met1 ;
        RECT 17.080 7.560 19.600 8.680 ;
      LAYER met1 ;
        RECT 19.600 8.400 23.800 8.680 ;
      LAYER met1 ;
        RECT 23.800 8.400 26.880 8.680 ;
      LAYER met1 ;
        RECT 12.880 7.280 17.360 7.560 ;
      LAYER met1 ;
        RECT 17.360 7.280 19.600 7.560 ;
      LAYER met1 ;
        RECT 19.600 7.280 23.520 8.400 ;
      LAYER met1 ;
        RECT 23.520 8.120 26.880 8.400 ;
      LAYER met1 ;
        RECT 26.880 8.120 35.840 8.680 ;
      LAYER met1 ;
        RECT 23.520 7.840 24.920 8.120 ;
      LAYER met1 ;
        RECT 24.920 7.840 25.760 8.120 ;
      LAYER met1 ;
        RECT 25.760 7.840 27.160 8.120 ;
      LAYER met1 ;
        RECT 27.160 7.840 35.840 8.120 ;
      LAYER met1 ;
        RECT 23.520 7.280 24.640 7.840 ;
      LAYER met1 ;
        RECT 12.880 2.800 17.640 7.280 ;
      LAYER met1 ;
        RECT 17.640 3.080 19.600 7.280 ;
      LAYER met1 ;
        RECT 19.600 3.920 22.960 7.280 ;
      LAYER met1 ;
        RECT 22.960 3.920 24.640 7.280 ;
      LAYER met1 ;
        RECT 19.600 3.640 23.240 3.920 ;
      LAYER met1 ;
        RECT 23.240 3.640 24.640 3.920 ;
      LAYER met1 ;
        RECT 19.600 3.080 23.520 3.640 ;
      LAYER met1 ;
        RECT 23.520 3.080 24.640 3.640 ;
      LAYER met1 ;
        RECT 24.640 3.080 25.760 7.840 ;
      LAYER met1 ;
        RECT 25.760 7.560 27.440 7.840 ;
      LAYER met1 ;
        RECT 27.440 7.560 35.840 7.840 ;
      LAYER met1 ;
        RECT 25.760 3.360 27.720 7.560 ;
      LAYER met1 ;
        RECT 27.720 3.360 35.840 7.560 ;
      LAYER met1 ;
        RECT 25.760 3.080 27.440 3.360 ;
      LAYER met1 ;
        RECT 27.440 3.080 35.840 3.360 ;
      LAYER met1 ;
        RECT 17.640 2.800 19.880 3.080 ;
      LAYER met1 ;
        RECT 19.880 2.800 23.520 3.080 ;
      LAYER met1 ;
        RECT 23.520 2.800 24.920 3.080 ;
      LAYER met1 ;
        RECT 24.920 2.800 25.760 3.080 ;
      LAYER met1 ;
        RECT 25.760 2.800 27.160 3.080 ;
      LAYER met1 ;
        RECT 27.160 2.800 35.840 3.080 ;
        RECT 12.880 0.840 17.080 2.800 ;
      LAYER met1 ;
        RECT 17.080 2.520 20.160 2.800 ;
      LAYER met1 ;
        RECT 20.160 2.520 23.520 2.800 ;
      LAYER met1 ;
        RECT 23.520 2.520 26.880 2.800 ;
        RECT 17.080 2.240 20.440 2.520 ;
      LAYER met1 ;
        RECT 20.440 2.240 23.800 2.520 ;
      LAYER met1 ;
        RECT 23.800 2.240 26.880 2.520 ;
        RECT 17.080 1.960 20.720 2.240 ;
      LAYER met1 ;
        RECT 20.720 1.960 24.080 2.240 ;
      LAYER met1 ;
        RECT 24.080 1.960 26.880 2.240 ;
        RECT 17.080 0.840 21.000 1.960 ;
      LAYER met1 ;
        RECT 21.000 0.840 24.360 1.960 ;
      LAYER met1 ;
        RECT 24.360 1.680 26.880 1.960 ;
      LAYER met1 ;
        RECT 26.880 1.680 35.840 2.800 ;
      LAYER met1 ;
        RECT 24.360 1.400 26.600 1.680 ;
      LAYER met1 ;
        RECT 26.600 1.400 35.840 1.680 ;
      LAYER met1 ;
        RECT 24.360 1.120 26.320 1.400 ;
      LAYER met1 ;
        RECT 26.320 1.120 35.840 1.400 ;
      LAYER met1 ;
        RECT 24.360 0.840 26.040 1.120 ;
      LAYER met1 ;
        RECT 26.040 0.840 35.840 1.120 ;
        RECT 0.000 0.000 35.840 0.840 ;
      LAYER met2 ;
        RECT 4.760 34.720 7.840 35.000 ;
        RECT 12.040 34.720 13.720 35.000 ;
        RECT 17.920 34.720 21.000 35.000 ;
        RECT 23.800 34.720 28.280 35.000 ;
        RECT 4.480 33.880 7.840 34.720 ;
        RECT 4.480 33.600 8.120 33.880 ;
        RECT 11.760 33.600 13.720 34.720 ;
        RECT 17.640 33.880 21.000 34.720 ;
        RECT 17.640 33.600 21.280 33.880 ;
        RECT 3.920 33.320 8.400 33.600 ;
        RECT 11.480 33.320 14.280 33.600 ;
        RECT 17.080 33.320 21.560 33.600 ;
        RECT 3.920 33.040 8.680 33.320 ;
        RECT 3.920 32.480 5.040 33.040 ;
        RECT 4.200 32.200 4.480 32.480 ;
        RECT 6.720 31.080 8.680 33.040 ;
        RECT 11.200 33.040 14.560 33.320 ;
        RECT 11.200 32.200 12.320 33.040 ;
        RECT 13.160 32.760 14.560 33.040 ;
        RECT 17.080 33.040 21.840 33.320 ;
        RECT 10.640 31.920 12.320 32.200 ;
        RECT 6.720 30.800 8.400 31.080 ;
        RECT 6.440 30.520 8.120 30.800 ;
        RECT 6.160 30.240 7.840 30.520 ;
        RECT 5.880 29.960 7.840 30.240 ;
        RECT 5.600 29.680 7.840 29.960 ;
        RECT 5.320 29.400 7.840 29.680 ;
        RECT 5.320 28.840 7.280 29.400 ;
        RECT 10.360 28.840 12.320 31.920 ;
        RECT 5.320 28.560 7.000 28.840 ;
        RECT 10.640 28.560 12.320 28.840 ;
        RECT 5.040 28.280 6.440 28.560 ;
        RECT 10.920 28.280 12.320 28.560 ;
        RECT 4.480 27.160 6.440 28.280 ;
        RECT 11.200 27.720 12.320 28.280 ;
        RECT 13.440 28.000 15.120 32.760 ;
        RECT 17.080 32.480 18.200 33.040 ;
        RECT 17.360 32.200 17.640 32.480 ;
        RECT 19.880 31.080 21.840 33.040 ;
        RECT 23.520 33.040 28.280 34.720 ;
        RECT 23.520 32.200 25.480 33.040 ;
        RECT 23.520 31.920 25.760 32.200 ;
        RECT 23.520 31.360 27.720 31.920 ;
        RECT 19.880 30.800 21.560 31.080 ;
        RECT 19.600 30.520 21.280 30.800 ;
        RECT 19.320 30.240 21.000 30.520 ;
        RECT 19.040 29.960 21.000 30.240 ;
        RECT 18.760 29.680 21.000 29.960 ;
        RECT 23.520 30.240 28.280 31.360 ;
        RECT 23.520 29.960 25.760 30.240 ;
        RECT 26.040 29.960 28.280 30.240 ;
        RECT 23.520 29.680 25.480 29.960 ;
        RECT 26.320 29.680 28.280 29.960 ;
        RECT 18.480 29.400 21.000 29.680 ;
        RECT 23.800 29.400 25.200 29.680 ;
        RECT 26.600 29.400 28.280 29.680 ;
        RECT 18.480 28.840 20.440 29.400 ;
        RECT 18.480 28.560 20.160 28.840 ;
        RECT 27.160 28.560 28.280 29.400 ;
        RECT 18.200 28.280 19.600 28.560 ;
        RECT 26.880 28.280 28.280 28.560 ;
        RECT 13.160 27.720 14.840 28.000 ;
        RECT 7.560 27.440 8.400 27.720 ;
        RECT 7.560 27.160 8.680 27.440 ;
        RECT 11.200 27.160 14.560 27.720 ;
        RECT 17.640 27.160 19.600 28.280 ;
        RECT 23.520 28.000 24.640 28.280 ;
        RECT 23.520 27.720 24.920 28.000 ;
        RECT 20.720 27.440 21.560 27.720 ;
        RECT 23.520 27.440 25.200 27.720 ;
        RECT 20.720 27.160 21.840 27.440 ;
        RECT 23.800 27.160 25.480 27.440 ;
        RECT 26.600 27.160 28.280 28.280 ;
        RECT 4.200 26.880 6.720 27.160 ;
        RECT 7.280 26.880 8.680 27.160 ;
        RECT 3.920 26.040 8.680 26.880 ;
        RECT 11.760 26.600 14.560 27.160 ;
        RECT 17.360 26.880 19.880 27.160 ;
        RECT 20.440 26.880 21.840 27.160 ;
        RECT 24.080 26.880 25.760 27.160 ;
        RECT 26.320 26.880 27.720 27.160 ;
        RECT 11.760 26.320 14.280 26.600 ;
        RECT 11.760 26.040 13.720 26.320 ;
        RECT 3.920 25.760 8.400 26.040 ;
        RECT 12.040 25.760 13.720 26.040 ;
        RECT 17.080 26.040 21.840 26.880 ;
        RECT 24.360 26.040 27.720 26.880 ;
        RECT 17.080 25.760 21.560 26.040 ;
        RECT 24.360 25.760 27.440 26.040 ;
        RECT 3.080 22.960 8.680 24.640 ;
        RECT 11.760 24.080 18.200 24.640 ;
        RECT 3.360 22.680 8.680 22.960 ;
        RECT 11.200 22.960 18.200 24.080 ;
        RECT 11.200 22.680 14.280 22.960 ;
        RECT 15.680 22.680 18.200 22.960 ;
        RECT 3.640 22.400 8.680 22.680 ;
        RECT 10.640 22.400 13.720 22.680 ;
        RECT 3.920 22.120 8.680 22.400 ;
        RECT 10.360 22.120 13.720 22.400 ;
        RECT 16.240 22.400 18.480 22.680 ;
        RECT 4.200 21.840 7.280 22.120 ;
        RECT 0.840 14.280 3.360 15.120 ;
        RECT 0.840 13.720 3.640 14.280 ;
        RECT 4.480 13.720 7.280 21.840 ;
        RECT 10.360 21.560 13.160 22.120 ;
        RECT 10.360 20.160 12.880 21.560 ;
        RECT 16.240 20.720 18.760 22.400 ;
        RECT 10.360 19.600 13.160 20.160 ;
        RECT 10.360 19.320 13.720 19.600 ;
        RECT 10.640 19.040 13.720 19.320 ;
        RECT 16.240 19.040 17.360 19.600 ;
        RECT 19.880 19.320 22.400 24.640 ;
        RECT 25.760 23.520 28.280 24.640 ;
        RECT 25.480 23.240 28.280 23.520 ;
        RECT 25.200 22.960 28.280 23.240 ;
        RECT 24.920 22.680 28.000 22.960 ;
        RECT 24.920 21.280 27.720 22.680 ;
        RECT 24.640 21.000 27.720 21.280 ;
        RECT 23.520 20.720 27.720 21.000 ;
        RECT 23.520 20.440 26.600 20.720 ;
        RECT 23.520 20.160 26.320 20.440 ;
        RECT 19.880 19.040 22.680 19.320 ;
        RECT 23.520 19.040 26.040 20.160 ;
        RECT 10.920 18.760 14.000 19.040 ;
        RECT 15.960 18.760 17.640 19.040 ;
        RECT 19.880 18.760 22.960 19.040 ;
        RECT 23.240 18.760 26.040 19.040 ;
        RECT 11.200 17.640 18.200 18.760 ;
        RECT 19.880 18.480 26.040 18.760 ;
        RECT 19.880 18.200 24.920 18.480 ;
        RECT 19.880 17.640 24.640 18.200 ;
        RECT 11.760 17.360 18.480 17.640 ;
        RECT 19.880 17.360 24.920 17.640 ;
        RECT 11.760 17.080 18.760 17.360 ;
        RECT 15.960 16.800 18.760 17.080 ;
        RECT 10.360 14.280 12.880 15.120 ;
        RECT 10.360 13.720 13.160 14.280 ;
        RECT 16.240 14.000 18.760 16.800 ;
        RECT 15.960 13.720 18.760 14.000 ;
        RECT 0.840 13.440 7.000 13.720 ;
        RECT 10.360 13.440 18.760 13.720 ;
        RECT 19.880 17.080 26.040 17.360 ;
        RECT 19.880 16.800 22.960 17.080 ;
        RECT 23.240 16.800 26.040 17.080 ;
        RECT 19.880 16.520 22.680 16.800 ;
        RECT 1.120 13.160 6.720 13.440 ;
        RECT 10.640 13.160 18.480 13.440 ;
        RECT 1.680 12.040 6.440 13.160 ;
        RECT 1.960 11.760 6.440 12.040 ;
        RECT 11.200 11.760 18.200 13.160 ;
        RECT 2.240 11.480 6.440 11.760 ;
        RECT 2.520 11.200 6.440 11.480 ;
        RECT 11.760 11.200 18.200 11.760 ;
        RECT 19.880 11.200 22.400 16.520 ;
        RECT 23.520 15.680 26.040 16.800 ;
        RECT 23.520 15.400 26.320 15.680 ;
        RECT 23.520 15.120 26.600 15.400 ;
        RECT 23.520 14.840 27.720 15.120 ;
        RECT 24.640 14.560 27.720 14.840 ;
        RECT 24.920 14.000 27.720 14.560 ;
        RECT 24.920 13.720 28.000 14.000 ;
        RECT 24.920 13.440 28.280 13.720 ;
        RECT 25.480 13.160 28.280 13.440 ;
        RECT 25.760 11.200 28.280 13.160 ;
        RECT 3.080 9.520 7.840 10.080 ;
        RECT 9.800 9.800 14.280 10.080 ;
        RECT 9.800 9.520 14.560 9.800 ;
        RECT 18.480 9.520 19.600 10.080 ;
        RECT 3.080 8.960 8.400 9.520 ;
        RECT 9.800 9.240 14.840 9.520 ;
        RECT 17.920 9.240 19.600 9.520 ;
        RECT 9.800 8.960 15.120 9.240 ;
        RECT 3.080 8.680 8.120 8.960 ;
        RECT 9.800 8.680 14.840 8.960 ;
        RECT 17.640 8.680 19.600 9.240 ;
        RECT 24.360 8.960 26.040 10.080 ;
        RECT 24.080 8.680 26.320 8.960 ;
        RECT 3.080 8.400 7.840 8.680 ;
        RECT 9.800 8.400 14.560 8.680 ;
        RECT 3.360 8.120 7.560 8.400 ;
        RECT 9.800 8.120 14.280 8.400 ;
        RECT 4.480 1.120 6.440 8.120 ;
        RECT 10.920 7.840 13.160 8.120 ;
        RECT 4.760 0.840 6.160 1.120 ;
        RECT 11.200 0.840 12.880 7.840 ;
        RECT 17.080 7.560 19.600 8.680 ;
        RECT 23.800 8.400 26.880 8.680 ;
        RECT 17.360 7.280 19.600 7.560 ;
        RECT 23.520 8.120 26.880 8.400 ;
        RECT 23.520 7.840 24.920 8.120 ;
        RECT 25.760 7.840 27.160 8.120 ;
        RECT 23.520 7.280 24.640 7.840 ;
        RECT 17.640 3.080 19.600 7.280 ;
        RECT 22.960 3.920 24.640 7.280 ;
        RECT 23.240 3.640 24.640 3.920 ;
        RECT 23.520 3.080 24.640 3.640 ;
        RECT 25.760 7.560 27.440 7.840 ;
        RECT 25.760 3.360 27.720 7.560 ;
        RECT 25.760 3.080 27.440 3.360 ;
        RECT 17.640 2.800 19.880 3.080 ;
        RECT 23.520 2.800 24.920 3.080 ;
        RECT 25.760 2.800 27.160 3.080 ;
        RECT 17.080 2.520 20.160 2.800 ;
        RECT 23.520 2.520 26.880 2.800 ;
        RECT 17.080 2.240 20.440 2.520 ;
        RECT 23.800 2.240 26.880 2.520 ;
        RECT 17.080 1.960 20.720 2.240 ;
        RECT 24.080 1.960 26.880 2.240 ;
        RECT 17.080 0.840 21.000 1.960 ;
        RECT 24.360 1.680 26.880 1.960 ;
        RECT 24.360 1.400 26.600 1.680 ;
        RECT 24.360 1.120 26.320 1.400 ;
        RECT 24.360 0.840 26.040 1.120 ;
      LAYER met3 ;
        RECT 4.760 34.720 7.840 35.000 ;
        RECT 12.040 34.720 13.720 35.000 ;
        RECT 17.920 34.720 21.000 35.000 ;
        RECT 23.800 34.720 28.280 35.000 ;
        RECT 4.480 33.880 7.840 34.720 ;
        RECT 4.480 33.600 8.120 33.880 ;
        RECT 11.760 33.600 13.720 34.720 ;
        RECT 17.640 33.880 21.000 34.720 ;
        RECT 17.640 33.600 21.280 33.880 ;
        RECT 3.920 33.320 8.400 33.600 ;
        RECT 11.480 33.320 14.280 33.600 ;
        RECT 17.080 33.320 21.560 33.600 ;
        RECT 3.920 33.040 8.680 33.320 ;
        RECT 3.920 32.480 5.040 33.040 ;
        RECT 4.200 32.200 4.480 32.480 ;
        RECT 6.720 31.080 8.680 33.040 ;
        RECT 11.200 33.040 14.560 33.320 ;
        RECT 11.200 32.200 12.320 33.040 ;
        RECT 13.160 32.760 14.560 33.040 ;
        RECT 17.080 33.040 21.840 33.320 ;
        RECT 10.640 31.920 12.320 32.200 ;
        RECT 6.720 30.800 8.400 31.080 ;
        RECT 6.440 30.520 8.120 30.800 ;
        RECT 6.160 30.240 7.840 30.520 ;
        RECT 5.880 29.960 7.840 30.240 ;
        RECT 5.600 29.680 7.840 29.960 ;
        RECT 5.320 29.400 7.840 29.680 ;
        RECT 5.320 28.840 7.280 29.400 ;
        RECT 10.360 28.840 12.320 31.920 ;
        RECT 5.320 28.560 7.000 28.840 ;
        RECT 10.640 28.560 12.320 28.840 ;
        RECT 5.040 28.280 6.440 28.560 ;
        RECT 10.920 28.280 12.320 28.560 ;
        RECT 4.480 27.160 6.440 28.280 ;
        RECT 11.200 27.720 12.320 28.280 ;
        RECT 13.440 28.000 15.120 32.760 ;
        RECT 17.080 32.480 18.200 33.040 ;
        RECT 17.360 32.200 17.640 32.480 ;
        RECT 19.880 31.080 21.840 33.040 ;
        RECT 23.520 33.040 28.280 34.720 ;
        RECT 23.520 32.200 25.480 33.040 ;
        RECT 23.520 31.920 25.760 32.200 ;
        RECT 23.520 31.360 27.720 31.920 ;
        RECT 19.880 30.800 21.560 31.080 ;
        RECT 19.600 30.520 21.280 30.800 ;
        RECT 19.320 30.240 21.000 30.520 ;
        RECT 19.040 29.960 21.000 30.240 ;
        RECT 18.760 29.680 21.000 29.960 ;
        RECT 23.520 30.240 28.280 31.360 ;
        RECT 23.520 29.960 25.760 30.240 ;
        RECT 26.040 29.960 28.280 30.240 ;
        RECT 23.520 29.680 25.480 29.960 ;
        RECT 26.320 29.680 28.280 29.960 ;
        RECT 18.480 29.400 21.000 29.680 ;
        RECT 23.800 29.400 25.200 29.680 ;
        RECT 26.600 29.400 28.280 29.680 ;
        RECT 18.480 28.840 20.440 29.400 ;
        RECT 18.480 28.560 20.160 28.840 ;
        RECT 27.160 28.560 28.280 29.400 ;
        RECT 18.200 28.280 19.600 28.560 ;
        RECT 26.880 28.280 28.280 28.560 ;
        RECT 13.160 27.720 14.840 28.000 ;
        RECT 7.560 27.440 8.400 27.720 ;
        RECT 7.560 27.160 8.680 27.440 ;
        RECT 11.200 27.160 14.560 27.720 ;
        RECT 17.640 27.160 19.600 28.280 ;
        RECT 23.520 28.000 24.640 28.280 ;
        RECT 23.520 27.720 24.920 28.000 ;
        RECT 20.720 27.440 21.560 27.720 ;
        RECT 23.520 27.440 25.200 27.720 ;
        RECT 20.720 27.160 21.840 27.440 ;
        RECT 23.800 27.160 25.480 27.440 ;
        RECT 26.600 27.160 28.280 28.280 ;
        RECT 4.200 26.880 6.720 27.160 ;
        RECT 7.280 26.880 8.680 27.160 ;
        RECT 3.920 26.040 8.680 26.880 ;
        RECT 11.760 26.600 14.560 27.160 ;
        RECT 17.360 26.880 19.880 27.160 ;
        RECT 20.440 26.880 21.840 27.160 ;
        RECT 24.080 26.880 25.760 27.160 ;
        RECT 26.320 26.880 27.720 27.160 ;
        RECT 11.760 26.320 14.280 26.600 ;
        RECT 11.760 26.040 13.720 26.320 ;
        RECT 3.920 25.760 8.400 26.040 ;
        RECT 12.040 25.760 13.720 26.040 ;
        RECT 17.080 26.040 21.840 26.880 ;
        RECT 24.360 26.040 27.720 26.880 ;
        RECT 17.080 25.760 21.560 26.040 ;
        RECT 24.360 25.760 27.440 26.040 ;
        RECT 3.080 22.960 8.680 24.640 ;
        RECT 11.760 24.080 18.200 24.640 ;
        RECT 3.360 22.680 8.680 22.960 ;
        RECT 11.200 22.960 18.200 24.080 ;
        RECT 11.200 22.680 14.280 22.960 ;
        RECT 15.680 22.680 18.200 22.960 ;
        RECT 3.640 22.400 8.680 22.680 ;
        RECT 10.640 22.400 13.720 22.680 ;
        RECT 3.920 22.120 8.680 22.400 ;
        RECT 10.360 22.120 13.720 22.400 ;
        RECT 16.240 22.400 18.480 22.680 ;
        RECT 4.200 21.840 7.280 22.120 ;
        RECT 0.840 14.280 3.360 15.120 ;
        RECT 0.840 13.720 3.640 14.280 ;
        RECT 4.480 13.720 7.280 21.840 ;
        RECT 10.360 21.560 13.160 22.120 ;
        RECT 10.360 20.160 12.880 21.560 ;
        RECT 16.240 20.720 18.760 22.400 ;
        RECT 10.360 19.600 13.160 20.160 ;
        RECT 10.360 19.320 13.720 19.600 ;
        RECT 10.640 19.040 13.720 19.320 ;
        RECT 16.240 19.040 17.360 19.600 ;
        RECT 19.880 19.320 22.400 24.640 ;
        RECT 25.760 23.520 28.280 24.640 ;
        RECT 25.480 23.240 28.280 23.520 ;
        RECT 25.200 22.960 28.280 23.240 ;
        RECT 24.920 22.680 28.000 22.960 ;
        RECT 24.920 21.280 27.720 22.680 ;
        RECT 24.640 21.000 27.720 21.280 ;
        RECT 23.520 20.720 27.720 21.000 ;
        RECT 23.520 20.440 26.600 20.720 ;
        RECT 23.520 20.160 26.320 20.440 ;
        RECT 19.880 19.040 22.680 19.320 ;
        RECT 23.520 19.040 26.040 20.160 ;
        RECT 10.920 18.760 14.000 19.040 ;
        RECT 15.960 18.760 17.640 19.040 ;
        RECT 19.880 18.760 22.960 19.040 ;
        RECT 23.240 18.760 26.040 19.040 ;
        RECT 11.200 17.640 18.200 18.760 ;
        RECT 19.880 18.480 26.040 18.760 ;
        RECT 19.880 18.200 24.920 18.480 ;
        RECT 19.880 17.640 24.640 18.200 ;
        RECT 11.760 17.360 18.480 17.640 ;
        RECT 19.880 17.360 24.920 17.640 ;
        RECT 11.760 17.080 18.760 17.360 ;
        RECT 15.960 16.800 18.760 17.080 ;
        RECT 10.360 14.280 12.880 15.120 ;
        RECT 10.360 13.720 13.160 14.280 ;
        RECT 16.240 14.000 18.760 16.800 ;
        RECT 15.960 13.720 18.760 14.000 ;
        RECT 0.840 13.440 7.000 13.720 ;
        RECT 10.360 13.440 18.760 13.720 ;
        RECT 19.880 17.080 26.040 17.360 ;
        RECT 19.880 16.800 22.960 17.080 ;
        RECT 23.240 16.800 26.040 17.080 ;
        RECT 19.880 16.520 22.680 16.800 ;
        RECT 1.120 13.160 6.720 13.440 ;
        RECT 10.640 13.160 18.480 13.440 ;
        RECT 1.680 12.040 6.440 13.160 ;
        RECT 1.960 11.760 6.440 12.040 ;
        RECT 11.200 11.760 18.200 13.160 ;
        RECT 2.240 11.480 6.440 11.760 ;
        RECT 2.520 11.200 6.440 11.480 ;
        RECT 11.760 11.200 18.200 11.760 ;
        RECT 19.880 11.200 22.400 16.520 ;
        RECT 23.520 15.680 26.040 16.800 ;
        RECT 23.520 15.400 26.320 15.680 ;
        RECT 23.520 15.120 26.600 15.400 ;
        RECT 23.520 14.840 27.720 15.120 ;
        RECT 24.640 14.560 27.720 14.840 ;
        RECT 24.920 14.000 27.720 14.560 ;
        RECT 24.920 13.720 28.000 14.000 ;
        RECT 24.920 13.440 28.280 13.720 ;
        RECT 25.480 13.160 28.280 13.440 ;
        RECT 25.760 11.200 28.280 13.160 ;
        RECT 3.080 9.520 7.840 10.080 ;
        RECT 9.800 9.800 14.280 10.080 ;
        RECT 9.800 9.520 14.560 9.800 ;
        RECT 18.480 9.520 19.600 10.080 ;
        RECT 3.080 8.960 8.400 9.520 ;
        RECT 9.800 9.240 14.840 9.520 ;
        RECT 17.920 9.240 19.600 9.520 ;
        RECT 9.800 8.960 15.120 9.240 ;
        RECT 3.080 8.680 8.120 8.960 ;
        RECT 9.800 8.680 14.840 8.960 ;
        RECT 17.640 8.680 19.600 9.240 ;
        RECT 24.360 8.960 26.040 10.080 ;
        RECT 24.080 8.680 26.320 8.960 ;
        RECT 3.080 8.400 7.840 8.680 ;
        RECT 9.800 8.400 14.560 8.680 ;
        RECT 3.360 8.120 7.560 8.400 ;
        RECT 9.800 8.120 14.280 8.400 ;
        RECT 4.480 1.120 6.440 8.120 ;
        RECT 10.920 7.840 13.160 8.120 ;
        RECT 4.760 0.840 6.160 1.120 ;
        RECT 11.200 0.840 12.880 7.840 ;
        RECT 17.080 7.560 19.600 8.680 ;
        RECT 23.800 8.400 26.880 8.680 ;
        RECT 17.360 7.280 19.600 7.560 ;
        RECT 23.520 8.120 26.880 8.400 ;
        RECT 23.520 7.840 24.920 8.120 ;
        RECT 25.760 7.840 27.160 8.120 ;
        RECT 23.520 7.280 24.640 7.840 ;
        RECT 17.640 3.080 19.600 7.280 ;
        RECT 22.960 3.920 24.640 7.280 ;
        RECT 23.240 3.640 24.640 3.920 ;
        RECT 23.520 3.080 24.640 3.640 ;
        RECT 25.760 7.560 27.440 7.840 ;
        RECT 25.760 3.360 27.720 7.560 ;
        RECT 25.760 3.080 27.440 3.360 ;
        RECT 17.640 2.800 19.880 3.080 ;
        RECT 23.520 2.800 24.920 3.080 ;
        RECT 25.760 2.800 27.160 3.080 ;
        RECT 17.080 2.520 20.160 2.800 ;
        RECT 23.520 2.520 26.880 2.800 ;
        RECT 17.080 2.240 20.440 2.520 ;
        RECT 23.800 2.240 26.880 2.520 ;
        RECT 17.080 1.960 20.720 2.240 ;
        RECT 24.080 1.960 26.880 2.240 ;
        RECT 17.080 0.840 21.000 1.960 ;
        RECT 24.360 1.680 26.880 1.960 ;
        RECT 24.360 1.400 26.600 1.680 ;
        RECT 24.360 1.120 26.320 1.400 ;
        RECT 24.360 0.840 26.040 1.120 ;
      LAYER met4 ;
        RECT 4.760 34.720 7.840 35.000 ;
        RECT 12.040 34.720 13.720 35.000 ;
        RECT 17.920 34.720 21.000 35.000 ;
        RECT 23.800 34.720 28.280 35.000 ;
        RECT 4.480 33.880 7.840 34.720 ;
        RECT 4.480 33.600 8.120 33.880 ;
        RECT 11.760 33.600 13.720 34.720 ;
        RECT 17.640 33.880 21.000 34.720 ;
        RECT 17.640 33.600 21.280 33.880 ;
        RECT 3.920 33.320 8.400 33.600 ;
        RECT 11.480 33.320 14.280 33.600 ;
        RECT 17.080 33.320 21.560 33.600 ;
        RECT 3.920 33.040 8.680 33.320 ;
        RECT 3.920 32.480 5.040 33.040 ;
        RECT 4.200 32.200 4.480 32.480 ;
        RECT 6.720 31.080 8.680 33.040 ;
        RECT 11.200 33.040 14.560 33.320 ;
        RECT 11.200 32.200 12.320 33.040 ;
        RECT 13.160 32.760 14.560 33.040 ;
        RECT 17.080 33.040 21.840 33.320 ;
        RECT 10.640 31.920 12.320 32.200 ;
        RECT 6.720 30.800 8.400 31.080 ;
        RECT 6.440 30.520 8.120 30.800 ;
        RECT 6.160 30.240 7.840 30.520 ;
        RECT 5.880 29.960 7.840 30.240 ;
        RECT 5.600 29.680 7.840 29.960 ;
        RECT 5.320 29.400 7.840 29.680 ;
        RECT 5.320 28.840 7.280 29.400 ;
        RECT 10.360 28.840 12.320 31.920 ;
        RECT 5.320 28.560 7.000 28.840 ;
        RECT 10.640 28.560 12.320 28.840 ;
        RECT 5.040 28.280 6.440 28.560 ;
        RECT 10.920 28.280 12.320 28.560 ;
        RECT 4.480 27.160 6.440 28.280 ;
        RECT 11.200 27.720 12.320 28.280 ;
        RECT 13.440 28.000 15.120 32.760 ;
        RECT 17.080 32.480 18.200 33.040 ;
        RECT 17.360 32.200 17.640 32.480 ;
        RECT 19.880 31.080 21.840 33.040 ;
        RECT 23.520 33.040 28.280 34.720 ;
        RECT 23.520 32.200 25.480 33.040 ;
        RECT 23.520 31.920 25.760 32.200 ;
        RECT 23.520 31.360 27.720 31.920 ;
        RECT 19.880 30.800 21.560 31.080 ;
        RECT 19.600 30.520 21.280 30.800 ;
        RECT 19.320 30.240 21.000 30.520 ;
        RECT 19.040 29.960 21.000 30.240 ;
        RECT 18.760 29.680 21.000 29.960 ;
        RECT 23.520 30.240 28.280 31.360 ;
        RECT 23.520 29.960 25.760 30.240 ;
        RECT 26.040 29.960 28.280 30.240 ;
        RECT 23.520 29.680 25.480 29.960 ;
        RECT 26.320 29.680 28.280 29.960 ;
        RECT 18.480 29.400 21.000 29.680 ;
        RECT 23.800 29.400 25.200 29.680 ;
        RECT 26.600 29.400 28.280 29.680 ;
        RECT 18.480 28.840 20.440 29.400 ;
        RECT 18.480 28.560 20.160 28.840 ;
        RECT 27.160 28.560 28.280 29.400 ;
        RECT 18.200 28.280 19.600 28.560 ;
        RECT 26.880 28.280 28.280 28.560 ;
        RECT 13.160 27.720 14.840 28.000 ;
        RECT 7.560 27.440 8.400 27.720 ;
        RECT 7.560 27.160 8.680 27.440 ;
        RECT 11.200 27.160 14.560 27.720 ;
        RECT 17.640 27.160 19.600 28.280 ;
        RECT 23.520 28.000 24.640 28.280 ;
        RECT 23.520 27.720 24.920 28.000 ;
        RECT 20.720 27.440 21.560 27.720 ;
        RECT 23.520 27.440 25.200 27.720 ;
        RECT 20.720 27.160 21.840 27.440 ;
        RECT 23.800 27.160 25.480 27.440 ;
        RECT 26.600 27.160 28.280 28.280 ;
        RECT 4.200 26.880 6.720 27.160 ;
        RECT 7.280 26.880 8.680 27.160 ;
        RECT 3.920 26.040 8.680 26.880 ;
        RECT 11.760 26.600 14.560 27.160 ;
        RECT 17.360 26.880 19.880 27.160 ;
        RECT 20.440 26.880 21.840 27.160 ;
        RECT 24.080 26.880 25.760 27.160 ;
        RECT 26.320 26.880 27.720 27.160 ;
        RECT 11.760 26.320 14.280 26.600 ;
        RECT 11.760 26.040 13.720 26.320 ;
        RECT 3.920 25.760 8.400 26.040 ;
        RECT 12.040 25.760 13.720 26.040 ;
        RECT 17.080 26.040 21.840 26.880 ;
        RECT 24.360 26.040 27.720 26.880 ;
        RECT 17.080 25.760 21.560 26.040 ;
        RECT 24.360 25.760 27.440 26.040 ;
        RECT 3.080 22.960 8.680 24.640 ;
        RECT 11.760 24.080 18.200 24.640 ;
        RECT 3.360 22.680 8.680 22.960 ;
        RECT 11.200 22.960 18.200 24.080 ;
        RECT 11.200 22.680 14.280 22.960 ;
        RECT 15.680 22.680 18.200 22.960 ;
        RECT 3.640 22.400 8.680 22.680 ;
        RECT 10.640 22.400 13.720 22.680 ;
        RECT 3.920 22.120 8.680 22.400 ;
        RECT 10.360 22.120 13.720 22.400 ;
        RECT 16.240 22.400 18.480 22.680 ;
        RECT 4.200 21.840 7.280 22.120 ;
        RECT 0.840 14.280 3.360 15.120 ;
        RECT 0.840 13.720 3.640 14.280 ;
        RECT 4.480 13.720 7.280 21.840 ;
        RECT 10.360 21.560 13.160 22.120 ;
        RECT 10.360 20.160 12.880 21.560 ;
        RECT 16.240 20.720 18.760 22.400 ;
        RECT 10.360 19.600 13.160 20.160 ;
        RECT 10.360 19.320 13.720 19.600 ;
        RECT 10.640 19.040 13.720 19.320 ;
        RECT 16.240 19.040 17.360 19.600 ;
        RECT 19.880 19.320 22.400 24.640 ;
        RECT 25.760 23.520 28.280 24.640 ;
        RECT 25.480 23.240 28.280 23.520 ;
        RECT 25.200 22.960 28.280 23.240 ;
        RECT 24.920 22.680 28.000 22.960 ;
        RECT 24.920 21.280 27.720 22.680 ;
        RECT 24.640 21.000 27.720 21.280 ;
        RECT 23.520 20.720 27.720 21.000 ;
        RECT 23.520 20.440 26.600 20.720 ;
        RECT 23.520 20.160 26.320 20.440 ;
        RECT 19.880 19.040 22.680 19.320 ;
        RECT 23.520 19.040 26.040 20.160 ;
        RECT 10.920 18.760 14.000 19.040 ;
        RECT 15.960 18.760 17.640 19.040 ;
        RECT 19.880 18.760 22.960 19.040 ;
        RECT 23.240 18.760 26.040 19.040 ;
        RECT 11.200 17.640 18.200 18.760 ;
        RECT 19.880 18.480 26.040 18.760 ;
        RECT 19.880 18.200 24.920 18.480 ;
        RECT 19.880 17.640 24.640 18.200 ;
        RECT 11.760 17.360 18.480 17.640 ;
        RECT 19.880 17.360 24.920 17.640 ;
        RECT 11.760 17.080 18.760 17.360 ;
        RECT 15.960 16.800 18.760 17.080 ;
        RECT 10.360 14.280 12.880 15.120 ;
        RECT 10.360 13.720 13.160 14.280 ;
        RECT 16.240 14.000 18.760 16.800 ;
        RECT 15.960 13.720 18.760 14.000 ;
        RECT 0.840 13.440 7.000 13.720 ;
        RECT 10.360 13.440 18.760 13.720 ;
        RECT 19.880 17.080 26.040 17.360 ;
        RECT 19.880 16.800 22.960 17.080 ;
        RECT 23.240 16.800 26.040 17.080 ;
        RECT 19.880 16.520 22.680 16.800 ;
        RECT 1.120 13.160 6.720 13.440 ;
        RECT 10.640 13.160 18.480 13.440 ;
        RECT 1.680 12.040 6.440 13.160 ;
        RECT 1.960 11.760 6.440 12.040 ;
        RECT 11.200 11.760 18.200 13.160 ;
        RECT 2.240 11.480 6.440 11.760 ;
        RECT 2.520 11.200 6.440 11.480 ;
        RECT 11.760 11.200 18.200 11.760 ;
        RECT 19.880 11.200 22.400 16.520 ;
        RECT 23.520 15.680 26.040 16.800 ;
        RECT 23.520 15.400 26.320 15.680 ;
        RECT 23.520 15.120 26.600 15.400 ;
        RECT 23.520 14.840 27.720 15.120 ;
        RECT 24.640 14.560 27.720 14.840 ;
        RECT 24.920 14.000 27.720 14.560 ;
        RECT 24.920 13.720 28.000 14.000 ;
        RECT 24.920 13.440 28.280 13.720 ;
        RECT 25.480 13.160 28.280 13.440 ;
        RECT 25.760 11.200 28.280 13.160 ;
        RECT 3.080 9.520 7.840 10.080 ;
        RECT 9.800 9.800 14.280 10.080 ;
        RECT 9.800 9.520 14.560 9.800 ;
        RECT 18.480 9.520 19.600 10.080 ;
        RECT 3.080 8.960 8.400 9.520 ;
        RECT 9.800 9.240 14.840 9.520 ;
        RECT 17.920 9.240 19.600 9.520 ;
        RECT 9.800 8.960 15.120 9.240 ;
        RECT 3.080 8.680 8.120 8.960 ;
        RECT 9.800 8.680 14.840 8.960 ;
        RECT 17.640 8.680 19.600 9.240 ;
        RECT 24.360 8.960 26.040 10.080 ;
        RECT 24.080 8.680 26.320 8.960 ;
        RECT 3.080 8.400 7.840 8.680 ;
        RECT 9.800 8.400 14.560 8.680 ;
        RECT 3.360 8.120 7.560 8.400 ;
        RECT 9.800 8.120 14.280 8.400 ;
        RECT 4.480 1.120 6.440 8.120 ;
        RECT 10.920 7.840 13.160 8.120 ;
        RECT 4.760 0.840 6.160 1.120 ;
        RECT 11.200 0.840 12.880 7.840 ;
        RECT 17.080 7.560 19.600 8.680 ;
        RECT 23.800 8.400 26.880 8.680 ;
        RECT 17.360 7.280 19.600 7.560 ;
        RECT 23.520 8.120 26.880 8.400 ;
        RECT 23.520 7.840 24.920 8.120 ;
        RECT 25.760 7.840 27.160 8.120 ;
        RECT 23.520 7.280 24.640 7.840 ;
        RECT 17.640 3.080 19.600 7.280 ;
        RECT 22.960 3.920 24.640 7.280 ;
        RECT 23.240 3.640 24.640 3.920 ;
        RECT 23.520 3.080 24.640 3.640 ;
        RECT 25.760 7.560 27.440 7.840 ;
        RECT 25.760 3.360 27.720 7.560 ;
        RECT 25.760 3.080 27.440 3.360 ;
        RECT 17.640 2.800 19.880 3.080 ;
        RECT 23.520 2.800 24.920 3.080 ;
        RECT 25.760 2.800 27.160 3.080 ;
        RECT 17.080 2.520 20.160 2.800 ;
        RECT 23.520 2.520 26.880 2.800 ;
        RECT 17.080 2.240 20.440 2.520 ;
        RECT 23.800 2.240 26.880 2.520 ;
        RECT 17.080 1.960 20.720 2.240 ;
        RECT 24.080 1.960 26.880 2.240 ;
        RECT 17.080 0.840 21.000 1.960 ;
        RECT 24.360 1.680 26.880 1.960 ;
        RECT 24.360 1.400 26.600 1.680 ;
        RECT 24.360 1.120 26.320 1.400 ;
        RECT 24.360 0.840 26.040 1.120 ;
  END
END my_logo
END LIBRARY

