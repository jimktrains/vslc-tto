module tt_um_jimktrains_vslc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire clknet_0_clk;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire \cur_addr[0] ;
 wire \cur_addr[1] ;
 wire \cur_addr[2] ;
 wire \cur_addr[3] ;
 wire \cur_addr[4] ;
 wire \cur_addr[5] ;
 wire \cur_addr[6] ;
 wire \cur_addr[7] ;
 wire \cycle_end_addr[0] ;
 wire \cycle_end_addr[1] ;
 wire \cycle_end_addr[2] ;
 wire \cycle_end_addr[3] ;
 wire \cycle_end_addr[4] ;
 wire \cycle_end_addr[5] ;
 wire \cycle_end_addr[6] ;
 wire \cycle_end_addr[7] ;
 wire \cycle_start_addr[0] ;
 wire \cycle_start_addr[1] ;
 wire \cycle_start_addr[2] ;
 wire \cycle_start_addr[3] ;
 wire \cycle_start_addr[4] ;
 wire \cycle_start_addr[5] ;
 wire \cycle_start_addr[6] ;
 wire \cycle_start_addr[7] ;
 wire eeprom_copi;
 wire eeprom_cs;
 wire eeprom_oe_copi;
 wire eeprom_sck;
 wire \fetch_count[0] ;
 wire \fetch_count[1] ;
 wire \fetch_count[2] ;
 wire \fetch_prev_state[0] ;
 wire \fetch_prev_state[1] ;
 wire \fetch_prev_state[2] ;
 wire \fetch_prev_state[3] ;
 wire \fetch_state[0] ;
 wire \fetch_state[1] ;
 wire \fetch_state[2] ;
 wire \fetch_state[3] ;
 wire \instr[0] ;
 wire \instr[1] ;
 wire \instr[2] ;
 wire \instr[3] ;
 wire \instr[4] ;
 wire \instr[5] ;
 wire \instr[6] ;
 wire \instr[7] ;
 wire \stack[0] ;
 wire \stack[10] ;
 wire \stack[11] ;
 wire \stack[12] ;
 wire \stack[13] ;
 wire \stack[14] ;
 wire \stack[15] ;
 wire \stack[1] ;
 wire \stack[2] ;
 wire \stack[3] ;
 wire \stack[4] ;
 wire \stack[5] ;
 wire \stack[6] ;
 wire \stack[7] ;
 wire \stack[8] ;
 wire \stack[9] ;
 wire stack_out;
 wire \timer_clock_counter[0] ;
 wire \timer_clock_counter[10] ;
 wire \timer_clock_counter[11] ;
 wire \timer_clock_counter[12] ;
 wire \timer_clock_counter[13] ;
 wire \timer_clock_counter[14] ;
 wire \timer_clock_counter[15] ;
 wire \timer_clock_counter[1] ;
 wire \timer_clock_counter[2] ;
 wire \timer_clock_counter[3] ;
 wire \timer_clock_counter[4] ;
 wire \timer_clock_counter[5] ;
 wire \timer_clock_counter[6] ;
 wire \timer_clock_counter[7] ;
 wire \timer_clock_counter[8] ;
 wire \timer_clock_counter[9] ;
 wire \timer_clock_divisor[0] ;
 wire \timer_clock_divisor[1] ;
 wire \timer_clock_divisor[2] ;
 wire \timer_clock_divisor[3] ;
 wire \timer_counter[0] ;
 wire \timer_counter[10] ;
 wire \timer_counter[11] ;
 wire \timer_counter[12] ;
 wire \timer_counter[13] ;
 wire \timer_counter[14] ;
 wire \timer_counter[15] ;
 wire \timer_counter[1] ;
 wire \timer_counter[2] ;
 wire \timer_counter[3] ;
 wire \timer_counter[4] ;
 wire \timer_counter[5] ;
 wire \timer_counter[6] ;
 wire \timer_counter[7] ;
 wire \timer_counter[8] ;
 wire \timer_counter[9] ;
 wire timer_enabled;
 wire timer_mode;
 wire timer_out;
 wire \timer_period_a[0] ;
 wire \timer_period_a[10] ;
 wire \timer_period_a[11] ;
 wire \timer_period_a[12] ;
 wire \timer_period_a[13] ;
 wire \timer_period_a[14] ;
 wire \timer_period_a[15] ;
 wire \timer_period_a[1] ;
 wire \timer_period_a[2] ;
 wire \timer_period_a[3] ;
 wire \timer_period_a[4] ;
 wire \timer_period_a[5] ;
 wire \timer_period_a[6] ;
 wire \timer_period_a[7] ;
 wire \timer_period_a[8] ;
 wire \timer_period_a[9] ;
 wire \timer_period_b[0] ;
 wire \timer_period_b[10] ;
 wire \timer_period_b[11] ;
 wire \timer_period_b[12] ;
 wire \timer_period_b[13] ;
 wire \timer_period_b[14] ;
 wire \timer_period_b[15] ;
 wire \timer_period_b[1] ;
 wire \timer_period_b[2] ;
 wire \timer_period_b[3] ;
 wire \timer_period_b[4] ;
 wire \timer_period_b[5] ;
 wire \timer_period_b[6] ;
 wire \timer_period_b[7] ;
 wire \timer_period_b[8] ;
 wire \timer_period_b[9] ;
 wire timer_phase;
 wire \ui_in_reg[0] ;
 wire \ui_in_reg[1] ;
 wire \ui_in_reg[2] ;
 wire \ui_in_reg[3] ;
 wire \ui_in_reg[4] ;
 wire \ui_in_reg[5] ;
 wire \ui_in_reg[6] ;
 wire \ui_in_reg[7] ;
 wire \uio_in_reg[3] ;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net71;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;

 sky130_fd_sc_hd__inv_2 _0754_ (.A(net54),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(timer_phase),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(\timer_counter[13] ),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(\timer_counter[10] ),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(\timer_counter[9] ),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(\timer_counter[8] ),
    .Y(_0330_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(\timer_counter[7] ),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(\timer_counter[6] ),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(\timer_counter[2] ),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(net44),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(net46),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(net49),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(\cur_addr[7] ),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(net240),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(\cur_addr[5] ),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(net247),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(\cur_addr[3] ),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(\cur_addr[2] ),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(\fetch_count[2] ),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(\timer_period_a[0] ),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(\timer_period_a[6] ),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(\timer_period_a[11] ),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(\timer_period_a[14] ),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(\timer_period_b[0] ),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(\timer_period_b[1] ),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(\timer_period_b[4] ),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(\timer_period_b[8] ),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _1367__3 (.A(clknet_4_7_0_clk),
    .Y(net72));
 sky130_fd_sc_hd__nand3_1 _0782_ (.A(\fetch_count[2] ),
    .B(\fetch_count[1] ),
    .C(\fetch_count[0] ),
    .Y(_0352_));
 sky130_fd_sc_hd__or3b_4 _0783_ (.A(\fetch_prev_state[2] ),
    .B(_0352_),
    .C_N(\fetch_prev_state[3] ),
    .X(_0353_));
 sky130_fd_sc_hd__nor3_4 _0784_ (.A(\fetch_prev_state[1] ),
    .B(\fetch_prev_state[0] ),
    .C(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__mux4_1 _0785_ (.A0(\timer_clock_counter[12] ),
    .A1(\timer_clock_counter[13] ),
    .A2(\timer_clock_counter[14] ),
    .A3(\timer_clock_counter[15] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0355_));
 sky130_fd_sc_hd__mux4_1 _0786_ (.A0(\timer_clock_counter[8] ),
    .A1(\timer_clock_counter[9] ),
    .A2(\timer_clock_counter[10] ),
    .A3(\timer_clock_counter[11] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0356_));
 sky130_fd_sc_hd__nand2b_1 _0787_ (.A_N(\timer_clock_divisor[2] ),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__a21boi_1 _0788_ (.A1(\timer_clock_divisor[2] ),
    .A2(_0355_),
    .B1_N(\timer_clock_divisor[3] ),
    .Y(_0358_));
 sky130_fd_sc_hd__mux4_1 _0789_ (.A0(\timer_clock_counter[0] ),
    .A1(\timer_clock_counter[1] ),
    .A2(\timer_clock_counter[2] ),
    .A3(\timer_clock_counter[3] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0359_));
 sky130_fd_sc_hd__mux4_1 _0790_ (.A0(\timer_clock_counter[4] ),
    .A1(\timer_clock_counter[5] ),
    .A2(\timer_clock_counter[6] ),
    .A3(\timer_clock_counter[7] ),
    .S0(\timer_clock_divisor[0] ),
    .S1(\timer_clock_divisor[1] ),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(_0359_),
    .A1(_0360_),
    .S(\timer_clock_divisor[2] ),
    .X(_0361_));
 sky130_fd_sc_hd__o2bb2a_2 _0792_ (.A1_N(_0357_),
    .A2_N(_0358_),
    .B1(_0361_),
    .B2(\timer_clock_divisor[3] ),
    .X(_0362_));
 sky130_fd_sc_hd__and2b_1 _0793_ (.A_N(\timer_counter[3] ),
    .B(\timer_period_b[3] ),
    .X(_0363_));
 sky130_fd_sc_hd__and2b_1 _0794_ (.A_N(\timer_counter[5] ),
    .B(\timer_period_b[5] ),
    .X(_0364_));
 sky130_fd_sc_hd__and2b_1 _0795_ (.A_N(\timer_period_b[12] ),
    .B(\timer_counter[12] ),
    .X(_0365_));
 sky130_fd_sc_hd__and2b_1 _0796_ (.A_N(\timer_period_b[9] ),
    .B(\timer_counter[9] ),
    .X(_0366_));
 sky130_fd_sc_hd__and2b_1 _0797_ (.A_N(\timer_counter[1] ),
    .B(\timer_period_b[1] ),
    .X(_0367_));
 sky130_fd_sc_hd__and2b_1 _0798_ (.A_N(\timer_counter[2] ),
    .B(\timer_period_b[2] ),
    .X(_0368_));
 sky130_fd_sc_hd__xor2_1 _0799_ (.A(\timer_counter[15] ),
    .B(\timer_period_b[15] ),
    .X(_0369_));
 sky130_fd_sc_hd__xor2_1 _0800_ (.A(\timer_counter[11] ),
    .B(\timer_period_b[11] ),
    .X(_0370_));
 sky130_fd_sc_hd__and2b_1 _0801_ (.A_N(\timer_period_b[5] ),
    .B(\timer_counter[5] ),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_1 _0802_ (.A(_0332_),
    .B(\timer_period_b[6] ),
    .Y(_0372_));
 sky130_fd_sc_hd__and2b_1 _0803_ (.A_N(\timer_period_b[3] ),
    .B(\timer_counter[3] ),
    .X(_0373_));
 sky130_fd_sc_hd__and2b_1 _0804_ (.A_N(\timer_counter[12] ),
    .B(\timer_period_b[12] ),
    .X(_0374_));
 sky130_fd_sc_hd__and2b_1 _0805_ (.A_N(\timer_counter[10] ),
    .B(\timer_period_b[10] ),
    .X(_0375_));
 sky130_fd_sc_hd__and2b_1 _0806_ (.A_N(\timer_counter[7] ),
    .B(\timer_period_b[7] ),
    .X(_0376_));
 sky130_fd_sc_hd__nor2_1 _0807_ (.A(\timer_counter[4] ),
    .B(_0350_),
    .Y(_0377_));
 sky130_fd_sc_hd__and2b_1 _0808_ (.A_N(\timer_period_b[1] ),
    .B(\timer_counter[1] ),
    .X(_0378_));
 sky130_fd_sc_hd__and2b_1 _0809_ (.A_N(\timer_period_b[2] ),
    .B(\timer_counter[2] ),
    .X(_0379_));
 sky130_fd_sc_hd__and2b_1 _0810_ (.A_N(\timer_counter[8] ),
    .B(\timer_period_b[8] ),
    .X(_0380_));
 sky130_fd_sc_hd__a22o_1 _0811_ (.A1(_0332_),
    .A2(\timer_period_b[6] ),
    .B1(\timer_period_b[9] ),
    .B2(_0329_),
    .X(_0381_));
 sky130_fd_sc_hd__a2111o_1 _0812_ (.A1(\timer_counter[0] ),
    .A2(_0348_),
    .B1(_0369_),
    .C1(_0381_),
    .D1(_0326_),
    .X(_0382_));
 sky130_fd_sc_hd__or3_1 _0813_ (.A(_0364_),
    .B(_0366_),
    .C(_0379_),
    .X(_0383_));
 sky130_fd_sc_hd__xor2_1 _0814_ (.A(\timer_counter[14] ),
    .B(\timer_period_b[14] ),
    .X(_0384_));
 sky130_fd_sc_hd__a221o_1 _0815_ (.A1(\timer_counter[8] ),
    .A2(_0351_),
    .B1(\timer_period_b[13] ),
    .B2(_0327_),
    .C1(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__o22ai_1 _0816_ (.A1(\timer_counter[0] ),
    .A2(_0348_),
    .B1(\timer_period_b[7] ),
    .B2(_0331_),
    .Y(_0386_));
 sky130_fd_sc_hd__nor2_1 _0817_ (.A(_0327_),
    .B(\timer_period_b[13] ),
    .Y(_0387_));
 sky130_fd_sc_hd__or4_1 _0818_ (.A(_0383_),
    .B(_0385_),
    .C(_0386_),
    .D(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__or4_1 _0819_ (.A(_0370_),
    .B(_0376_),
    .C(_0378_),
    .D(_0380_),
    .X(_0389_));
 sky130_fd_sc_hd__or3_1 _0820_ (.A(_0363_),
    .B(_0367_),
    .C(_0373_),
    .X(_0390_));
 sky130_fd_sc_hd__a2bb2o_1 _0821_ (.A1_N(_0328_),
    .A2_N(\timer_period_b[10] ),
    .B1(\timer_counter[4] ),
    .B2(_0350_),
    .X(_0391_));
 sky130_fd_sc_hd__or4_1 _0822_ (.A(_0365_),
    .B(_0389_),
    .C(_0390_),
    .D(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__or3_1 _0823_ (.A(_0368_),
    .B(_0371_),
    .C(_0375_),
    .X(_0393_));
 sky130_fd_sc_hd__or4_1 _0824_ (.A(_0372_),
    .B(_0374_),
    .C(_0377_),
    .D(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__nor4_1 _0825_ (.A(_0382_),
    .B(_0388_),
    .C(_0392_),
    .D(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__and2_1 _0826_ (.A(timer_mode),
    .B(net18),
    .X(_0396_));
 sky130_fd_sc_hd__and3_2 _0827_ (.A(timer_mode),
    .B(_0362_),
    .C(net18),
    .X(_0397_));
 sky130_fd_sc_hd__a2111o_1 _0828_ (.A1(\timer_counter[0] ),
    .A2(_0348_),
    .B1(_0371_),
    .C1(_0375_),
    .D1(_0377_),
    .X(_0398_));
 sky130_fd_sc_hd__or4_1 _0829_ (.A(_0364_),
    .B(_0366_),
    .C(_0368_),
    .D(_0379_),
    .X(_0399_));
 sky130_fd_sc_hd__or4_1 _0830_ (.A(_0372_),
    .B(_0381_),
    .C(_0398_),
    .D(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _0831_ (.A(_0326_),
    .B(_0365_),
    .C(_0376_),
    .D(_0380_),
    .X(_0401_));
 sky130_fd_sc_hd__or4_1 _0832_ (.A(_0374_),
    .B(_0387_),
    .C(_0391_),
    .D(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__or4_1 _0833_ (.A(_0369_),
    .B(_0385_),
    .C(_0386_),
    .D(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__or4_1 _0834_ (.A(_0363_),
    .B(_0367_),
    .C(_0373_),
    .D(_0378_),
    .X(_0404_));
 sky130_fd_sc_hd__or4_1 _0835_ (.A(_0370_),
    .B(_0400_),
    .C(_0403_),
    .D(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__nor2_2 _0836_ (.A(_0354_),
    .B(_0397_),
    .Y(_0406_));
 sky130_fd_sc_hd__a32o_1 _0837_ (.A1(net30),
    .A2(\timer_period_b[15] ),
    .A3(_0406_),
    .B1(_0354_),
    .B2(net34),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _0838_ (.A(net51),
    .B(_0407_),
    .X(_0285_));
 sky130_fd_sc_hd__a32o_1 _0839_ (.A1(net30),
    .A2(\timer_period_b[14] ),
    .A3(_0406_),
    .B1(_0354_),
    .B2(net35),
    .X(_0408_));
 sky130_fd_sc_hd__and2_1 _0840_ (.A(net52),
    .B(_0408_),
    .X(_0284_));
 sky130_fd_sc_hd__a32o_1 _0841_ (.A1(net30),
    .A2(\timer_period_b[13] ),
    .A3(_0406_),
    .B1(_0354_),
    .B2(net38),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _0842_ (.A(net58),
    .B(_0409_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_1 _0843_ (.A(net52),
    .B(net39),
    .X(_0410_));
 sky130_fd_sc_hd__nand2_1 _0844_ (.A(net52),
    .B(net39),
    .Y(_0411_));
 sky130_fd_sc_hd__and2_1 _0845_ (.A(net52),
    .B(net30),
    .X(_0412_));
 sky130_fd_sc_hd__nand2_1 _0846_ (.A(net51),
    .B(net30),
    .Y(_0413_));
 sky130_fd_sc_hd__a32o_1 _0847_ (.A1(net233),
    .A2(_0406_),
    .A3(_0412_),
    .B1(_0410_),
    .B2(_0354_),
    .X(_0282_));
 sky130_fd_sc_hd__a32o_1 _0848_ (.A1(net31),
    .A2(\timer_period_b[11] ),
    .A3(_0406_),
    .B1(_0354_),
    .B2(net42),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _0849_ (.A(net58),
    .B(_0414_),
    .X(_0281_));
 sky130_fd_sc_hd__a32o_1 _0850_ (.A1(net31),
    .A2(\timer_period_b[10] ),
    .A3(_0406_),
    .B1(_0354_),
    .B2(net44),
    .X(_0415_));
 sky130_fd_sc_hd__and2_1 _0851_ (.A(net58),
    .B(_0415_),
    .X(_0280_));
 sky130_fd_sc_hd__a32o_1 _0852_ (.A1(net30),
    .A2(\timer_period_b[9] ),
    .A3(_0406_),
    .B1(_0354_),
    .B2(net45),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(net51),
    .B(_0416_),
    .X(_0279_));
 sky130_fd_sc_hd__a32o_1 _0854_ (.A1(net30),
    .A2(\timer_period_b[8] ),
    .A3(_0406_),
    .B1(_0354_),
    .B2(net48),
    .X(_0417_));
 sky130_fd_sc_hd__and2_1 _0855_ (.A(net51),
    .B(_0417_),
    .X(_0278_));
 sky130_fd_sc_hd__nor3b_1 _0856_ (.A(_0353_),
    .B(\fetch_prev_state[1] ),
    .C_N(\fetch_prev_state[0] ),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_2 _0857_ (.A(_0397_),
    .B(net19),
    .Y(_0419_));
 sky130_fd_sc_hd__a32o_1 _0858_ (.A1(net31),
    .A2(\timer_period_b[7] ),
    .A3(_0419_),
    .B1(net19),
    .B2(net34),
    .X(_0420_));
 sky130_fd_sc_hd__and2_1 _0859_ (.A(net58),
    .B(_0420_),
    .X(_0277_));
 sky130_fd_sc_hd__a32o_1 _0860_ (.A1(net31),
    .A2(\timer_period_b[6] ),
    .A3(_0419_),
    .B1(net19),
    .B2(net35),
    .X(_0421_));
 sky130_fd_sc_hd__and2_1 _0861_ (.A(net58),
    .B(_0421_),
    .X(_0276_));
 sky130_fd_sc_hd__a32o_1 _0862_ (.A1(net31),
    .A2(\timer_period_b[5] ),
    .A3(_0419_),
    .B1(net19),
    .B2(net38),
    .X(_0422_));
 sky130_fd_sc_hd__and2_1 _0863_ (.A(net58),
    .B(_0422_),
    .X(_0275_));
 sky130_fd_sc_hd__a32o_1 _0864_ (.A1(net236),
    .A2(_0412_),
    .A3(_0419_),
    .B1(net19),
    .B2(_0410_),
    .X(_0274_));
 sky130_fd_sc_hd__a32o_1 _0865_ (.A1(net32),
    .A2(\timer_period_b[3] ),
    .A3(_0419_),
    .B1(net19),
    .B2(net42),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _0866_ (.A(net59),
    .B(_0423_),
    .X(_0273_));
 sky130_fd_sc_hd__a32o_1 _0867_ (.A1(net31),
    .A2(\timer_period_b[2] ),
    .A3(_0419_),
    .B1(net19),
    .B2(net44),
    .X(_0424_));
 sky130_fd_sc_hd__and2_1 _0868_ (.A(net59),
    .B(_0424_),
    .X(_0272_));
 sky130_fd_sc_hd__a32o_1 _0869_ (.A1(net32),
    .A2(_0349_),
    .A3(_0419_),
    .B1(net19),
    .B2(_0335_),
    .X(_0425_));
 sky130_fd_sc_hd__nand2_1 _0870_ (.A(net59),
    .B(_0425_),
    .Y(_0271_));
 sky130_fd_sc_hd__a32o_1 _0871_ (.A1(net31),
    .A2(\timer_period_b[0] ),
    .A3(_0419_),
    .B1(net19),
    .B2(net49),
    .X(_0426_));
 sky130_fd_sc_hd__and2_1 _0872_ (.A(net58),
    .B(_0426_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _0873_ (.A1(\timer_counter[11] ),
    .A2(_0346_),
    .B1(_0347_),
    .B2(\timer_counter[14] ),
    .X(_0427_));
 sky130_fd_sc_hd__xor2_1 _0874_ (.A(\timer_counter[4] ),
    .B(\timer_period_a[4] ),
    .X(_0428_));
 sky130_fd_sc_hd__a221o_1 _0875_ (.A1(_0332_),
    .A2(\timer_period_a[6] ),
    .B1(\timer_period_a[7] ),
    .B2(_0331_),
    .C1(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_1 _0876_ (.A(\timer_counter[1] ),
    .B(\timer_period_a[1] ),
    .Y(_0430_));
 sky130_fd_sc_hd__or2_1 _0877_ (.A(\timer_counter[1] ),
    .B(\timer_period_a[1] ),
    .X(_0431_));
 sky130_fd_sc_hd__xor2_1 _0878_ (.A(\timer_counter[15] ),
    .B(\timer_period_a[15] ),
    .X(_0432_));
 sky130_fd_sc_hd__a211o_1 _0879_ (.A1(_0430_),
    .A2(_0431_),
    .B1(_0432_),
    .C1(_0429_),
    .X(_0433_));
 sky130_fd_sc_hd__a211o_1 _0880_ (.A1(_0333_),
    .A2(\timer_period_a[2] ),
    .B1(_0427_),
    .C1(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__xor2_1 _0881_ (.A(\timer_counter[0] ),
    .B(\timer_period_a[0] ),
    .X(_0435_));
 sky130_fd_sc_hd__or2_1 _0882_ (.A(\timer_counter[3] ),
    .B(\timer_period_a[3] ),
    .X(_0436_));
 sky130_fd_sc_hd__nand2_1 _0883_ (.A(\timer_counter[3] ),
    .B(\timer_period_a[3] ),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _0884_ (.A(\timer_counter[5] ),
    .B(\timer_period_a[5] ),
    .Y(_0438_));
 sky130_fd_sc_hd__or2_1 _0885_ (.A(\timer_counter[5] ),
    .B(\timer_period_a[5] ),
    .X(_0439_));
 sky130_fd_sc_hd__a221o_1 _0886_ (.A1(_0436_),
    .A2(_0437_),
    .B1(_0438_),
    .B2(_0439_),
    .C1(_0435_),
    .X(_0440_));
 sky130_fd_sc_hd__a2bb2o_1 _0887_ (.A1_N(_0330_),
    .A2_N(\timer_period_a[8] ),
    .B1(\timer_period_a[10] ),
    .B2(_0328_),
    .X(_0441_));
 sky130_fd_sc_hd__a221o_1 _0888_ (.A1(\timer_counter[6] ),
    .A2(_0345_),
    .B1(\timer_period_a[8] ),
    .B2(_0330_),
    .C1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__or2_1 _0889_ (.A(\timer_counter[9] ),
    .B(\timer_period_a[9] ),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _0890_ (.A(\timer_counter[9] ),
    .B(\timer_period_a[9] ),
    .Y(_0444_));
 sky130_fd_sc_hd__a221o_1 _0891_ (.A1(_0327_),
    .A2(\timer_period_a[13] ),
    .B1(_0443_),
    .B2(_0444_),
    .C1(timer_phase),
    .X(_0445_));
 sky130_fd_sc_hd__o22a_1 _0892_ (.A1(_0331_),
    .A2(\timer_period_a[7] ),
    .B1(_0346_),
    .B2(\timer_counter[11] ),
    .X(_0446_));
 sky130_fd_sc_hd__o221a_1 _0893_ (.A1(_0333_),
    .A2(\timer_period_a[2] ),
    .B1(\timer_period_a[13] ),
    .B2(_0327_),
    .C1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__xnor2_1 _0894_ (.A(\timer_counter[12] ),
    .B(\timer_period_a[12] ),
    .Y(_0448_));
 sky130_fd_sc_hd__o221a_1 _0895_ (.A1(_0328_),
    .A2(\timer_period_a[10] ),
    .B1(_0347_),
    .B2(\timer_counter[14] ),
    .C1(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__and4bb_1 _0896_ (.A_N(_0442_),
    .B_N(_0445_),
    .C(_0447_),
    .D(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__or3b_1 _0897_ (.A(_0434_),
    .B(_0440_),
    .C_N(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__a21boi_2 _0898_ (.A1(_0405_),
    .A2(_0451_),
    .B1_N(_0362_),
    .Y(_0452_));
 sky130_fd_sc_hd__a21oi_1 _0899_ (.A1(timer_phase),
    .A2(_0452_),
    .B1(_0413_),
    .Y(_0453_));
 sky130_fd_sc_hd__o21a_1 _0900_ (.A1(net249),
    .A2(_0452_),
    .B1(_0453_),
    .X(_0269_));
 sky130_fd_sc_hd__or3b_4 _0901_ (.A(_0352_),
    .B(\fetch_prev_state[3] ),
    .C_N(\fetch_prev_state[2] ),
    .X(_0454_));
 sky130_fd_sc_hd__or3b_2 _0902_ (.A(_0454_),
    .B(\fetch_prev_state[1] ),
    .C_N(\fetch_prev_state[0] ),
    .X(_0455_));
 sky130_fd_sc_hd__or4b_1 _0903_ (.A(net33),
    .B(net35),
    .C(\stack[0] ),
    .D_N(net37),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _0904_ (.A(net38),
    .B(net39),
    .Y(_0457_));
 sky130_fd_sc_hd__nor3_1 _0905_ (.A(net33),
    .B(net35),
    .C(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__or3_1 _0906_ (.A(net33),
    .B(net36),
    .C(_0457_),
    .X(_0459_));
 sky130_fd_sc_hd__or4b_1 _0907_ (.A(net41),
    .B(_0455_),
    .C(net22),
    .D_N(_0456_),
    .X(_0460_));
 sky130_fd_sc_hd__or4b_1 _0908_ (.A(net33),
    .B(_0455_),
    .C(net35),
    .D_N(net37),
    .X(_0461_));
 sky130_fd_sc_hd__o31ai_1 _0909_ (.A1(net41),
    .A2(\stack[0] ),
    .A3(_0461_),
    .B1(_0397_),
    .Y(_0462_));
 sky130_fd_sc_hd__and3_1 _0910_ (.A(net30),
    .B(_0460_),
    .C(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_1 _0911_ (.A(net38),
    .B(net39),
    .Y(_0464_));
 sky130_fd_sc_hd__and2b_1 _0912_ (.A_N(net39),
    .B(net38),
    .X(_0465_));
 sky130_fd_sc_hd__nand2b_2 _0913_ (.A_N(net40),
    .B(net38),
    .Y(_0466_));
 sky130_fd_sc_hd__or2_1 _0914_ (.A(\stack[0] ),
    .B(net28),
    .X(_0467_));
 sky130_fd_sc_hd__and3b_1 _0915_ (.A_N(_0460_),
    .B(_0464_),
    .C(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__o21a_1 _0916_ (.A1(_0463_),
    .A2(_0468_),
    .B1(net61),
    .X(_0268_));
 sky130_fd_sc_hd__nor3b_2 _0917_ (.A(\fetch_prev_state[0] ),
    .B(_0454_),
    .C_N(\fetch_prev_state[1] ),
    .Y(_0469_));
 sky130_fd_sc_hd__nand2b_1 _0918_ (.A_N(\fetch_prev_state[0] ),
    .B(\fetch_prev_state[1] ),
    .Y(_0470_));
 sky130_fd_sc_hd__o21ba_1 _0919_ (.A1(_0454_),
    .A2(_0470_),
    .B1_N(_0397_),
    .X(_0471_));
 sky130_fd_sc_hd__and3_1 _0920_ (.A(net29),
    .B(\timer_period_a[15] ),
    .C(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(net34),
    .B(_0469_),
    .X(_0473_));
 sky130_fd_sc_hd__o21a_1 _0922_ (.A1(_0472_),
    .A2(_0473_),
    .B1(net51),
    .X(_0267_));
 sky130_fd_sc_hd__and3_1 _0923_ (.A(net30),
    .B(\timer_period_a[14] ),
    .C(_0471_),
    .X(_0474_));
 sky130_fd_sc_hd__and2_1 _0924_ (.A(net36),
    .B(_0469_),
    .X(_0475_));
 sky130_fd_sc_hd__o21a_1 _0925_ (.A1(_0474_),
    .A2(_0475_),
    .B1(net52),
    .X(_0266_));
 sky130_fd_sc_hd__and3_1 _0926_ (.A(net29),
    .B(\timer_period_a[13] ),
    .C(_0471_),
    .X(_0476_));
 sky130_fd_sc_hd__and2_1 _0927_ (.A(net37),
    .B(_0469_),
    .X(_0477_));
 sky130_fd_sc_hd__o21a_1 _0928_ (.A1(_0476_),
    .A2(_0477_),
    .B1(net51),
    .X(_0265_));
 sky130_fd_sc_hd__and3_1 _0929_ (.A(\timer_period_a[12] ),
    .B(_0412_),
    .C(_0471_),
    .X(_0478_));
 sky130_fd_sc_hd__a21o_1 _0930_ (.A1(_0410_),
    .A2(_0469_),
    .B1(_0478_),
    .X(_0264_));
 sky130_fd_sc_hd__and3_1 _0931_ (.A(net29),
    .B(\timer_period_a[11] ),
    .C(_0471_),
    .X(_0479_));
 sky130_fd_sc_hd__and2_1 _0932_ (.A(net41),
    .B(_0469_),
    .X(_0480_));
 sky130_fd_sc_hd__o21a_1 _0933_ (.A1(_0479_),
    .A2(_0480_),
    .B1(net51),
    .X(_0263_));
 sky130_fd_sc_hd__and3_1 _0934_ (.A(net29),
    .B(\timer_period_a[10] ),
    .C(_0471_),
    .X(_0481_));
 sky130_fd_sc_hd__and2_1 _0935_ (.A(net43),
    .B(_0469_),
    .X(_0482_));
 sky130_fd_sc_hd__o21a_1 _0936_ (.A1(_0481_),
    .A2(_0482_),
    .B1(net51),
    .X(_0262_));
 sky130_fd_sc_hd__and3_1 _0937_ (.A(net29),
    .B(\timer_period_a[9] ),
    .C(_0471_),
    .X(_0483_));
 sky130_fd_sc_hd__and2_1 _0938_ (.A(net45),
    .B(_0469_),
    .X(_0484_));
 sky130_fd_sc_hd__o21a_1 _0939_ (.A1(_0483_),
    .A2(_0484_),
    .B1(net51),
    .X(_0261_));
 sky130_fd_sc_hd__and3_1 _0940_ (.A(net29),
    .B(\timer_period_a[8] ),
    .C(_0471_),
    .X(_0485_));
 sky130_fd_sc_hd__and2_1 _0941_ (.A(net48),
    .B(_0469_),
    .X(_0486_));
 sky130_fd_sc_hd__o21a_1 _0942_ (.A1(_0485_),
    .A2(_0486_),
    .B1(net51),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_1 _0943_ (.A(\fetch_prev_state[1] ),
    .B(\fetch_prev_state[0] ),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_4 _0944_ (.A(_0454_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_2 _0945_ (.A(_0397_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__a32o_1 _0946_ (.A1(net31),
    .A2(\timer_period_a[7] ),
    .A3(_0489_),
    .B1(_0488_),
    .B2(net33),
    .X(_0490_));
 sky130_fd_sc_hd__and2_1 _0947_ (.A(net58),
    .B(_0490_),
    .X(_0259_));
 sky130_fd_sc_hd__a32o_1 _0948_ (.A1(net31),
    .A2(\timer_period_a[6] ),
    .A3(_0489_),
    .B1(_0488_),
    .B2(net35),
    .X(_0491_));
 sky130_fd_sc_hd__and2_1 _0949_ (.A(net58),
    .B(_0491_),
    .X(_0258_));
 sky130_fd_sc_hd__a32o_1 _0950_ (.A1(net32),
    .A2(\timer_period_a[5] ),
    .A3(_0489_),
    .B1(_0488_),
    .B2(net38),
    .X(_0492_));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(net59),
    .B(_0492_),
    .X(_0257_));
 sky130_fd_sc_hd__a32o_1 _0952_ (.A1(net219),
    .A2(_0412_),
    .A3(_0489_),
    .B1(_0488_),
    .B2(_0410_),
    .X(_0256_));
 sky130_fd_sc_hd__a32o_1 _0953_ (.A1(net32),
    .A2(\timer_period_a[3] ),
    .A3(_0489_),
    .B1(_0488_),
    .B2(net42),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _0954_ (.A(net59),
    .B(_0493_),
    .X(_0255_));
 sky130_fd_sc_hd__a32o_1 _0955_ (.A1(net31),
    .A2(\timer_period_a[2] ),
    .A3(_0489_),
    .B1(_0488_),
    .B2(net44),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _0956_ (.A(net58),
    .B(_0494_),
    .X(_0254_));
 sky130_fd_sc_hd__a32o_1 _0957_ (.A1(net32),
    .A2(\timer_period_a[1] ),
    .A3(_0489_),
    .B1(_0488_),
    .B2(\instr[1] ),
    .X(_0495_));
 sky130_fd_sc_hd__and2_1 _0958_ (.A(net59),
    .B(_0495_),
    .X(_0253_));
 sky130_fd_sc_hd__a32o_1 _0959_ (.A1(net32),
    .A2(_0344_),
    .A3(_0489_),
    .B1(_0488_),
    .B2(_0336_),
    .X(_0496_));
 sky130_fd_sc_hd__nand2_1 _0960_ (.A(net59),
    .B(_0496_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2b_1 _0961_ (.A_N(net34),
    .B(net36),
    .Y(_0497_));
 sky130_fd_sc_hd__nor4_1 _0962_ (.A(net37),
    .B(net39),
    .C(_0455_),
    .D(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__nor2_1 _0963_ (.A(_0397_),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__a32o_1 _0964_ (.A1(net29),
    .A2(\timer_clock_divisor[3] ),
    .A3(_0499_),
    .B1(net17),
    .B2(net41),
    .X(_0500_));
 sky130_fd_sc_hd__and2_1 _0965_ (.A(net53),
    .B(_0500_),
    .X(_0251_));
 sky130_fd_sc_hd__a32o_1 _0966_ (.A1(net29),
    .A2(\timer_clock_divisor[2] ),
    .A3(_0499_),
    .B1(net17),
    .B2(net43),
    .X(_0501_));
 sky130_fd_sc_hd__and2_1 _0967_ (.A(net53),
    .B(_0501_),
    .X(_0250_));
 sky130_fd_sc_hd__a32o_1 _0968_ (.A1(net29),
    .A2(\timer_clock_divisor[1] ),
    .A3(_0499_),
    .B1(net17),
    .B2(net45),
    .X(_0502_));
 sky130_fd_sc_hd__and2_1 _0969_ (.A(net53),
    .B(_0502_),
    .X(_0249_));
 sky130_fd_sc_hd__a32o_1 _0970_ (.A1(net29),
    .A2(\timer_clock_divisor[0] ),
    .A3(_0499_),
    .B1(net17),
    .B2(net48),
    .X(_0503_));
 sky130_fd_sc_hd__and2_1 _0971_ (.A(net53),
    .B(_0503_),
    .X(_0248_));
 sky130_fd_sc_hd__and3_1 _0972_ (.A(\timer_counter[2] ),
    .B(\timer_counter[1] ),
    .C(\timer_counter[0] ),
    .X(_0504_));
 sky130_fd_sc_hd__and4_1 _0973_ (.A(\timer_counter[8] ),
    .B(\timer_counter[7] ),
    .C(\timer_counter[6] ),
    .D(\timer_counter[3] ),
    .X(_0505_));
 sky130_fd_sc_hd__and4_1 _0974_ (.A(\timer_counter[5] ),
    .B(\timer_counter[4] ),
    .C(_0504_),
    .D(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_1 _0975_ (.A(_0362_),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__nor2_1 _0976_ (.A(_0329_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__and4_2 _0977_ (.A(\timer_counter[10] ),
    .B(\timer_counter[9] ),
    .C(_0362_),
    .D(_0506_),
    .X(_0509_));
 sky130_fd_sc_hd__inv_2 _0978_ (.A(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(net261),
    .B(_0509_),
    .Y(_0511_));
 sky130_fd_sc_hd__and3_1 _0980_ (.A(\timer_counter[12] ),
    .B(\timer_counter[11] ),
    .C(_0509_),
    .X(_0512_));
 sky130_fd_sc_hd__and4_1 _0981_ (.A(\timer_counter[13] ),
    .B(\timer_counter[12] ),
    .C(\timer_counter[11] ),
    .D(_0509_),
    .X(_0513_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_1 _0983_ (.A(\timer_counter[14] ),
    .B(_0513_),
    .Y(_0515_));
 sky130_fd_sc_hd__nor2_1 _0984_ (.A(_0413_),
    .B(_0452_),
    .Y(_0516_));
 sky130_fd_sc_hd__xnor2_1 _0985_ (.A(\timer_counter[15] ),
    .B(_0515_),
    .Y(_0517_));
 sky130_fd_sc_hd__and2_1 _0986_ (.A(net11),
    .B(_0517_),
    .X(_0247_));
 sky130_fd_sc_hd__o211a_1 _0987_ (.A1(\timer_counter[14] ),
    .A2(_0513_),
    .B1(_0515_),
    .C1(net11),
    .X(_0246_));
 sky130_fd_sc_hd__o211a_1 _0988_ (.A1(net237),
    .A2(_0512_),
    .B1(_0514_),
    .C1(net11),
    .X(_0245_));
 sky130_fd_sc_hd__a21o_1 _0989_ (.A1(\timer_counter[11] ),
    .A2(_0509_),
    .B1(\timer_counter[12] ),
    .X(_0518_));
 sky130_fd_sc_hd__and3b_1 _0990_ (.A_N(_0512_),
    .B(net11),
    .C(_0518_),
    .X(_0244_));
 sky130_fd_sc_hd__o211a_1 _0991_ (.A1(\timer_counter[11] ),
    .A2(_0509_),
    .B1(_0511_),
    .C1(net11),
    .X(_0243_));
 sky130_fd_sc_hd__o211a_1 _0992_ (.A1(net250),
    .A2(_0508_),
    .B1(_0510_),
    .C1(net11),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(_0329_),
    .B(_0507_),
    .Y(_0519_));
 sky130_fd_sc_hd__and3b_1 _0994_ (.A_N(_0508_),
    .B(net11),
    .C(_0519_),
    .X(_0241_));
 sky130_fd_sc_hd__and2_1 _0995_ (.A(\timer_counter[0] ),
    .B(_0362_),
    .X(_0520_));
 sky130_fd_sc_hd__and3_1 _0996_ (.A(\timer_counter[1] ),
    .B(\timer_counter[0] ),
    .C(_0362_),
    .X(_0521_));
 sky130_fd_sc_hd__and2_1 _0997_ (.A(_0362_),
    .B(_0504_),
    .X(_0522_));
 sky130_fd_sc_hd__and3_1 _0998_ (.A(\timer_counter[3] ),
    .B(_0362_),
    .C(_0504_),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _0999_ (.A(\timer_counter[4] ),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__and3_1 _1000_ (.A(\timer_counter[5] ),
    .B(\timer_counter[4] ),
    .C(_0523_),
    .X(_0525_));
 sky130_fd_sc_hd__and3_1 _1001_ (.A(\timer_counter[6] ),
    .B(\timer_counter[5] ),
    .C(_0524_),
    .X(_0526_));
 sky130_fd_sc_hd__and2_1 _1002_ (.A(\timer_counter[7] ),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__o211a_1 _1003_ (.A1(\timer_counter[8] ),
    .A2(_0527_),
    .B1(net12),
    .C1(_0507_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _1004_ (.A(\timer_counter[7] ),
    .B(_0526_),
    .X(_0528_));
 sky130_fd_sc_hd__and3b_1 _1005_ (.A_N(_0527_),
    .B(_0528_),
    .C(net11),
    .X(_0239_));
 sky130_fd_sc_hd__or2_1 _1006_ (.A(\timer_counter[6] ),
    .B(_0525_),
    .X(_0529_));
 sky130_fd_sc_hd__and3b_1 _1007_ (.A_N(_0526_),
    .B(_0529_),
    .C(net11),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _1008_ (.A(\timer_counter[5] ),
    .B(_0524_),
    .X(_0530_));
 sky130_fd_sc_hd__and3b_1 _1009_ (.A_N(_0525_),
    .B(_0530_),
    .C(net11),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(\timer_counter[4] ),
    .B(_0523_),
    .X(_0531_));
 sky130_fd_sc_hd__and3b_1 _1011_ (.A_N(_0524_),
    .B(_0531_),
    .C(net12),
    .X(_0236_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(\timer_counter[3] ),
    .B(_0522_),
    .X(_0532_));
 sky130_fd_sc_hd__and3b_1 _1013_ (.A_N(_0523_),
    .B(_0532_),
    .C(net12),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _1014_ (.A(\timer_counter[2] ),
    .B(_0521_),
    .X(_0533_));
 sky130_fd_sc_hd__and3b_1 _1015_ (.A_N(_0522_),
    .B(_0533_),
    .C(net12),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _1016_ (.A(\timer_counter[1] ),
    .B(_0520_),
    .X(_0534_));
 sky130_fd_sc_hd__and3b_1 _1017_ (.A_N(_0521_),
    .B(_0534_),
    .C(net12),
    .X(_0233_));
 sky130_fd_sc_hd__or2_1 _1018_ (.A(\timer_counter[0] ),
    .B(_0362_),
    .X(_0535_));
 sky130_fd_sc_hd__and3b_1 _1019_ (.A_N(_0520_),
    .B(_0535_),
    .C(net12),
    .X(_0232_));
 sky130_fd_sc_hd__nand3_1 _1020_ (.A(\timer_clock_counter[0] ),
    .B(\timer_clock_counter[1] ),
    .C(\timer_clock_counter[2] ),
    .Y(_0536_));
 sky130_fd_sc_hd__and4_1 _1021_ (.A(\timer_clock_counter[0] ),
    .B(\timer_clock_counter[1] ),
    .C(\timer_clock_counter[2] ),
    .D(\timer_clock_counter[3] ),
    .X(_0537_));
 sky130_fd_sc_hd__and3_1 _1022_ (.A(\timer_clock_counter[4] ),
    .B(\timer_clock_counter[5] ),
    .C(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__and4_1 _1023_ (.A(\timer_clock_counter[4] ),
    .B(\timer_clock_counter[5] ),
    .C(\timer_clock_counter[6] ),
    .D(_0537_),
    .X(_0539_));
 sky130_fd_sc_hd__and2_1 _1024_ (.A(\timer_clock_counter[7] ),
    .B(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__and3_1 _1025_ (.A(\timer_clock_counter[7] ),
    .B(\timer_clock_counter[8] ),
    .C(_0539_),
    .X(_0541_));
 sky130_fd_sc_hd__and2_1 _1026_ (.A(\timer_clock_counter[9] ),
    .B(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__and3_1 _1027_ (.A(\timer_clock_counter[10] ),
    .B(\timer_clock_counter[11] ),
    .C(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__and2_1 _1028_ (.A(\timer_clock_counter[12] ),
    .B(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__and3_1 _1029_ (.A(\timer_clock_counter[13] ),
    .B(\timer_clock_counter[14] ),
    .C(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__nor2_1 _1030_ (.A(_0362_),
    .B(_0413_),
    .Y(_0546_));
 sky130_fd_sc_hd__o21a_1 _1031_ (.A1(net214),
    .A2(_0545_),
    .B1(net15),
    .X(_0231_));
 sky130_fd_sc_hd__a31o_1 _1032_ (.A1(\timer_clock_counter[12] ),
    .A2(\timer_clock_counter[13] ),
    .A3(_0543_),
    .B1(\timer_clock_counter[14] ),
    .X(_0547_));
 sky130_fd_sc_hd__and3b_1 _1033_ (.A_N(_0545_),
    .B(net15),
    .C(_0547_),
    .X(_0230_));
 sky130_fd_sc_hd__o21ai_1 _1034_ (.A1(net217),
    .A2(_0544_),
    .B1(net15),
    .Y(_0548_));
 sky130_fd_sc_hd__a21oi_1 _1035_ (.A1(net217),
    .A2(_0544_),
    .B1(_0548_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ai_1 _1036_ (.A1(net238),
    .A2(_0543_),
    .B1(net15),
    .Y(_0549_));
 sky130_fd_sc_hd__nor2_1 _1037_ (.A(_0544_),
    .B(_0549_),
    .Y(_0228_));
 sky130_fd_sc_hd__a31o_1 _1038_ (.A1(\timer_clock_counter[9] ),
    .A2(\timer_clock_counter[10] ),
    .A3(_0541_),
    .B1(\timer_clock_counter[11] ),
    .X(_0550_));
 sky130_fd_sc_hd__and3b_1 _1039_ (.A_N(_0543_),
    .B(net15),
    .C(_0550_),
    .X(_0227_));
 sky130_fd_sc_hd__o21ai_1 _1040_ (.A1(net218),
    .A2(_0542_),
    .B1(net15),
    .Y(_0551_));
 sky130_fd_sc_hd__a21oi_1 _1041_ (.A1(net218),
    .A2(_0542_),
    .B1(_0551_),
    .Y(_0226_));
 sky130_fd_sc_hd__o21ai_1 _1042_ (.A1(net244),
    .A2(_0541_),
    .B1(net15),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_1 _1043_ (.A(_0542_),
    .B(_0552_),
    .Y(_0225_));
 sky130_fd_sc_hd__o21ai_1 _1044_ (.A1(net227),
    .A2(_0540_),
    .B1(net16),
    .Y(_0553_));
 sky130_fd_sc_hd__nor2_1 _1045_ (.A(_0541_),
    .B(_0553_),
    .Y(_0224_));
 sky130_fd_sc_hd__o21ai_1 _1046_ (.A1(net241),
    .A2(_0539_),
    .B1(net15),
    .Y(_0554_));
 sky130_fd_sc_hd__nor2_1 _1047_ (.A(_0540_),
    .B(_0554_),
    .Y(_0223_));
 sky130_fd_sc_hd__o21ai_1 _1048_ (.A1(net220),
    .A2(_0538_),
    .B1(net15),
    .Y(_0555_));
 sky130_fd_sc_hd__nor2_1 _1049_ (.A(_0539_),
    .B(_0555_),
    .Y(_0222_));
 sky130_fd_sc_hd__a21o_1 _1050_ (.A1(\timer_clock_counter[4] ),
    .A2(_0537_),
    .B1(\timer_clock_counter[5] ),
    .X(_0556_));
 sky130_fd_sc_hd__and3b_1 _1051_ (.A_N(_0538_),
    .B(net15),
    .C(_0556_),
    .X(_0221_));
 sky130_fd_sc_hd__o21ai_1 _1052_ (.A1(\timer_clock_counter[4] ),
    .A2(_0537_),
    .B1(net16),
    .Y(_0557_));
 sky130_fd_sc_hd__a21oi_1 _1053_ (.A1(net228),
    .A2(_0537_),
    .B1(_0557_),
    .Y(_0220_));
 sky130_fd_sc_hd__a31o_1 _1054_ (.A1(\timer_clock_counter[0] ),
    .A2(\timer_clock_counter[1] ),
    .A3(\timer_clock_counter[2] ),
    .B1(\timer_clock_counter[3] ),
    .X(_0558_));
 sky130_fd_sc_hd__and3b_1 _1055_ (.A_N(_0537_),
    .B(net16),
    .C(_0558_),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_1 _1056_ (.A1(\timer_clock_counter[0] ),
    .A2(\timer_clock_counter[1] ),
    .B1(\timer_clock_counter[2] ),
    .X(_0559_));
 sky130_fd_sc_hd__and3_1 _1057_ (.A(_0536_),
    .B(net16),
    .C(_0559_),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1058_ (.A1(\timer_clock_counter[0] ),
    .A2(\timer_clock_counter[1] ),
    .B1(net16),
    .Y(_0560_));
 sky130_fd_sc_hd__a21oi_1 _1059_ (.A1(net242),
    .A2(\timer_clock_counter[1] ),
    .B1(_0560_),
    .Y(_0217_));
 sky130_fd_sc_hd__and2b_1 _1060_ (.A_N(\timer_clock_counter[0] ),
    .B(net16),
    .X(_0216_));
 sky130_fd_sc_hd__nor2_1 _1061_ (.A(net35),
    .B(_0455_),
    .Y(_0561_));
 sky130_fd_sc_hd__or2_1 _1062_ (.A(net35),
    .B(_0455_),
    .X(_0562_));
 sky130_fd_sc_hd__or3b_1 _1063_ (.A(_0562_),
    .B(\stack[14] ),
    .C_N(_0457_),
    .X(_0563_));
 sky130_fd_sc_hd__a21o_1 _1064_ (.A1(_0457_),
    .A2(_0561_),
    .B1(\stack[15] ),
    .X(_0564_));
 sky130_fd_sc_hd__and3_1 _1065_ (.A(net61),
    .B(_0563_),
    .C(_0564_),
    .X(_0215_));
 sky130_fd_sc_hd__and2b_1 _1066_ (.A_N(\fetch_state[2] ),
    .B(\fetch_state[3] ),
    .X(_0565_));
 sky130_fd_sc_hd__nor2_1 _1067_ (.A(net50),
    .B(\fetch_state[0] ),
    .Y(_0566_));
 sky130_fd_sc_hd__or2_1 _1068_ (.A(net50),
    .B(\fetch_state[0] ),
    .X(_0567_));
 sky130_fd_sc_hd__and2b_1 _1069_ (.A_N(\fetch_state[3] ),
    .B(\fetch_state[2] ),
    .X(_0568_));
 sky130_fd_sc_hd__a21oi_2 _1070_ (.A1(_0567_),
    .A2(_0568_),
    .B1(_0565_),
    .Y(_0569_));
 sky130_fd_sc_hd__a21o_2 _1071_ (.A1(_0567_),
    .A2(_0568_),
    .B1(_0565_),
    .X(_0570_));
 sky130_fd_sc_hd__or2_1 _1072_ (.A(net36),
    .B(_0569_),
    .X(_0571_));
 sky130_fd_sc_hd__o211a_1 _1073_ (.A1(net34),
    .A2(net20),
    .B1(_0571_),
    .C1(net55),
    .X(_0214_));
 sky130_fd_sc_hd__or2_1 _1074_ (.A(net37),
    .B(_0569_),
    .X(_0572_));
 sky130_fd_sc_hd__o211a_1 _1075_ (.A1(net36),
    .A2(net20),
    .B1(_0572_),
    .C1(net55),
    .X(_0213_));
 sky130_fd_sc_hd__or2_1 _1076_ (.A(net39),
    .B(_0569_),
    .X(_0573_));
 sky130_fd_sc_hd__o211a_1 _1077_ (.A1(net37),
    .A2(net20),
    .B1(_0573_),
    .C1(net55),
    .X(_0212_));
 sky130_fd_sc_hd__or2_1 _1078_ (.A(net41),
    .B(_0569_),
    .X(_0574_));
 sky130_fd_sc_hd__o211a_1 _1079_ (.A1(net39),
    .A2(net20),
    .B1(_0574_),
    .C1(net55),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_1 _1080_ (.A(_0334_),
    .B(net20),
    .Y(_0575_));
 sky130_fd_sc_hd__o211a_1 _1081_ (.A1(net42),
    .A2(net20),
    .B1(_0575_),
    .C1(net61),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _1082_ (.A(_0335_),
    .B(_0570_),
    .Y(_0576_));
 sky130_fd_sc_hd__o211a_1 _1083_ (.A1(net44),
    .A2(net20),
    .B1(_0576_),
    .C1(net59),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _1084_ (.A(_0336_),
    .B(_0570_),
    .Y(_0577_));
 sky130_fd_sc_hd__o211a_1 _1085_ (.A1(net239),
    .A2(_0570_),
    .B1(_0577_),
    .C1(net59),
    .X(_0208_));
 sky130_fd_sc_hd__or2_1 _1086_ (.A(\uio_in_reg[3] ),
    .B(_0569_),
    .X(_0578_));
 sky130_fd_sc_hd__o211a_1 _1087_ (.A1(net47),
    .A2(net20),
    .B1(_0578_),
    .C1(net55),
    .X(_0207_));
 sky130_fd_sc_hd__nor2_1 _1088_ (.A(_0353_),
    .B(_0470_),
    .Y(_0579_));
 sky130_fd_sc_hd__or2_2 _1089_ (.A(_0353_),
    .B(_0470_),
    .X(_0580_));
 sky130_fd_sc_hd__or2_1 _1090_ (.A(\cycle_end_addr[7] ),
    .B(_0579_),
    .X(_0581_));
 sky130_fd_sc_hd__o211a_1 _1091_ (.A1(net34),
    .A2(_0580_),
    .B1(_0581_),
    .C1(net52),
    .X(_0206_));
 sky130_fd_sc_hd__or2_1 _1092_ (.A(\cycle_end_addr[6] ),
    .B(_0579_),
    .X(_0582_));
 sky130_fd_sc_hd__o211a_1 _1093_ (.A1(net36),
    .A2(_0580_),
    .B1(_0582_),
    .C1(net53),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _1094_ (.A(\cycle_end_addr[5] ),
    .B(_0579_),
    .X(_0583_));
 sky130_fd_sc_hd__o211a_1 _1095_ (.A1(net37),
    .A2(_0580_),
    .B1(_0583_),
    .C1(net53),
    .X(_0204_));
 sky130_fd_sc_hd__or2_1 _1096_ (.A(\cycle_end_addr[4] ),
    .B(_0579_),
    .X(_0584_));
 sky130_fd_sc_hd__o211a_1 _1097_ (.A1(net39),
    .A2(_0580_),
    .B1(_0584_),
    .C1(net52),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _1098_ (.A(\cycle_end_addr[3] ),
    .B(_0579_),
    .X(_0585_));
 sky130_fd_sc_hd__o211a_1 _1099_ (.A1(net41),
    .A2(_0580_),
    .B1(_0585_),
    .C1(net53),
    .X(_0202_));
 sky130_fd_sc_hd__or2_1 _1100_ (.A(\cycle_end_addr[2] ),
    .B(_0579_),
    .X(_0586_));
 sky130_fd_sc_hd__o211a_1 _1101_ (.A1(net43),
    .A2(_0580_),
    .B1(_0586_),
    .C1(net53),
    .X(_0201_));
 sky130_fd_sc_hd__or2_1 _1102_ (.A(net266),
    .B(_0579_),
    .X(_0587_));
 sky130_fd_sc_hd__o211a_1 _1103_ (.A1(net45),
    .A2(_0580_),
    .B1(_0587_),
    .C1(net53),
    .X(_0200_));
 sky130_fd_sc_hd__or2_1 _1104_ (.A(net248),
    .B(_0579_),
    .X(_0588_));
 sky130_fd_sc_hd__o211a_1 _1105_ (.A1(net48),
    .A2(_0580_),
    .B1(_0588_),
    .C1(net53),
    .X(_0199_));
 sky130_fd_sc_hd__nor2_1 _1106_ (.A(_0353_),
    .B(_0487_),
    .Y(_0589_));
 sky130_fd_sc_hd__or2_2 _1107_ (.A(_0353_),
    .B(_0487_),
    .X(_0590_));
 sky130_fd_sc_hd__or2_1 _1108_ (.A(net260),
    .B(_0589_),
    .X(_0591_));
 sky130_fd_sc_hd__o211a_1 _1109_ (.A1(net34),
    .A2(_0590_),
    .B1(_0591_),
    .C1(net55),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _1110_ (.A(net256),
    .B(_0589_),
    .X(_0592_));
 sky130_fd_sc_hd__o211a_1 _1111_ (.A1(net36),
    .A2(_0590_),
    .B1(_0592_),
    .C1(net55),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _1112_ (.A(net263),
    .B(_0589_),
    .X(_0593_));
 sky130_fd_sc_hd__o211a_1 _1113_ (.A1(net37),
    .A2(_0590_),
    .B1(_0593_),
    .C1(net55),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _1114_ (.A(net262),
    .B(_0589_),
    .X(_0594_));
 sky130_fd_sc_hd__o211a_1 _1115_ (.A1(net39),
    .A2(_0590_),
    .B1(_0594_),
    .C1(net55),
    .X(_0195_));
 sky130_fd_sc_hd__or2_1 _1116_ (.A(net264),
    .B(_0589_),
    .X(_0595_));
 sky130_fd_sc_hd__o211a_1 _1117_ (.A1(net42),
    .A2(_0590_),
    .B1(_0595_),
    .C1(net55),
    .X(_0194_));
 sky130_fd_sc_hd__or2_1 _1118_ (.A(net270),
    .B(_0589_),
    .X(_0596_));
 sky130_fd_sc_hd__o211a_1 _1119_ (.A1(net43),
    .A2(_0590_),
    .B1(_0596_),
    .C1(net56),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _1120_ (.A(net269),
    .B(_0589_),
    .X(_0597_));
 sky130_fd_sc_hd__o211a_1 _1121_ (.A1(net45),
    .A2(_0590_),
    .B1(_0597_),
    .C1(net54),
    .X(_0192_));
 sky130_fd_sc_hd__or2_1 _1122_ (.A(net258),
    .B(_0589_),
    .X(_0598_));
 sky130_fd_sc_hd__o211a_1 _1123_ (.A1(net47),
    .A2(_0590_),
    .B1(_0598_),
    .C1(net54),
    .X(_0191_));
 sky130_fd_sc_hd__and2b_1 _1124_ (.A_N(\fetch_state[0] ),
    .B(net50),
    .X(_0599_));
 sky130_fd_sc_hd__or2_2 _1125_ (.A(\fetch_state[3] ),
    .B(\fetch_state[2] ),
    .X(_0600_));
 sky130_fd_sc_hd__nor2_1 _1126_ (.A(_0599_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__or3_2 _1127_ (.A(\fetch_count[2] ),
    .B(\fetch_count[1] ),
    .C(\fetch_count[0] ),
    .X(_0602_));
 sky130_fd_sc_hd__o21ai_4 _1128_ (.A1(_0599_),
    .A2(_0600_),
    .B1(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_2 _1129_ (.A(net54),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__and4_1 _1130_ (.A(net54),
    .B(\cur_addr[0] ),
    .C(net20),
    .D(_0603_),
    .X(_0605_));
 sky130_fd_sc_hd__and3_1 _1131_ (.A(\cur_addr[2] ),
    .B(\cur_addr[1] ),
    .C(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__and2_1 _1132_ (.A(\cur_addr[3] ),
    .B(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__and3_1 _1133_ (.A(\cur_addr[5] ),
    .B(\cur_addr[4] ),
    .C(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__nand2_1 _1134_ (.A(\cur_addr[6] ),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__xnor2_1 _1135_ (.A(net222),
    .B(_0609_),
    .Y(_0190_));
 sky130_fd_sc_hd__xnor2_1 _1136_ (.A(_0338_),
    .B(_0608_),
    .Y(_0189_));
 sky130_fd_sc_hd__a21oi_1 _1137_ (.A1(\cur_addr[4] ),
    .A2(_0607_),
    .B1(net234),
    .Y(_0610_));
 sky130_fd_sc_hd__nor2_1 _1138_ (.A(_0608_),
    .B(net235),
    .Y(_0188_));
 sky130_fd_sc_hd__xnor2_1 _1139_ (.A(_0340_),
    .B(_0607_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _1140_ (.A(net231),
    .B(_0606_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _1141_ (.A(_0607_),
    .B(_0611_),
    .Y(_0186_));
 sky130_fd_sc_hd__a21oi_1 _1142_ (.A1(net271),
    .A2(_0605_),
    .B1(net232),
    .Y(_0612_));
 sky130_fd_sc_hd__nor2_1 _1143_ (.A(_0606_),
    .B(_0612_),
    .Y(_0185_));
 sky130_fd_sc_hd__xor2_1 _1144_ (.A(net246),
    .B(_0605_),
    .X(_0184_));
 sky130_fd_sc_hd__o21ba_1 _1145_ (.A1(_0569_),
    .A2(_0604_),
    .B1_N(\cur_addr[0] ),
    .X(_0613_));
 sky130_fd_sc_hd__nor2_1 _1146_ (.A(_0605_),
    .B(_0613_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand2_1 _1147_ (.A(net45),
    .B(net47),
    .Y(_0614_));
 sky130_fd_sc_hd__or4bb_1 _1148_ (.A(net33),
    .B(net35),
    .C_N(net37),
    .D_N(net40),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_2 _1149_ (.A(net45),
    .B(net47),
    .Y(_0616_));
 sky130_fd_sc_hd__and2b_2 _1150_ (.A_N(net49),
    .B(net46),
    .X(_0617_));
 sky130_fd_sc_hd__and3_1 _1151_ (.A(net46),
    .B(net47),
    .C(uo_out[3]),
    .X(_0618_));
 sky130_fd_sc_hd__and2b_2 _1152_ (.A_N(net45),
    .B(net47),
    .X(_0619_));
 sky130_fd_sc_hd__a21o_1 _1153_ (.A1(uo_out[2]),
    .A2(_0617_),
    .B1(net44),
    .X(_0620_));
 sky130_fd_sc_hd__a221o_1 _1154_ (.A1(uo_out[0]),
    .A2(_0616_),
    .B1(_0619_),
    .B2(uo_out[1]),
    .C1(_0618_),
    .X(_0621_));
 sky130_fd_sc_hd__mux4_1 _1155_ (.A0(uo_out[4]),
    .A1(uo_out[5]),
    .A2(uo_out[6]),
    .A3(uo_out[7]),
    .S0(net47),
    .S1(net45),
    .X(_0622_));
 sky130_fd_sc_hd__o22ai_1 _1156_ (.A1(_0620_),
    .A2(_0621_),
    .B1(_0622_),
    .B2(_0334_),
    .Y(_0623_));
 sky130_fd_sc_hd__a2bb2o_2 _1157_ (.A1_N(_0456_),
    .A2_N(_0623_),
    .B1(_0615_),
    .B2(\stack[0] ),
    .X(_0624_));
 sky130_fd_sc_hd__and2b_1 _1158_ (.A_N(net35),
    .B(net33),
    .X(_0625_));
 sky130_fd_sc_hd__nand2b_1 _1159_ (.A_N(net36),
    .B(net34),
    .Y(_0626_));
 sky130_fd_sc_hd__a31o_1 _1160_ (.A1(net43),
    .A2(net45),
    .A3(net47),
    .B1(uo_out[7]),
    .X(_0627_));
 sky130_fd_sc_hd__o311a_1 _1161_ (.A1(_0334_),
    .A2(_0614_),
    .A3(_0624_),
    .B1(net24),
    .C1(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__or3_1 _1162_ (.A(net33),
    .B(net37),
    .C(net40),
    .X(_0629_));
 sky130_fd_sc_hd__o211a_2 _1163_ (.A1(net41),
    .A2(net22),
    .B1(_0561_),
    .C1(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__a21bo_1 _1164_ (.A1(net41),
    .A2(net26),
    .B1_N(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__o221a_1 _1165_ (.A1(uo_out[7]),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0628_),
    .C1(net56),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _1166_ (.A(net43),
    .B(_0617_),
    .Y(_0632_));
 sky130_fd_sc_hd__a21o_1 _1167_ (.A1(net43),
    .A2(_0617_),
    .B1(uo_out[6]),
    .X(_0633_));
 sky130_fd_sc_hd__o211a_1 _1168_ (.A1(_0624_),
    .A2(_0632_),
    .B1(_0633_),
    .C1(net24),
    .X(_0634_));
 sky130_fd_sc_hd__o21ai_1 _1169_ (.A1(_0334_),
    .A2(net24),
    .B1(_0630_),
    .Y(_0635_));
 sky130_fd_sc_hd__o221a_1 _1170_ (.A1(uo_out[6]),
    .A2(_0630_),
    .B1(_0634_),
    .B2(_0635_),
    .C1(net56),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _1171_ (.A(net43),
    .B(_0619_),
    .Y(_0636_));
 sky130_fd_sc_hd__mux2_1 _1172_ (.A0(_0624_),
    .A1(uo_out[5]),
    .S(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _1173_ (.A0(net46),
    .A1(_0637_),
    .S(net24),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _1174_ (.A0(uo_out[5]),
    .A1(_0638_),
    .S(_0630_),
    .X(_0639_));
 sky130_fd_sc_hd__and2_1 _1175_ (.A(net56),
    .B(_0639_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _1176_ (.A(net44),
    .B(_0616_),
    .Y(_0640_));
 sky130_fd_sc_hd__mux2_1 _1177_ (.A0(_0624_),
    .A1(uo_out[4]),
    .S(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(net48),
    .A1(_0641_),
    .S(net24),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _1179_ (.A0(uo_out[4]),
    .A1(_0642_),
    .S(_0630_),
    .X(_0643_));
 sky130_fd_sc_hd__and2_1 _1180_ (.A(net56),
    .B(_0643_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _1181_ (.A0(\fetch_state[3] ),
    .A1(net216),
    .S(_0604_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(\fetch_state[2] ),
    .A1(net225),
    .S(_0604_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _1183_ (.A0(net50),
    .A1(net268),
    .S(_0604_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(net255),
    .A1(\fetch_prev_state[0] ),
    .S(_0604_),
    .X(_0175_));
 sky130_fd_sc_hd__nand2_1 _1185_ (.A(\fetch_state[3] ),
    .B(\fetch_state[2] ),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2_1 _1186_ (.A(_0567_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__or2_1 _1187_ (.A(_0567_),
    .B(_0644_),
    .X(_0646_));
 sky130_fd_sc_hd__nand2_1 _1188_ (.A(net50),
    .B(\fetch_state[0] ),
    .Y(_0647_));
 sky130_fd_sc_hd__or2_1 _1189_ (.A(_0600_),
    .B(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__nand2b_1 _1190_ (.A_N(net50),
    .B(\fetch_state[0] ),
    .Y(_0649_));
 sky130_fd_sc_hd__o21ai_1 _1191_ (.A1(net50),
    .A2(_0644_),
    .B1(_0648_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _1192_ (.A(net20),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__or2_1 _1193_ (.A(\fetch_count[0] ),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or2_1 _1194_ (.A(\fetch_count[1] ),
    .B(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__nand2_1 _1195_ (.A(net251),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__o211ai_1 _1196_ (.A1(_0602_),
    .A2(_0651_),
    .B1(_0654_),
    .C1(net54),
    .Y(_0174_));
 sky130_fd_sc_hd__nand2_1 _1197_ (.A(net54),
    .B(_0653_),
    .Y(_0655_));
 sky130_fd_sc_hd__a21o_1 _1198_ (.A1(\fetch_count[1] ),
    .A2(_0652_),
    .B1(_0655_),
    .X(_0173_));
 sky130_fd_sc_hd__nand2_1 _1199_ (.A(net54),
    .B(_0652_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21o_1 _1200_ (.A1(\fetch_count[0] ),
    .A2(_0651_),
    .B1(_0656_),
    .X(_0172_));
 sky130_fd_sc_hd__or4_2 _1201_ (.A(net42),
    .B(net43),
    .C(_0464_),
    .D(_0497_),
    .X(_0657_));
 sky130_fd_sc_hd__inv_2 _1202_ (.A(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__nand2_1 _1203_ (.A(_0619_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__and3b_1 _1204_ (.A_N(net50),
    .B(\fetch_state[0] ),
    .C(_0568_),
    .X(_0660_));
 sky130_fd_sc_hd__or4_1 _1205_ (.A(\cur_addr[3] ),
    .B(\cur_addr[2] ),
    .C(\cur_addr[1] ),
    .D(\cur_addr[0] ),
    .X(_0661_));
 sky130_fd_sc_hd__or4_1 _1206_ (.A(\cur_addr[7] ),
    .B(\cur_addr[6] ),
    .C(\cur_addr[5] ),
    .D(\cur_addr[4] ),
    .X(_0662_));
 sky130_fd_sc_hd__nor2_1 _1207_ (.A(_0661_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2b_1 _1208_ (.A_N(\cycle_end_addr[1] ),
    .B(\cur_addr[1] ),
    .Y(_0664_));
 sky130_fd_sc_hd__and2b_1 _1209_ (.A_N(\cur_addr[1] ),
    .B(\cycle_end_addr[1] ),
    .X(_0665_));
 sky130_fd_sc_hd__nand2b_1 _1210_ (.A_N(\cycle_end_addr[0] ),
    .B(\cur_addr[0] ),
    .Y(_0666_));
 sky130_fd_sc_hd__a221o_1 _1211_ (.A1(\cycle_end_addr[2] ),
    .A2(_0342_),
    .B1(_0664_),
    .B2(_0666_),
    .C1(_0665_),
    .X(_0667_));
 sky130_fd_sc_hd__o22a_1 _1212_ (.A1(\cycle_end_addr[3] ),
    .A2(_0341_),
    .B1(_0342_),
    .B2(\cycle_end_addr[2] ),
    .X(_0668_));
 sky130_fd_sc_hd__a22o_1 _1213_ (.A1(\cycle_end_addr[4] ),
    .A2(_0340_),
    .B1(_0341_),
    .B2(\cycle_end_addr[3] ),
    .X(_0669_));
 sky130_fd_sc_hd__a21o_1 _1214_ (.A1(_0667_),
    .A2(_0668_),
    .B1(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__o22a_1 _1215_ (.A1(\cycle_end_addr[5] ),
    .A2(_0339_),
    .B1(_0340_),
    .B2(\cycle_end_addr[4] ),
    .X(_0671_));
 sky130_fd_sc_hd__a22o_1 _1216_ (.A1(\cycle_end_addr[6] ),
    .A2(_0338_),
    .B1(_0339_),
    .B2(\cycle_end_addr[5] ),
    .X(_0672_));
 sky130_fd_sc_hd__a21o_1 _1217_ (.A1(_0670_),
    .A2(_0671_),
    .B1(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__o22a_1 _1218_ (.A1(\cycle_end_addr[7] ),
    .A2(_0337_),
    .B1(_0338_),
    .B2(\cycle_end_addr[6] ),
    .X(_0674_));
 sky130_fd_sc_hd__a22o_1 _1219_ (.A1(\cycle_end_addr[7] ),
    .A2(_0337_),
    .B1(_0673_),
    .B2(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__nand2b_1 _1220_ (.A_N(_0663_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__and3b_1 _1221_ (.A_N(_0663_),
    .B(_0675_),
    .C(_0660_),
    .X(_0677_));
 sky130_fd_sc_hd__or4_1 _1222_ (.A(\cycle_start_addr[3] ),
    .B(\cycle_start_addr[2] ),
    .C(\cycle_start_addr[1] ),
    .D(\cycle_start_addr[0] ),
    .X(_0678_));
 sky130_fd_sc_hd__or4_1 _1223_ (.A(\cycle_start_addr[7] ),
    .B(\cycle_start_addr[6] ),
    .C(\cycle_start_addr[5] ),
    .D(\cycle_start_addr[4] ),
    .X(_0679_));
 sky130_fd_sc_hd__nor2_1 _1224_ (.A(_0678_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__a32o_1 _1225_ (.A1(net50),
    .A2(\fetch_state[0] ),
    .A3(_0565_),
    .B1(_0645_),
    .B2(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__o211ai_1 _1226_ (.A1(_0644_),
    .A2(_0649_),
    .B1(_0648_),
    .C1(_0603_),
    .Y(_0682_));
 sky130_fd_sc_hd__a211o_1 _1227_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0681_),
    .C1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__a31o_1 _1228_ (.A1(_0619_),
    .A2(_0658_),
    .A3(_0677_),
    .B1(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__o211a_1 _1229_ (.A1(\fetch_state[3] ),
    .A2(_0603_),
    .B1(_0684_),
    .C1(net57),
    .X(_0171_));
 sky130_fd_sc_hd__a32o_1 _1230_ (.A1(_0565_),
    .A2(_0567_),
    .A3(_0647_),
    .B1(_0568_),
    .B2(net50),
    .X(_0685_));
 sky130_fd_sc_hd__nor2_1 _1231_ (.A(_0646_),
    .B(_0680_),
    .Y(_0686_));
 sky130_fd_sc_hd__a2111o_1 _1232_ (.A1(_0659_),
    .A2(_0677_),
    .B1(_0682_),
    .C1(_0685_),
    .D1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__o211a_1 _1233_ (.A1(net267),
    .A2(_0603_),
    .B1(_0687_),
    .C1(net54),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _1234_ (.A(_0568_),
    .B(_0599_),
    .X(_0688_));
 sky130_fd_sc_hd__nor2_1 _1235_ (.A(_0600_),
    .B(_0649_),
    .Y(_0689_));
 sky130_fd_sc_hd__or4b_1 _1236_ (.A(_0681_),
    .B(_0688_),
    .C(_0689_),
    .D_N(_0603_),
    .X(_0690_));
 sky130_fd_sc_hd__a31o_1 _1237_ (.A1(_0616_),
    .A2(_0658_),
    .A3(_0677_),
    .B1(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__o211a_1 _1238_ (.A1(net215),
    .A2(_0603_),
    .B1(_0691_),
    .C1(net57),
    .X(_0169_));
 sky130_fd_sc_hd__o31a_1 _1239_ (.A1(net46),
    .A2(_0657_),
    .A3(_0676_),
    .B1(_0660_),
    .X(_0692_));
 sky130_fd_sc_hd__a2111o_1 _1240_ (.A1(\fetch_state[3] ),
    .A2(_0566_),
    .B1(_0601_),
    .C1(_0602_),
    .D1(_0685_),
    .X(_0693_));
 sky130_fd_sc_hd__o221a_1 _1241_ (.A1(\fetch_state[0] ),
    .A2(_0603_),
    .B1(_0692_),
    .B2(_0693_),
    .C1(net54),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _1242_ (.A(_0325_),
    .B(net230),
    .X(_0167_));
 sky130_fd_sc_hd__or4_1 _1243_ (.A(\timer_period_b[1] ),
    .B(\timer_period_b[2] ),
    .C(\timer_period_b[3] ),
    .D(\timer_period_b[4] ),
    .X(_0694_));
 sky130_fd_sc_hd__or3_1 _1244_ (.A(timer_mode),
    .B(\timer_period_b[0] ),
    .C(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__or4_1 _1245_ (.A(\timer_period_b[9] ),
    .B(\timer_period_b[10] ),
    .C(\timer_period_b[11] ),
    .D(\timer_period_b[12] ),
    .X(_0696_));
 sky130_fd_sc_hd__or4_1 _1246_ (.A(\timer_period_b[5] ),
    .B(\timer_period_b[6] ),
    .C(\timer_period_b[7] ),
    .D(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__or4_1 _1247_ (.A(\timer_period_b[8] ),
    .B(\timer_period_b[13] ),
    .C(\timer_period_b[14] ),
    .D(\timer_period_b[15] ),
    .X(_0698_));
 sky130_fd_sc_hd__or4_1 _1248_ (.A(_0405_),
    .B(_0695_),
    .C(_0697_),
    .D(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__a21o_1 _1249_ (.A1(_0452_),
    .A2(_0699_),
    .B1(timer_out),
    .X(_0700_));
 sky130_fd_sc_hd__o211ai_1 _1250_ (.A1(timer_out),
    .A2(_0396_),
    .B1(_0452_),
    .C1(_0699_),
    .Y(_0701_));
 sky130_fd_sc_hd__and3_1 _1251_ (.A(_0412_),
    .B(_0700_),
    .C(_0701_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _1252_ (.A0(\cycle_start_addr[0] ),
    .A1(\cycle_start_addr[1] ),
    .S(\fetch_count[0] ),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _1253_ (.A0(\cycle_start_addr[2] ),
    .A1(\cycle_start_addr[3] ),
    .S(\fetch_count[0] ),
    .X(_0703_));
 sky130_fd_sc_hd__a21bo_1 _1254_ (.A1(_0645_),
    .A2(_0703_),
    .B1_N(\fetch_count[1] ),
    .X(_0704_));
 sky130_fd_sc_hd__o311a_1 _1255_ (.A1(\fetch_count[1] ),
    .A2(_0646_),
    .A3(_0702_),
    .B1(_0704_),
    .C1(_0343_),
    .X(_0705_));
 sky130_fd_sc_hd__mux4_1 _1256_ (.A0(\cycle_start_addr[4] ),
    .A1(\cycle_start_addr[5] ),
    .A2(\cycle_start_addr[6] ),
    .A3(\cycle_start_addr[7] ),
    .S0(\fetch_count[0] ),
    .S1(\fetch_count[1] ),
    .X(_0706_));
 sky130_fd_sc_hd__or3b_1 _1257_ (.A(_0343_),
    .B(_0646_),
    .C_N(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_1 _1258_ (.A(_0650_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__o221a_1 _1259_ (.A1(net221),
    .A2(_0650_),
    .B1(_0705_),
    .B2(_0708_),
    .C1(net57),
    .X(_0165_));
 sky130_fd_sc_hd__nand2_1 _1260_ (.A(net41),
    .B(_0623_),
    .Y(_0709_));
 sky130_fd_sc_hd__a311o_1 _1261_ (.A1(net46),
    .A2(net49),
    .A3(\ui_in_reg[7] ),
    .B1(_0334_),
    .C1(net42),
    .X(_0710_));
 sky130_fd_sc_hd__a22o_1 _1262_ (.A1(\ui_in_reg[4] ),
    .A2(_0616_),
    .B1(_0617_),
    .B2(\ui_in_reg[6] ),
    .X(_0711_));
 sky130_fd_sc_hd__a211o_1 _1263_ (.A1(\ui_in_reg[5] ),
    .A2(_0619_),
    .B1(_0710_),
    .C1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__and3_1 _1264_ (.A(net46),
    .B(net49),
    .C(\ui_in_reg[3] ),
    .X(_0713_));
 sky130_fd_sc_hd__a221o_1 _1265_ (.A1(\ui_in_reg[0] ),
    .A2(_0616_),
    .B1(_0619_),
    .B2(\ui_in_reg[1] ),
    .C1(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__a2111o_1 _1266_ (.A1(\ui_in_reg[2] ),
    .A2(_0617_),
    .B1(_0714_),
    .C1(net44),
    .D1(net42),
    .X(_0715_));
 sky130_fd_sc_hd__and3_1 _1267_ (.A(net21),
    .B(_0712_),
    .C(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__a221o_1 _1268_ (.A1(\stack[1] ),
    .A2(_0458_),
    .B1(_0709_),
    .B2(_0716_),
    .C1(net26),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _1269_ (.A0(net41),
    .A1(net44),
    .S(\stack[0] ),
    .X(_0718_));
 sky130_fd_sc_hd__and2b_1 _1270_ (.A_N(\stack[1] ),
    .B(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _1271_ (.A0(net46),
    .A1(net47),
    .S(\stack[0] ),
    .X(_0720_));
 sky130_fd_sc_hd__a211o_1 _1272_ (.A1(\stack[1] ),
    .A2(_0720_),
    .B1(_0719_),
    .C1(net24),
    .X(_0721_));
 sky130_fd_sc_hd__a21o_1 _1273_ (.A1(_0717_),
    .A2(_0721_),
    .B1(_0562_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_1 _1274_ (.A1(\stack[0] ),
    .A2(_0561_),
    .B1(_0722_),
    .C1(net61),
    .X(_0164_));
 sky130_fd_sc_hd__a21oi_2 _1275_ (.A1(net33),
    .A2(net40),
    .B1(_0562_),
    .Y(_0723_));
 sky130_fd_sc_hd__a21o_1 _1276_ (.A1(net33),
    .A2(net40),
    .B1(_0562_),
    .X(_0724_));
 sky130_fd_sc_hd__or2_1 _1277_ (.A(\stack[13] ),
    .B(net28),
    .X(_0725_));
 sky130_fd_sc_hd__o211a_1 _1278_ (.A1(\stack[15] ),
    .A2(net27),
    .B1(net25),
    .C1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _1279_ (.A0(\stack[15] ),
    .A1(\stack[13] ),
    .S(net21),
    .X(_0727_));
 sky130_fd_sc_hd__a211o_1 _1280_ (.A1(net23),
    .A2(_0727_),
    .B1(_0726_),
    .C1(net13),
    .X(_0728_));
 sky130_fd_sc_hd__o211a_1 _1281_ (.A1(net245),
    .A2(net14),
    .B1(_0728_),
    .C1(net60),
    .X(_0163_));
 sky130_fd_sc_hd__or2_1 _1282_ (.A(\stack[12] ),
    .B(net28),
    .X(_0729_));
 sky130_fd_sc_hd__o211a_1 _1283_ (.A1(\stack[14] ),
    .A2(net27),
    .B1(net25),
    .C1(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(\stack[14] ),
    .A1(\stack[12] ),
    .S(net21),
    .X(_0731_));
 sky130_fd_sc_hd__a211o_1 _1285_ (.A1(net23),
    .A2(_0731_),
    .B1(_0730_),
    .C1(net13),
    .X(_0732_));
 sky130_fd_sc_hd__o211a_1 _1286_ (.A1(net252),
    .A2(net14),
    .B1(_0732_),
    .C1(net60),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _1287_ (.A(\stack[11] ),
    .B(net28),
    .X(_0733_));
 sky130_fd_sc_hd__o211a_1 _1288_ (.A1(\stack[13] ),
    .A2(net27),
    .B1(net26),
    .C1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _1289_ (.A0(\stack[13] ),
    .A1(\stack[11] ),
    .S(net21),
    .X(_0735_));
 sky130_fd_sc_hd__a211o_1 _1290_ (.A1(net23),
    .A2(_0735_),
    .B1(_0734_),
    .C1(_0724_),
    .X(_0736_));
 sky130_fd_sc_hd__o211a_1 _1291_ (.A1(net257),
    .A2(net14),
    .B1(_0736_),
    .C1(net60),
    .X(_0161_));
 sky130_fd_sc_hd__or2_1 _1292_ (.A(\stack[10] ),
    .B(net28),
    .X(_0737_));
 sky130_fd_sc_hd__o211a_1 _1293_ (.A1(\stack[12] ),
    .A2(net27),
    .B1(net25),
    .C1(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _1294_ (.A0(\stack[12] ),
    .A1(\stack[10] ),
    .S(net22),
    .X(_0739_));
 sky130_fd_sc_hd__a211o_1 _1295_ (.A1(net23),
    .A2(_0739_),
    .B1(_0738_),
    .C1(_0724_),
    .X(_0740_));
 sky130_fd_sc_hd__o211a_1 _1296_ (.A1(net254),
    .A2(net14),
    .B1(_0740_),
    .C1(net60),
    .X(_0160_));
 sky130_fd_sc_hd__or2_1 _1297_ (.A(\stack[9] ),
    .B(net28),
    .X(_0741_));
 sky130_fd_sc_hd__o211a_1 _1298_ (.A1(\stack[11] ),
    .A2(_0466_),
    .B1(net25),
    .C1(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _1299_ (.A0(\stack[11] ),
    .A1(\stack[9] ),
    .S(net22),
    .X(_0743_));
 sky130_fd_sc_hd__a211o_1 _1300_ (.A1(_0626_),
    .A2(_0743_),
    .B1(_0742_),
    .C1(_0724_),
    .X(_0744_));
 sky130_fd_sc_hd__o211a_1 _1301_ (.A1(net265),
    .A2(_0723_),
    .B1(_0744_),
    .C1(net60),
    .X(_0159_));
 sky130_fd_sc_hd__or2_1 _1302_ (.A(\stack[8] ),
    .B(_0465_),
    .X(_0745_));
 sky130_fd_sc_hd__o211a_1 _1303_ (.A1(\stack[10] ),
    .A2(_0466_),
    .B1(net25),
    .C1(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _1304_ (.A0(\stack[10] ),
    .A1(\stack[8] ),
    .S(net22),
    .X(_0747_));
 sky130_fd_sc_hd__a211o_1 _1305_ (.A1(net24),
    .A2(_0747_),
    .B1(_0746_),
    .C1(_0724_),
    .X(_0748_));
 sky130_fd_sc_hd__o211a_1 _1306_ (.A1(net253),
    .A2(_0723_),
    .B1(_0748_),
    .C1(net60),
    .X(_0158_));
 sky130_fd_sc_hd__or2_1 _1307_ (.A(\stack[7] ),
    .B(_0465_),
    .X(_0749_));
 sky130_fd_sc_hd__o211a_1 _1308_ (.A1(\stack[9] ),
    .A2(net27),
    .B1(net25),
    .C1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _1309_ (.A0(\stack[9] ),
    .A1(\stack[7] ),
    .S(net21),
    .X(_0751_));
 sky130_fd_sc_hd__a211o_1 _1310_ (.A1(net24),
    .A2(_0751_),
    .B1(_0750_),
    .C1(net13),
    .X(_0752_));
 sky130_fd_sc_hd__o211a_1 _1311_ (.A1(net259),
    .A2(_0723_),
    .B1(_0752_),
    .C1(net60),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _1312_ (.A(\stack[6] ),
    .B(net28),
    .X(_0753_));
 sky130_fd_sc_hd__o211a_1 _1313_ (.A1(\stack[8] ),
    .A2(net27),
    .B1(net25),
    .C1(_0753_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _1314_ (.A0(\stack[8] ),
    .A1(\stack[6] ),
    .S(net21),
    .X(_0287_));
 sky130_fd_sc_hd__a211o_1 _1315_ (.A1(net23),
    .A2(_0287_),
    .B1(_0286_),
    .C1(net13),
    .X(_0288_));
 sky130_fd_sc_hd__o211a_1 _1316_ (.A1(\stack[7] ),
    .A2(_0723_),
    .B1(_0288_),
    .C1(net60),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _1317_ (.A(\stack[5] ),
    .B(_0465_),
    .X(_0289_));
 sky130_fd_sc_hd__o211a_1 _1318_ (.A1(\stack[7] ),
    .A2(_0466_),
    .B1(net26),
    .C1(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1319_ (.A0(\stack[7] ),
    .A1(\stack[5] ),
    .S(net21),
    .X(_0291_));
 sky130_fd_sc_hd__a211o_1 _1320_ (.A1(net23),
    .A2(_0291_),
    .B1(_0290_),
    .C1(net13),
    .X(_0292_));
 sky130_fd_sc_hd__o211a_1 _1321_ (.A1(\stack[6] ),
    .A2(net14),
    .B1(_0292_),
    .C1(net60),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _1322_ (.A(\stack[4] ),
    .B(_0465_),
    .X(_0293_));
 sky130_fd_sc_hd__o211a_1 _1323_ (.A1(\stack[6] ),
    .A2(_0466_),
    .B1(net25),
    .C1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(\stack[6] ),
    .A1(\stack[4] ),
    .S(net21),
    .X(_0295_));
 sky130_fd_sc_hd__a211o_1 _1325_ (.A1(net23),
    .A2(_0295_),
    .B1(_0294_),
    .C1(net13),
    .X(_0296_));
 sky130_fd_sc_hd__o211a_1 _1326_ (.A1(\stack[5] ),
    .A2(net14),
    .B1(_0296_),
    .C1(net62),
    .X(_0154_));
 sky130_fd_sc_hd__or2_1 _1327_ (.A(\stack[3] ),
    .B(net28),
    .X(_0297_));
 sky130_fd_sc_hd__o211a_1 _1328_ (.A1(\stack[5] ),
    .A2(net27),
    .B1(net25),
    .C1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _1329_ (.A0(\stack[5] ),
    .A1(\stack[3] ),
    .S(net21),
    .X(_0299_));
 sky130_fd_sc_hd__a211o_1 _1330_ (.A1(net23),
    .A2(_0299_),
    .B1(_0298_),
    .C1(net13),
    .X(_0300_));
 sky130_fd_sc_hd__o211a_1 _1331_ (.A1(\stack[4] ),
    .A2(net14),
    .B1(_0300_),
    .C1(net62),
    .X(_0153_));
 sky130_fd_sc_hd__or2_1 _1332_ (.A(\stack[2] ),
    .B(net28),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_1 _1333_ (.A1(\stack[4] ),
    .A2(net27),
    .B1(net25),
    .C1(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _1334_ (.A0(\stack[4] ),
    .A1(\stack[2] ),
    .S(net21),
    .X(_0303_));
 sky130_fd_sc_hd__a211o_1 _1335_ (.A1(net23),
    .A2(_0303_),
    .B1(_0302_),
    .C1(net13),
    .X(_0304_));
 sky130_fd_sc_hd__o211a_1 _1336_ (.A1(\stack[3] ),
    .A2(net14),
    .B1(_0304_),
    .C1(net60),
    .X(_0152_));
 sky130_fd_sc_hd__or2_1 _1337_ (.A(\stack[1] ),
    .B(net28),
    .X(_0305_));
 sky130_fd_sc_hd__o211a_1 _1338_ (.A1(\stack[3] ),
    .A2(net27),
    .B1(net26),
    .C1(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(\stack[3] ),
    .A1(\stack[1] ),
    .S(net22),
    .X(_0307_));
 sky130_fd_sc_hd__a211o_1 _1340_ (.A1(net23),
    .A2(_0307_),
    .B1(_0306_),
    .C1(net13),
    .X(_0308_));
 sky130_fd_sc_hd__o211a_1 _1341_ (.A1(\stack[2] ),
    .A2(net14),
    .B1(_0308_),
    .C1(net61),
    .X(_0151_));
 sky130_fd_sc_hd__o211a_1 _1342_ (.A1(\stack[2] ),
    .A2(net27),
    .B1(_0467_),
    .C1(net26),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _1343_ (.A0(\stack[0] ),
    .A1(\stack[2] ),
    .S(_0458_),
    .X(_0310_));
 sky130_fd_sc_hd__a211o_1 _1344_ (.A1(net24),
    .A2(_0310_),
    .B1(_0309_),
    .C1(net13),
    .X(_0311_));
 sky130_fd_sc_hd__o211a_1 _1345_ (.A1(\stack[1] ),
    .A2(net14),
    .B1(_0311_),
    .C1(net61),
    .X(_0150_));
 sky130_fd_sc_hd__or4_1 _1346_ (.A(net38),
    .B(_0411_),
    .C(_0455_),
    .D(_0497_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _1347_ (.A0(net48),
    .A1(net229),
    .S(_0312_),
    .X(_0149_));
 sky130_fd_sc_hd__and4bb_2 _1348_ (.A_N(net43),
    .B_N(_0455_),
    .C(_0458_),
    .D(net42),
    .X(_0313_));
 sky130_fd_sc_hd__and3_1 _1349_ (.A(net46),
    .B(net47),
    .C(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(uo_out[3]),
    .A1(_0624_),
    .S(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__and2_1 _1351_ (.A(net61),
    .B(_0315_),
    .X(_0148_));
 sky130_fd_sc_hd__nand2_1 _1352_ (.A(_0617_),
    .B(_0313_),
    .Y(_0316_));
 sky130_fd_sc_hd__a21o_1 _1353_ (.A1(_0617_),
    .A2(_0313_),
    .B1(uo_out[2]),
    .X(_0317_));
 sky130_fd_sc_hd__o211a_1 _1354_ (.A1(_0624_),
    .A2(_0316_),
    .B1(_0317_),
    .C1(net61),
    .X(_0147_));
 sky130_fd_sc_hd__nand2_1 _1355_ (.A(_0619_),
    .B(_0313_),
    .Y(_0318_));
 sky130_fd_sc_hd__a21o_1 _1356_ (.A1(_0619_),
    .A2(_0313_),
    .B1(uo_out[1]),
    .X(_0319_));
 sky130_fd_sc_hd__o211a_1 _1357_ (.A1(_0624_),
    .A2(_0318_),
    .B1(_0319_),
    .C1(net61),
    .X(_0146_));
 sky130_fd_sc_hd__nand2_1 _1358_ (.A(_0616_),
    .B(_0313_),
    .Y(_0320_));
 sky130_fd_sc_hd__a21o_1 _1359_ (.A1(_0616_),
    .A2(_0313_),
    .B1(uo_out[0]),
    .X(_0321_));
 sky130_fd_sc_hd__o211a_1 _1360_ (.A1(_0624_),
    .A2(_0320_),
    .B1(_0321_),
    .C1(net61),
    .X(_0145_));
 sky130_fd_sc_hd__mux4_1 _1361_ (.A0(\stack[3] ),
    .A1(\stack[2] ),
    .A2(\stack[1] ),
    .A3(\stack[0] ),
    .S0(\fetch_count[0] ),
    .S1(\fetch_count[1] ),
    .X(_0322_));
 sky130_fd_sc_hd__mux4_1 _1362_ (.A0(\stack[7] ),
    .A1(\stack[6] ),
    .A2(\stack[5] ),
    .A3(\stack[4] ),
    .S0(\fetch_count[0] ),
    .S1(\fetch_count[1] ),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _1363_ (.A(\fetch_count[2] ),
    .B(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__o211a_1 _1364_ (.A1(_0343_),
    .A2(_0322_),
    .B1(_0324_),
    .C1(net56),
    .X(_0144_));
 sky130_fd_sc_hd__a211o_1 _1365_ (.A1(net224),
    .A2(_0648_),
    .B1(_0689_),
    .C1(_0325_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_2 _1366_ (.A(eeprom_cs),
    .B(net71),
    .Y(eeprom_sck));
 sky130_fd_sc_hd__inv_2 _1368__4 (.A(clknet_4_13_0_clk),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _1369__5 (.A(clknet_4_13_0_clk),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _1370__6 (.A(clknet_4_13_0_clk),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _1371__7 (.A(clknet_4_13_0_clk),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _1372__8 (.A(clknet_4_12_0_clk),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _1373__9 (.A(clknet_4_13_0_clk),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _1374__10 (.A(clknet_4_13_0_clk),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _1375__11 (.A(clknet_4_14_0_clk),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _1376__12 (.A(clknet_4_13_0_clk),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _1377__13 (.A(clknet_4_15_0_clk),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _1378__14 (.A(clknet_4_15_0_clk),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _1379__15 (.A(clknet_4_15_0_clk),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _1380__16 (.A(clknet_4_14_0_clk),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _1381__17 (.A(clknet_4_14_0_clk),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _1382__18 (.A(clknet_4_14_0_clk),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _1383__19 (.A(clknet_4_14_0_clk),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _1384__20 (.A(clknet_4_14_0_clk),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _1385__21 (.A(clknet_4_14_0_clk),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _1386__22 (.A(clknet_4_14_0_clk),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _1387__23 (.A(clknet_4_12_0_clk),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _1388__24 (.A(clknet_4_7_0_clk),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _1389__25 (.A(clknet_4_3_0_clk),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _1390__26 (.A(clknet_4_5_0_clk),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _1391__27 (.A(clknet_4_4_0_clk),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _1392__28 (.A(clknet_4_5_0_clk),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _1393__29 (.A(clknet_4_5_0_clk),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _1394__30 (.A(clknet_4_5_0_clk),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _1395__31 (.A(clknet_4_5_0_clk),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _1396__32 (.A(clknet_4_5_0_clk),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _1397__33 (.A(clknet_4_5_0_clk),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _1398__34 (.A(clknet_4_5_0_clk),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _1399__35 (.A(clknet_4_4_0_clk),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _1400__36 (.A(clknet_4_4_0_clk),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _1401__37 (.A(clknet_4_5_0_clk),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _1402__38 (.A(clknet_4_7_0_clk),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _1403__39 (.A(clknet_4_7_0_clk),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _1404__40 (.A(clknet_4_7_0_clk),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _1405__41 (.A(clknet_4_7_0_clk),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _1406__42 (.A(clknet_4_4_0_clk),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _1407__43 (.A(clknet_4_4_0_clk),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _1408__44 (.A(clknet_4_4_0_clk),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _1409__45 (.A(clknet_4_4_0_clk),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _1410__46 (.A(clknet_4_1_0_clk),
    .Y(net115));
 sky130_fd_sc_hd__inv_2 _1411__47 (.A(clknet_4_1_0_clk),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _1412__48 (.A(clknet_4_1_0_clk),
    .Y(net117));
 sky130_fd_sc_hd__inv_2 _1413__49 (.A(clknet_4_1_0_clk),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _1414__50 (.A(clknet_4_7_0_clk),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _1415__51 (.A(clknet_4_7_0_clk),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _1416__52 (.A(clknet_4_7_0_clk),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _1417__53 (.A(clknet_4_7_0_clk),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _1418__54 (.A(clknet_4_6_0_clk),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _1419__55 (.A(clknet_4_6_0_clk),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _1420__56 (.A(clknet_4_7_0_clk),
    .Y(net125));
 sky130_fd_sc_hd__inv_2 _1421__57 (.A(clknet_4_6_0_clk),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _1422__58 (.A(clknet_4_4_0_clk),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _1423__59 (.A(clknet_4_4_0_clk),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _1424__60 (.A(clknet_4_6_0_clk),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _1425__61 (.A(clknet_4_1_0_clk),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _1426__62 (.A(clknet_4_3_0_clk),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _1427__63 (.A(clknet_4_1_0_clk),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _1428__64 (.A(clknet_4_1_0_clk),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _1429__65 (.A(clknet_4_3_0_clk),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _1430__66 (.A(clknet_4_12_0_clk),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _1431__67 (.A(clknet_4_11_0_clk),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _1432__68 (.A(clknet_4_11_0_clk),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _1433__69 (.A(clknet_4_12_0_clk),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _1434__70 (.A(clknet_4_6_0_clk),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _1435__71 (.A(clknet_4_6_0_clk),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _1436__72 (.A(clknet_4_6_0_clk),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _1437__73 (.A(clknet_4_6_0_clk),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _1438__74 (.A(clknet_4_12_0_clk),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _1439__75 (.A(clknet_4_2_0_clk),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _1440__76 (.A(clknet_4_2_0_clk),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _1441__77 (.A(clknet_4_2_0_clk),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _1442__78 (.A(clknet_4_2_0_clk),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _1443__79 (.A(clknet_4_0_0_clk),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _1444__80 (.A(clknet_4_0_0_clk),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _1445__81 (.A(clknet_4_0_0_clk),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _1446__82 (.A(clknet_4_0_0_clk),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _1447__83 (.A(clknet_4_0_0_clk),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _1448__84 (.A(clknet_4_0_0_clk),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _1449__85 (.A(clknet_4_0_0_clk),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _1450__86 (.A(clknet_4_0_0_clk),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _1451__87 (.A(clknet_4_0_0_clk),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _1452__88 (.A(clknet_4_0_0_clk),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _1453__89 (.A(clknet_4_0_0_clk),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _1454__90 (.A(clknet_4_0_0_clk),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _1455__91 (.A(clknet_4_10_0_clk),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _1456__92 (.A(clknet_4_10_0_clk),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _1457__93 (.A(clknet_4_10_0_clk),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _1458__94 (.A(clknet_4_10_0_clk),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _1459__95 (.A(clknet_4_10_0_clk),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _1460__96 (.A(clknet_4_10_0_clk),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _1461__97 (.A(clknet_4_10_0_clk),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _1462__98 (.A(clknet_4_10_0_clk),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _1463__99 (.A(clknet_4_10_0_clk),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _1464__100 (.A(clknet_4_8_0_clk),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _1465__101 (.A(clknet_4_8_0_clk),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _1466__102 (.A(clknet_4_8_0_clk),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _1467__103 (.A(clknet_4_8_0_clk),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _1468__104 (.A(clknet_4_8_0_clk),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _1469__105 (.A(clknet_4_2_0_clk),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _1470__106 (.A(clknet_4_2_0_clk),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _1471__107 (.A(clknet_4_1_0_clk),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _1472__108 (.A(clknet_4_1_0_clk),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _1473__109 (.A(clknet_4_0_0_clk),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _1474__110 (.A(clknet_4_1_0_clk),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _1475__111 (.A(clknet_4_11_0_clk),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _1476__112 (.A(clknet_4_11_0_clk),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _1477__113 (.A(clknet_4_9_0_clk),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _1478__114 (.A(clknet_4_11_0_clk),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _1479__115 (.A(clknet_4_11_0_clk),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _1480__116 (.A(clknet_4_10_0_clk),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _1481__117 (.A(clknet_4_9_0_clk),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _1482__118 (.A(clknet_4_9_0_clk),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _1483__119 (.A(clknet_4_2_0_clk),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _1484__120 (.A(clknet_4_2_0_clk),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _1485__121 (.A(clknet_4_2_0_clk),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _1486__122 (.A(clknet_4_3_0_clk),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _1487__123 (.A(clknet_4_3_0_clk),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _1488__124 (.A(clknet_4_2_0_clk),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _1489__125 (.A(clknet_4_3_0_clk),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _1490__126 (.A(clknet_4_3_0_clk),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _1491__127 (.A(clknet_4_12_0_clk),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _1492__128 (.A(clknet_4_2_0_clk),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _1493__129 (.A(clknet_4_9_0_clk),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _1494__130 (.A(clknet_4_11_0_clk),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _1495__131 (.A(clknet_4_11_0_clk),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _1496__132 (.A(clknet_4_11_0_clk),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _1497__133 (.A(clknet_4_11_0_clk),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _1498__134 (.A(clknet_4_11_0_clk),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _1499__135 (.A(clknet_4_9_0_clk),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _1500__136 (.A(clknet_4_9_0_clk),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _1501__137 (.A(clknet_4_3_0_clk),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _1502__138 (.A(clknet_4_3_0_clk),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _1503__139 (.A(clknet_4_8_0_clk),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _1504__140 (.A(clknet_4_9_0_clk),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _1505__141 (.A(clknet_4_9_0_clk),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _1506__142 (.A(clknet_4_9_0_clk),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _1507__143 (.A(clknet_4_3_0_clk),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _1508__144 (.A(clknet_4_3_0_clk),
    .Y(net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _1509_ (.CLK(net70),
    .D(_0143_),
    .Q(eeprom_cs));
 sky130_fd_sc_hd__dfxtp_1 _1510_ (.CLK(net72),
    .D(_0144_),
    .Q(stack_out));
 sky130_fd_sc_hd__dfxtp_4 _1511_ (.CLK(net73),
    .D(_0145_),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_4 _1512_ (.CLK(net74),
    .D(_0146_),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_4 _1513_ (.CLK(net75),
    .D(_0147_),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_2 _1514_ (.CLK(net76),
    .D(_0148_),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_1 _1515_ (.CLK(net77),
    .D(_0149_),
    .Q(timer_mode));
 sky130_fd_sc_hd__dfxtp_1 _1516_ (.CLK(net78),
    .D(_0150_),
    .Q(\stack[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1517_ (.CLK(net79),
    .D(_0151_),
    .Q(\stack[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1518_ (.CLK(net80),
    .D(_0152_),
    .Q(\stack[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1519_ (.CLK(net81),
    .D(_0153_),
    .Q(\stack[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1520_ (.CLK(net82),
    .D(_0154_),
    .Q(\stack[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1521_ (.CLK(net83),
    .D(_0155_),
    .Q(\stack[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1522_ (.CLK(net84),
    .D(_0156_),
    .Q(\stack[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1523_ (.CLK(net85),
    .D(_0157_),
    .Q(\stack[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1524_ (.CLK(net86),
    .D(_0158_),
    .Q(\stack[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1525_ (.CLK(net87),
    .D(_0159_),
    .Q(\stack[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1526_ (.CLK(net88),
    .D(_0160_),
    .Q(\stack[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1527_ (.CLK(net89),
    .D(_0161_),
    .Q(\stack[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1528_ (.CLK(net90),
    .D(_0162_),
    .Q(\stack[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1529_ (.CLK(net91),
    .D(_0163_),
    .Q(\stack[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1530_ (.CLK(net92),
    .D(_0164_),
    .Q(\stack[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1531_ (.CLK(net93),
    .D(_0165_),
    .Q(eeprom_copi));
 sky130_fd_sc_hd__dfxtp_1 _1532_ (.CLK(net94),
    .D(_0166_),
    .Q(timer_out));
 sky130_fd_sc_hd__dfxtp_1 _1533_ (.CLK(clknet_4_13_0_clk),
    .D(net10),
    .Q(\uio_in_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1534_ (.CLK(clknet_4_15_0_clk),
    .D(net2),
    .Q(\ui_in_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1535_ (.CLK(clknet_4_15_0_clk),
    .D(net3),
    .Q(\ui_in_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1536_ (.CLK(clknet_4_15_0_clk),
    .D(net4),
    .Q(\ui_in_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1537_ (.CLK(clknet_4_15_0_clk),
    .D(net5),
    .Q(\ui_in_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1538_ (.CLK(clknet_4_15_0_clk),
    .D(net6),
    .Q(\ui_in_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1539_ (.CLK(clknet_4_15_0_clk),
    .D(net7),
    .Q(\ui_in_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1540_ (.CLK(clknet_4_15_0_clk),
    .D(net8),
    .Q(\ui_in_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1541_ (.CLK(clknet_4_15_0_clk),
    .D(net9),
    .Q(\ui_in_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1542_ (.CLK(net95),
    .D(_0167_),
    .Q(eeprom_oe_copi));
 sky130_fd_sc_hd__dfxtp_2 _1543_ (.CLK(net96),
    .D(_0168_),
    .Q(\fetch_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1544_ (.CLK(net97),
    .D(_0169_),
    .Q(\fetch_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1545_ (.CLK(net98),
    .D(_0170_),
    .Q(\fetch_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1546_ (.CLK(net99),
    .D(_0171_),
    .Q(\fetch_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1547_ (.CLK(net100),
    .D(_0172_),
    .Q(\fetch_count[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1548_ (.CLK(net101),
    .D(_0173_),
    .Q(\fetch_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1549_ (.CLK(net102),
    .D(_0174_),
    .Q(\fetch_count[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1550_ (.CLK(net103),
    .D(_0175_),
    .Q(\fetch_prev_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1551_ (.CLK(net104),
    .D(_0176_),
    .Q(\fetch_prev_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1552_ (.CLK(net105),
    .D(net226),
    .Q(\fetch_prev_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1553_ (.CLK(net106),
    .D(_0178_),
    .Q(\fetch_prev_state[3] ));
 sky130_fd_sc_hd__dfxtp_4 _1554_ (.CLK(net107),
    .D(_0179_),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_4 _1555_ (.CLK(net108),
    .D(_0180_),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_4 _1556_ (.CLK(net109),
    .D(_0181_),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_4 _1557_ (.CLK(net110),
    .D(_0182_),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfxtp_1 _1558_ (.CLK(net111),
    .D(_0183_),
    .Q(\cur_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1559_ (.CLK(net112),
    .D(_0184_),
    .Q(\cur_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1560_ (.CLK(net113),
    .D(_0185_),
    .Q(\cur_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1561_ (.CLK(net114),
    .D(_0186_),
    .Q(\cur_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1562_ (.CLK(net115),
    .D(_0187_),
    .Q(\cur_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1563_ (.CLK(net116),
    .D(_0188_),
    .Q(\cur_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1564_ (.CLK(net117),
    .D(_0189_),
    .Q(\cur_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1565_ (.CLK(net118),
    .D(net223),
    .Q(\cur_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1566_ (.CLK(net119),
    .D(_0191_),
    .Q(\cycle_start_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1567_ (.CLK(net120),
    .D(_0192_),
    .Q(\cycle_start_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1568_ (.CLK(net121),
    .D(_0193_),
    .Q(\cycle_start_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1569_ (.CLK(net122),
    .D(_0194_),
    .Q(\cycle_start_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1570_ (.CLK(net123),
    .D(_0195_),
    .Q(\cycle_start_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1571_ (.CLK(net124),
    .D(_0196_),
    .Q(\cycle_start_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1572_ (.CLK(net125),
    .D(_0197_),
    .Q(\cycle_start_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1573_ (.CLK(net126),
    .D(_0198_),
    .Q(\cycle_start_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1574_ (.CLK(net127),
    .D(_0199_),
    .Q(\cycle_end_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1575_ (.CLK(net128),
    .D(_0200_),
    .Q(\cycle_end_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1576_ (.CLK(net129),
    .D(_0201_),
    .Q(\cycle_end_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1577_ (.CLK(net130),
    .D(_0202_),
    .Q(\cycle_end_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1578_ (.CLK(net131),
    .D(_0203_),
    .Q(\cycle_end_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1579_ (.CLK(net132),
    .D(_0204_),
    .Q(\cycle_end_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1580_ (.CLK(net133),
    .D(_0205_),
    .Q(\cycle_end_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1581_ (.CLK(net134),
    .D(_0206_),
    .Q(\cycle_end_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1582_ (.CLK(net135),
    .D(_0207_),
    .Q(\instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1583_ (.CLK(net136),
    .D(_0208_),
    .Q(\instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1584_ (.CLK(net137),
    .D(_0209_),
    .Q(\instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1585_ (.CLK(net138),
    .D(_0210_),
    .Q(\instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1586_ (.CLK(net139),
    .D(_0211_),
    .Q(\instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1587_ (.CLK(net140),
    .D(_0212_),
    .Q(\instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1588_ (.CLK(net141),
    .D(_0213_),
    .Q(\instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1589_ (.CLK(net142),
    .D(_0214_),
    .Q(\instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1590_ (.CLK(net143),
    .D(_0215_),
    .Q(\stack[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1591_ (.CLK(net144),
    .D(_0216_),
    .Q(\timer_clock_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1592_ (.CLK(net145),
    .D(net243),
    .Q(\timer_clock_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1593_ (.CLK(net146),
    .D(_0218_),
    .Q(\timer_clock_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1594_ (.CLK(net147),
    .D(_0219_),
    .Q(\timer_clock_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1595_ (.CLK(net148),
    .D(_0220_),
    .Q(\timer_clock_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1596_ (.CLK(net149),
    .D(_0221_),
    .Q(\timer_clock_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1597_ (.CLK(net150),
    .D(_0222_),
    .Q(\timer_clock_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1598_ (.CLK(net151),
    .D(_0223_),
    .Q(\timer_clock_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1599_ (.CLK(net152),
    .D(_0224_),
    .Q(\timer_clock_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1600_ (.CLK(net153),
    .D(_0225_),
    .Q(\timer_clock_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1601_ (.CLK(net154),
    .D(_0226_),
    .Q(\timer_clock_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1602_ (.CLK(net155),
    .D(_0227_),
    .Q(\timer_clock_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1603_ (.CLK(net156),
    .D(_0228_),
    .Q(\timer_clock_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1604_ (.CLK(net157),
    .D(_0229_),
    .Q(\timer_clock_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1605_ (.CLK(net158),
    .D(_0230_),
    .Q(\timer_clock_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1606_ (.CLK(net159),
    .D(_0231_),
    .Q(\timer_clock_counter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1607_ (.CLK(net160),
    .D(_0232_),
    .Q(\timer_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1608_ (.CLK(net161),
    .D(_0233_),
    .Q(\timer_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1609_ (.CLK(net162),
    .D(_0234_),
    .Q(\timer_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1610_ (.CLK(net163),
    .D(_0235_),
    .Q(\timer_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1611_ (.CLK(net164),
    .D(_0236_),
    .Q(\timer_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1612_ (.CLK(net165),
    .D(_0237_),
    .Q(\timer_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1613_ (.CLK(net166),
    .D(_0238_),
    .Q(\timer_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1614_ (.CLK(net167),
    .D(_0239_),
    .Q(\timer_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1615_ (.CLK(net168),
    .D(_0240_),
    .Q(\timer_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1616_ (.CLK(net169),
    .D(_0241_),
    .Q(\timer_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1617_ (.CLK(net170),
    .D(_0242_),
    .Q(\timer_counter[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1618_ (.CLK(net171),
    .D(_0243_),
    .Q(\timer_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1619_ (.CLK(net172),
    .D(_0244_),
    .Q(\timer_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1620_ (.CLK(net173),
    .D(_0245_),
    .Q(\timer_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1621_ (.CLK(net174),
    .D(_0246_),
    .Q(\timer_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1622_ (.CLK(net175),
    .D(_0247_),
    .Q(\timer_counter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1623_ (.CLK(net176),
    .D(_0248_),
    .Q(\timer_clock_divisor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1624_ (.CLK(net177),
    .D(_0249_),
    .Q(\timer_clock_divisor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1625_ (.CLK(net178),
    .D(_0250_),
    .Q(\timer_clock_divisor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1626_ (.CLK(net179),
    .D(_0251_),
    .Q(\timer_clock_divisor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1627_ (.CLK(net180),
    .D(_0252_),
    .Q(\timer_period_a[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1628_ (.CLK(net181),
    .D(_0253_),
    .Q(\timer_period_a[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1629_ (.CLK(net182),
    .D(_0254_),
    .Q(\timer_period_a[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1630_ (.CLK(net183),
    .D(_0255_),
    .Q(\timer_period_a[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1631_ (.CLK(net184),
    .D(_0256_),
    .Q(\timer_period_a[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1632_ (.CLK(net185),
    .D(_0257_),
    .Q(\timer_period_a[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1633_ (.CLK(net186),
    .D(_0258_),
    .Q(\timer_period_a[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1634_ (.CLK(net187),
    .D(_0259_),
    .Q(\timer_period_a[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1635_ (.CLK(net188),
    .D(_0260_),
    .Q(\timer_period_a[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1636_ (.CLK(net189),
    .D(_0261_),
    .Q(\timer_period_a[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1637_ (.CLK(net190),
    .D(_0262_),
    .Q(\timer_period_a[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1638_ (.CLK(net191),
    .D(_0263_),
    .Q(\timer_period_a[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1639_ (.CLK(net192),
    .D(_0264_),
    .Q(\timer_period_a[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1640_ (.CLK(net193),
    .D(_0265_),
    .Q(\timer_period_a[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1641_ (.CLK(net194),
    .D(_0266_),
    .Q(\timer_period_a[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1642_ (.CLK(net195),
    .D(_0267_),
    .Q(\timer_period_a[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1643_ (.CLK(net196),
    .D(_0268_),
    .Q(timer_enabled));
 sky130_fd_sc_hd__dfxtp_1 _1644_ (.CLK(net197),
    .D(_0269_),
    .Q(timer_phase));
 sky130_fd_sc_hd__dfxtp_1 _1645_ (.CLK(net198),
    .D(_0270_),
    .Q(\timer_period_b[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1646_ (.CLK(net199),
    .D(_0271_),
    .Q(\timer_period_b[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1647_ (.CLK(net200),
    .D(_0272_),
    .Q(\timer_period_b[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1648_ (.CLK(net201),
    .D(_0273_),
    .Q(\timer_period_b[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1649_ (.CLK(net202),
    .D(_0274_),
    .Q(\timer_period_b[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1650_ (.CLK(net203),
    .D(_0275_),
    .Q(\timer_period_b[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1651_ (.CLK(net204),
    .D(_0276_),
    .Q(\timer_period_b[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1652_ (.CLK(net205),
    .D(_0277_),
    .Q(\timer_period_b[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1653_ (.CLK(net206),
    .D(_0278_),
    .Q(\timer_period_b[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1654_ (.CLK(net207),
    .D(_0279_),
    .Q(\timer_period_b[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1655_ (.CLK(net208),
    .D(_0280_),
    .Q(\timer_period_b[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1656_ (.CLK(net209),
    .D(_0281_),
    .Q(\timer_period_b[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1657_ (.CLK(net210),
    .D(_0282_),
    .Q(\timer_period_b[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1658_ (.CLK(net211),
    .D(_0283_),
    .Q(\timer_period_b[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1659_ (.CLK(net212),
    .D(_0284_),
    .Q(\timer_period_b[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1660_ (.CLK(net213),
    .D(_0285_),
    .Q(\timer_period_b[15] ));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_69 (.LO(net69));
 sky130_fd_sc_hd__inv_2 _0781__1 (.A(clknet_4_5_0_clk),
    .Y(net70));
 sky130_fd_sc_hd__buf_2 _1667_ (.A(eeprom_oe_copi),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__buf_2 _1668_ (.A(eeprom_oe_copi),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__buf_2 _1669_ (.A(eeprom_oe_copi),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__buf_2 _1670_ (.A(eeprom_oe_copi),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__buf_2 _1671_ (.A(eeprom_oe_copi),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__buf_2 _1672_ (.A(eeprom_sck),
    .X(uio_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _1673_ (.A(eeprom_cs),
    .X(uio_out[1]));
 sky130_fd_sc_hd__clkbuf_4 _1674_ (.A(eeprom_copi),
    .X(uio_out[2]));
 sky130_fd_sc_hd__clkbuf_4 _1675_ (.A(stack_out),
    .X(uio_out[6]));
 sky130_fd_sc_hd__clkbuf_4 _1676_ (.A(timer_out),
    .X(uio_out[7]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 fanout11 (.A(_0516_),
    .X(net11));
 sky130_fd_sc_hd__buf_1 fanout12 (.A(_0516_),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(_0724_),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(_0723_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout16 (.A(_0546_),
    .X(net16));
 sky130_fd_sc_hd__buf_1 wire17 (.A(_0498_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 wire18 (.A(_0395_),
    .X(net18));
 sky130_fd_sc_hd__buf_2 wire19 (.A(_0418_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(_0570_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(_0459_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(_0626_),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(_0625_),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(_0466_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 fanout28 (.A(_0465_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(timer_enabled),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(timer_enabled),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(timer_enabled),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(\instr[7] ),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(\instr[6] ),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(\instr[5] ),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(\instr[4] ),
    .X(net39));
 sky130_fd_sc_hd__buf_1 fanout40 (.A(\instr[4] ),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(\instr[3] ),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(\instr[2] ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(\instr[1] ),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(\instr[0] ),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(\fetch_state[1] ),
    .X(net50));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net63),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net63),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(net63),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net57),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net57),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net63),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(net62),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(net62),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net62),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(net1),
    .X(net63));
 sky130_fd_sc_hd__conb_1 tt_um_jimktrains_vslc_64 (.LO(net64));
 sky130_fd_sc_hd__inv_2 _0781__2 (.A(clknet_4_5_0_clk),
    .Y(net71));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__inv_4 clkload1 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_4 clkload2 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__inv_8 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__inv_4 clkload4 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_4 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__inv_16 clkload7 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__inv_8 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__inv_4 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_16 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_12 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__inv_16 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\timer_clock_counter[15] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\fetch_state[1] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\fetch_prev_state[3] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\timer_clock_counter[13] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\timer_clock_counter[10] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\timer_period_a[4] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\timer_clock_counter[6] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(eeprom_copi),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\cur_addr[7] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0190_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(eeprom_cs),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\fetch_prev_state[2] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0177_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\timer_clock_counter[8] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\timer_clock_counter[4] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(timer_mode),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(eeprom_oe_copi),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\cur_addr[3] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\cur_addr[2] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\timer_period_b[12] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\cur_addr[5] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0610_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\timer_period_b[4] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\timer_counter[13] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\timer_clock_counter[12] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\instr[1] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\cur_addr[6] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\timer_clock_counter[7] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\timer_clock_counter[0] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0217_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\timer_clock_counter[9] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\stack[14] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\cur_addr[1] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\cur_addr[4] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\cycle_end_addr[0] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(timer_phase),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\timer_counter[10] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\fetch_count[2] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\stack[13] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\stack[9] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\stack[11] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\fetch_state[0] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\cycle_start_addr[6] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\stack[12] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\cycle_start_addr[0] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\stack[8] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\cycle_start_addr[7] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\timer_counter[11] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\cycle_start_addr[4] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\cycle_start_addr[5] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\cycle_start_addr[3] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\stack[10] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\cycle_end_addr[1] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\fetch_state[2] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\fetch_prev_state[1] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\cycle_start_addr[1] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\cycle_start_addr[2] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\cur_addr[1] ),
    .X(net271));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 assign uio_oe[3] = net64;
 assign uio_oe[4] = net65;
 assign uio_oe[5] = net66;
 assign uio_out[3] = net67;
 assign uio_out[4] = net68;
 assign uio_out[5] = net69;
endmodule
