magic
tech sky130A
magscale 1 2
timestamp 1738303524
<< viali >>
rect 6101 21641 6135 21675
rect 8033 21641 8067 21675
rect 8401 21641 8435 21675
rect 8677 21641 8711 21675
rect 11713 21641 11747 21675
rect 12265 21641 12299 21675
rect 13001 21641 13035 21675
rect 18061 21641 18095 21675
rect 27905 21641 27939 21675
rect 7849 21505 7883 21539
rect 14105 21505 14139 21539
rect 24685 21505 24719 21539
rect 2237 21437 2271 21471
rect 2789 21437 2823 21471
rect 2973 21437 3007 21471
rect 5181 21437 5215 21471
rect 5457 21437 5491 21471
rect 6285 21437 6319 21471
rect 6469 21437 6503 21471
rect 6745 21437 6779 21471
rect 12909 21437 12943 21471
rect 17141 21437 17175 21471
rect 21557 21437 21591 21471
rect 22109 21437 22143 21471
rect 22201 21437 22235 21471
rect 23857 21437 23891 21471
rect 24409 21437 24443 21471
rect 26433 21437 26467 21471
rect 26709 21437 26743 21471
rect 27169 21437 27203 21471
rect 27721 21437 27755 21471
rect 28273 21437 28307 21471
rect 29009 21437 29043 21471
rect 5549 21369 5583 21403
rect 7021 21369 7055 21403
rect 7205 21369 7239 21403
rect 7297 21369 7331 21403
rect 13921 21369 13955 21403
rect 17877 21369 17911 21403
rect 18077 21369 18111 21403
rect 24952 21369 24986 21403
rect 29254 21369 29288 21403
rect 2145 21301 2179 21335
rect 2881 21301 2915 21335
rect 5273 21301 5307 21335
rect 6653 21301 6687 21335
rect 6837 21301 6871 21335
rect 12817 21301 12851 21335
rect 13553 21301 13587 21335
rect 14013 21301 14047 21335
rect 17049 21301 17083 21335
rect 18245 21301 18279 21335
rect 21465 21301 21499 21335
rect 21925 21301 21959 21335
rect 22385 21301 22419 21335
rect 24041 21301 24075 21335
rect 24593 21301 24627 21335
rect 26065 21301 26099 21335
rect 26617 21301 26651 21335
rect 26893 21301 26927 21335
rect 27353 21301 27387 21335
rect 28457 21301 28491 21335
rect 30389 21301 30423 21335
rect 3525 21097 3559 21131
rect 7205 21097 7239 21131
rect 8585 21097 8619 21131
rect 8953 21097 8987 21131
rect 9781 21097 9815 21131
rect 14749 21097 14783 21131
rect 18797 21097 18831 21131
rect 22661 21097 22695 21131
rect 25145 21097 25179 21131
rect 30139 21097 30173 21131
rect 6092 21029 6126 21063
rect 23940 21029 23974 21063
rect 28702 21029 28736 21063
rect 29929 21029 29963 21063
rect 1961 20961 1995 20995
rect 2228 20961 2262 20995
rect 3709 20961 3743 20995
rect 3893 20961 3927 20995
rect 4169 20961 4203 20995
rect 4721 20961 4755 20995
rect 4905 20961 4939 20995
rect 5825 20961 5859 20995
rect 7573 20961 7607 20995
rect 8033 20961 8067 20995
rect 8401 20961 8435 20995
rect 8769 20961 8803 20995
rect 9321 20961 9355 20995
rect 9505 20961 9539 20995
rect 9597 20961 9631 20995
rect 10425 20961 10459 20995
rect 11253 20961 11287 20995
rect 12633 20961 12667 20995
rect 16865 20961 16899 20995
rect 17132 20961 17166 20995
rect 18889 20961 18923 20995
rect 19436 20961 19470 20995
rect 19533 20961 19567 20995
rect 19625 20961 19659 20995
rect 19753 20961 19787 20995
rect 19901 20961 19935 20995
rect 20913 20961 20947 20995
rect 21281 20961 21315 20995
rect 25329 20961 25363 20995
rect 25513 20961 25547 20995
rect 27241 20961 27275 20995
rect 28457 20961 28491 20995
rect 9137 20893 9171 20927
rect 12909 20893 12943 20927
rect 14841 20893 14875 20927
rect 14933 20893 14967 20927
rect 18981 20893 19015 20927
rect 21557 20893 21591 20927
rect 23673 20893 23707 20927
rect 26985 20893 27019 20927
rect 4077 20825 4111 20859
rect 14381 20825 14415 20859
rect 18429 20825 18463 20859
rect 30297 20825 30331 20859
rect 3341 20757 3375 20791
rect 4813 20757 4847 20791
rect 7849 20757 7883 20791
rect 8217 20757 8251 20791
rect 10333 20757 10367 20791
rect 11529 20757 11563 20791
rect 14197 20757 14231 20791
rect 18245 20757 18279 20791
rect 19257 20757 19291 20791
rect 21005 20757 21039 20791
rect 25053 20757 25087 20791
rect 25697 20757 25731 20791
rect 28365 20757 28399 20791
rect 29837 20757 29871 20791
rect 30113 20757 30147 20791
rect 4813 20553 4847 20587
rect 7021 20553 7055 20587
rect 9597 20553 9631 20587
rect 13553 20553 13587 20587
rect 15025 20553 15059 20587
rect 17141 20553 17175 20587
rect 17969 20553 18003 20587
rect 18061 20553 18095 20587
rect 18889 20553 18923 20587
rect 21097 20553 21131 20587
rect 4629 20485 4663 20519
rect 9321 20485 9355 20519
rect 13369 20485 13403 20519
rect 18705 20485 18739 20519
rect 3249 20417 3283 20451
rect 5365 20417 5399 20451
rect 7665 20417 7699 20451
rect 12173 20417 12207 20451
rect 12817 20417 12851 20451
rect 14105 20417 14139 20451
rect 14381 20417 14415 20451
rect 14565 20417 14599 20451
rect 15209 20417 15243 20451
rect 15393 20417 15427 20451
rect 15853 20417 15887 20451
rect 16129 20417 16163 20451
rect 16246 20417 16280 20451
rect 17969 20417 18003 20451
rect 22569 20417 22603 20451
rect 24409 20417 24443 20451
rect 1317 20349 1351 20383
rect 1409 20349 1443 20383
rect 1593 20349 1627 20383
rect 5641 20349 5675 20383
rect 8125 20349 8159 20383
rect 8677 20349 8711 20383
rect 10977 20349 11011 20383
rect 11161 20349 11195 20383
rect 11253 20349 11287 20383
rect 11897 20349 11931 20383
rect 12357 20349 12391 20383
rect 13737 20349 13771 20383
rect 13921 20349 13955 20383
rect 14013 20349 14047 20383
rect 14197 20349 14231 20383
rect 16405 20349 16439 20383
rect 17325 20349 17359 20383
rect 17509 20349 17543 20383
rect 18153 20349 18187 20383
rect 20453 20349 20487 20383
rect 20637 20349 20671 20383
rect 20729 20349 20763 20383
rect 20821 20349 20855 20383
rect 21189 20349 21223 20383
rect 21465 20349 21499 20383
rect 23121 20349 23155 20383
rect 23397 20349 23431 20383
rect 24676 20349 24710 20383
rect 25881 20349 25915 20383
rect 26137 20349 26171 20383
rect 29009 20349 29043 20383
rect 29276 20349 29310 20383
rect 1860 20281 1894 20315
rect 3494 20281 3528 20315
rect 5908 20281 5942 20315
rect 8953 20281 8987 20315
rect 10710 20281 10744 20315
rect 12909 20281 12943 20315
rect 17049 20281 17083 20315
rect 17785 20281 17819 20315
rect 19073 20281 19107 20315
rect 2973 20213 3007 20247
rect 7113 20213 7147 20247
rect 7941 20213 7975 20247
rect 8769 20213 8803 20247
rect 9413 20213 9447 20247
rect 11989 20213 12023 20247
rect 12541 20213 12575 20247
rect 13001 20213 13035 20247
rect 14657 20213 14691 20247
rect 18873 20213 18907 20247
rect 22937 20213 22971 20247
rect 23305 20213 23339 20247
rect 25789 20213 25823 20247
rect 27261 20213 27295 20247
rect 30389 20213 30423 20247
rect 2329 20009 2363 20043
rect 2697 20009 2731 20043
rect 2973 20009 3007 20043
rect 5457 20009 5491 20043
rect 5825 20009 5859 20043
rect 6561 20009 6595 20043
rect 10977 20009 11011 20043
rect 13829 20009 13863 20043
rect 14565 20009 14599 20043
rect 19073 20009 19107 20043
rect 20913 20009 20947 20043
rect 21281 20009 21315 20043
rect 22017 20009 22051 20043
rect 22385 20009 22419 20043
rect 26433 20009 26467 20043
rect 28089 20009 28123 20043
rect 14473 19941 14507 19975
rect 19441 19941 19475 19975
rect 26709 19941 26743 19975
rect 29101 19941 29135 19975
rect 30113 19941 30147 19975
rect 2053 19873 2087 19907
rect 2237 19873 2271 19907
rect 2513 19873 2547 19907
rect 2789 19873 2823 19907
rect 3065 19873 3099 19907
rect 3341 19873 3375 19907
rect 3893 19873 3927 19907
rect 3985 19873 4019 19907
rect 4905 19873 4939 19907
rect 5365 19873 5399 19907
rect 6009 19873 6043 19907
rect 6101 19873 6135 19907
rect 6285 19873 6319 19907
rect 6377 19873 6411 19907
rect 6653 19873 6687 19907
rect 9137 19873 9171 19907
rect 9404 19873 9438 19907
rect 12265 19873 12299 19907
rect 12541 19873 12575 19907
rect 14933 19873 14967 19907
rect 15117 19873 15151 19907
rect 15485 19873 15519 19907
rect 15853 19873 15887 19907
rect 16129 19873 16163 19907
rect 16221 19873 16255 19907
rect 16405 19873 16439 19907
rect 16681 19873 16715 19907
rect 16865 19873 16899 19907
rect 18705 19873 18739 19907
rect 18889 19873 18923 19907
rect 18981 19873 19015 19907
rect 19257 19873 19291 19907
rect 19533 19873 19567 19907
rect 19625 19873 19659 19907
rect 20913 19873 20947 19907
rect 21097 19873 21131 19907
rect 21557 19873 21591 19907
rect 21649 19873 21683 19907
rect 21741 19873 21775 19907
rect 21925 19873 21959 19907
rect 22201 19873 22235 19907
rect 22477 19873 22511 19907
rect 24869 19873 24903 19907
rect 24961 19873 24995 19907
rect 25145 19873 25179 19907
rect 25237 19873 25271 19907
rect 25329 19873 25363 19907
rect 25789 19873 25823 19907
rect 25881 19873 25915 19907
rect 26065 19873 26099 19907
rect 26157 19873 26191 19907
rect 26617 19873 26651 19907
rect 26801 19873 26835 19907
rect 26985 19873 27019 19907
rect 27813 19873 27847 19907
rect 28181 19873 28215 19907
rect 28963 19873 28997 19907
rect 29193 19873 29227 19907
rect 29376 19873 29410 19907
rect 29469 19873 29503 19907
rect 29745 19873 29779 19907
rect 29929 19873 29963 19907
rect 2973 19805 3007 19839
rect 11529 19805 11563 19839
rect 14749 19805 14783 19839
rect 15025 19805 15059 19839
rect 10517 19737 10551 19771
rect 15301 19737 15335 19771
rect 25513 19737 25547 19771
rect 2145 19669 2179 19703
rect 3249 19669 3283 19703
rect 3617 19669 3651 19703
rect 3985 19669 4019 19703
rect 4813 19669 4847 19703
rect 14105 19669 14139 19703
rect 15761 19669 15795 19703
rect 16589 19669 16623 19703
rect 16773 19669 16807 19703
rect 18521 19669 18555 19703
rect 19717 19669 19751 19703
rect 25605 19669 25639 19703
rect 27445 19669 27479 19703
rect 27721 19669 27755 19703
rect 27905 19669 27939 19703
rect 28825 19669 28859 19703
rect 29653 19669 29687 19703
rect 4629 19465 4663 19499
rect 9965 19465 9999 19499
rect 16313 19465 16347 19499
rect 18797 19465 18831 19499
rect 21465 19465 21499 19499
rect 25881 19465 25915 19499
rect 27997 19465 28031 19499
rect 4353 19397 4387 19431
rect 7849 19397 7883 19431
rect 28089 19397 28123 19431
rect 8493 19329 8527 19363
rect 9413 19329 9447 19363
rect 9505 19329 9539 19363
rect 14197 19329 14231 19363
rect 14381 19329 14415 19363
rect 16773 19329 16807 19363
rect 20361 19329 20395 19363
rect 1869 19261 1903 19295
rect 2697 19261 2731 19295
rect 2881 19261 2915 19295
rect 2973 19261 3007 19295
rect 3249 19261 3283 19295
rect 4451 19261 4485 19295
rect 4629 19261 4663 19295
rect 7665 19261 7699 19295
rect 8401 19261 8435 19295
rect 8585 19261 8619 19295
rect 9045 19261 9079 19295
rect 9137 19261 9171 19295
rect 9321 19261 9355 19295
rect 9689 19261 9723 19295
rect 9873 19261 9907 19295
rect 10241 19261 10275 19295
rect 10333 19261 10367 19295
rect 10425 19261 10459 19295
rect 10609 19261 10643 19295
rect 10701 19263 10735 19297
rect 14749 19261 14783 19295
rect 15025 19261 15059 19295
rect 16497 19261 16531 19295
rect 16681 19261 16715 19295
rect 16865 19261 16899 19295
rect 17049 19261 17083 19295
rect 17877 19261 17911 19295
rect 18061 19261 18095 19295
rect 18153 19261 18187 19295
rect 18245 19261 18279 19295
rect 20085 19261 20119 19295
rect 21373 19261 21407 19295
rect 21557 19261 21591 19295
rect 24225 19261 24259 19295
rect 26709 19261 26743 19295
rect 28641 19261 28675 19295
rect 29009 19261 29043 19295
rect 29285 19261 29319 19295
rect 2513 19193 2547 19227
rect 3985 19193 4019 19227
rect 4169 19193 4203 19227
rect 7757 19193 7791 19227
rect 7941 19193 7975 19227
rect 8861 19193 8895 19227
rect 10793 19193 10827 19227
rect 14105 19193 14139 19227
rect 17233 19193 17267 19227
rect 18521 19193 18555 19227
rect 26065 19193 26099 19227
rect 28457 19193 28491 19227
rect 28733 19193 28767 19227
rect 29552 19193 29586 19227
rect 1777 19125 1811 19159
rect 3893 19125 3927 19159
rect 8677 19125 8711 19159
rect 13737 19125 13771 19159
rect 24317 19125 24351 19159
rect 25697 19125 25731 19159
rect 25865 19125 25899 19159
rect 26617 19125 26651 19159
rect 29101 19125 29135 19159
rect 30665 19125 30699 19159
rect 2973 18921 3007 18955
rect 5825 18921 5859 18955
rect 8677 18921 8711 18955
rect 14933 18921 14967 18955
rect 16773 18921 16807 18955
rect 18705 18921 18739 18955
rect 29285 18921 29319 18955
rect 1860 18853 1894 18887
rect 3065 18853 3099 18887
rect 9413 18853 9447 18887
rect 10977 18853 11011 18887
rect 11345 18853 11379 18887
rect 11437 18853 11471 18887
rect 22394 18853 22428 18887
rect 1593 18785 1627 18819
rect 3341 18785 3375 18819
rect 3433 18785 3467 18819
rect 3525 18785 3559 18819
rect 3709 18785 3743 18819
rect 5365 18785 5399 18819
rect 5549 18785 5583 18819
rect 6101 18785 6135 18819
rect 8861 18785 8895 18819
rect 9137 18785 9171 18819
rect 9321 18785 9355 18819
rect 10149 18785 10183 18819
rect 10517 18785 10551 18819
rect 11161 18785 11195 18819
rect 11621 18785 11655 18819
rect 12127 18785 12161 18819
rect 12265 18785 12299 18819
rect 12357 18785 12391 18819
rect 12541 18785 12575 18819
rect 12817 18785 12851 18819
rect 14841 18785 14875 18819
rect 15577 18785 15611 18819
rect 16129 18785 16163 18819
rect 16313 18785 16347 18819
rect 16405 18785 16439 18819
rect 16497 18785 16531 18819
rect 18705 18785 18739 18819
rect 18889 18785 18923 18819
rect 19533 18785 19567 18819
rect 25697 18785 25731 18819
rect 26433 18785 26467 18819
rect 26689 18785 26723 18819
rect 28641 18785 28675 18819
rect 28825 18785 28859 18819
rect 28917 18785 28951 18819
rect 29009 18785 29043 18819
rect 29377 18785 29411 18819
rect 29644 18785 29678 18819
rect 30849 18785 30883 18819
rect 4537 18717 4571 18751
rect 4721 18717 4755 18751
rect 4813 18717 4847 18751
rect 4905 18717 4939 18751
rect 4997 18717 5031 18751
rect 5825 18717 5859 18751
rect 8953 18717 8987 18751
rect 9597 18717 9631 18751
rect 9689 18717 9723 18751
rect 10057 18717 10091 18751
rect 15853 18717 15887 18751
rect 22661 18717 22695 18751
rect 24041 18717 24075 18751
rect 24685 18717 24719 18751
rect 24844 18717 24878 18751
rect 24961 18717 24995 18751
rect 25881 18717 25915 18751
rect 9045 18649 9079 18683
rect 11805 18649 11839 18683
rect 15761 18649 15795 18683
rect 25237 18649 25271 18683
rect 5181 18581 5215 18615
rect 6009 18581 6043 18615
rect 10241 18581 10275 18615
rect 10701 18581 10735 18615
rect 11897 18581 11931 18615
rect 12725 18581 12759 18615
rect 15669 18581 15703 18615
rect 19257 18581 19291 18615
rect 21281 18581 21315 18615
rect 27813 18581 27847 18615
rect 30757 18581 30791 18615
rect 31033 18581 31067 18615
rect 4813 18377 4847 18411
rect 5181 18377 5215 18411
rect 6561 18377 6595 18411
rect 20637 18377 20671 18411
rect 26249 18377 26283 18411
rect 28825 18377 28859 18411
rect 29837 18377 29871 18411
rect 29009 18309 29043 18343
rect 4261 18241 4295 18275
rect 5181 18241 5215 18275
rect 5641 18241 5675 18275
rect 5733 18241 5767 18275
rect 5917 18241 5951 18275
rect 6101 18241 6135 18275
rect 10057 18241 10091 18275
rect 11805 18241 11839 18275
rect 15669 18241 15703 18275
rect 16129 18241 16163 18275
rect 16405 18241 16439 18275
rect 16589 18241 16623 18275
rect 29469 18241 29503 18275
rect 29561 18241 29595 18275
rect 2881 18173 2915 18207
rect 3525 18173 3559 18207
rect 3985 18173 4019 18207
rect 4537 18173 4571 18207
rect 4721 18173 4755 18207
rect 4997 18173 5031 18207
rect 6009 18173 6043 18207
rect 6315 18173 6349 18207
rect 6469 18173 6503 18207
rect 6561 18173 6595 18207
rect 6745 18173 6779 18207
rect 8493 18173 8527 18207
rect 9413 18173 9447 18207
rect 10609 18173 10643 18207
rect 10701 18173 10735 18207
rect 10793 18173 10827 18207
rect 10977 18173 11011 18207
rect 11069 18173 11103 18207
rect 11437 18173 11471 18207
rect 12357 18173 12391 18207
rect 12909 18173 12943 18207
rect 13001 18173 13035 18207
rect 13093 18173 13127 18207
rect 13277 18173 13311 18207
rect 13553 18173 13587 18207
rect 15577 18173 15611 18207
rect 15761 18173 15795 18207
rect 15853 18173 15887 18207
rect 16037 18173 16071 18207
rect 16313 18173 16347 18207
rect 16497 18173 16531 18207
rect 18797 18173 18831 18207
rect 18981 18173 19015 18207
rect 19257 18173 19291 18207
rect 21281 18173 21315 18207
rect 22293 18173 22327 18207
rect 22477 18173 22511 18207
rect 22569 18173 22603 18207
rect 22661 18173 22695 18207
rect 23489 18173 23523 18207
rect 23581 18173 23615 18207
rect 23857 18173 23891 18207
rect 25513 18173 25547 18207
rect 25697 18173 25731 18207
rect 25789 18173 25823 18207
rect 25881 18173 25915 18207
rect 26525 18173 26559 18207
rect 26617 18173 26651 18207
rect 26709 18173 26743 18207
rect 26893 18173 26927 18207
rect 27997 18173 28031 18207
rect 28273 18173 28307 18207
rect 28365 18173 28399 18207
rect 28549 18173 28583 18207
rect 28641 18173 28675 18207
rect 30113 18173 30147 18207
rect 30205 18173 30239 18207
rect 30297 18173 30331 18207
rect 30481 18173 30515 18207
rect 3341 18105 3375 18139
rect 5457 18105 5491 18139
rect 9873 18105 9907 18139
rect 15025 18105 15059 18139
rect 15209 18105 15243 18139
rect 17141 18105 17175 18139
rect 19524 18105 19558 18139
rect 24124 18105 24158 18139
rect 27813 18105 27847 18139
rect 29377 18105 29411 18139
rect 2973 18037 3007 18071
rect 4721 18037 4755 18071
rect 5549 18037 5583 18071
rect 8585 18037 8619 18071
rect 8769 18037 8803 18071
rect 9505 18037 9539 18071
rect 9965 18037 9999 18071
rect 10333 18037 10367 18071
rect 12633 18037 12667 18071
rect 14197 18037 14231 18071
rect 15393 18037 15427 18071
rect 17049 18037 17083 18071
rect 18981 18037 19015 18071
rect 22937 18037 22971 18071
rect 25237 18037 25271 18071
rect 26157 18037 26191 18071
rect 28181 18037 28215 18071
rect 3985 17833 4019 17867
rect 5641 17833 5675 17867
rect 6929 17833 6963 17867
rect 8217 17833 8251 17867
rect 10057 17833 10091 17867
rect 10793 17833 10827 17867
rect 11437 17833 11471 17867
rect 13829 17833 13863 17867
rect 14197 17833 14231 17867
rect 16129 17833 16163 17867
rect 17049 17833 17083 17867
rect 19717 17833 19751 17867
rect 21097 17833 21131 17867
rect 24041 17833 24075 17867
rect 25237 17833 25271 17867
rect 25605 17833 25639 17867
rect 27445 17833 27479 17867
rect 29009 17833 29043 17867
rect 29561 17833 29595 17867
rect 29653 17833 29687 17867
rect 6561 17765 6595 17799
rect 8401 17765 8435 17799
rect 13645 17765 13679 17799
rect 19533 17765 19567 17799
rect 21373 17765 21407 17799
rect 22569 17765 22603 17799
rect 26433 17765 26467 17799
rect 27261 17765 27295 17799
rect 2697 17697 2731 17731
rect 2789 17697 2823 17731
rect 2881 17697 2915 17731
rect 3065 17697 3099 17731
rect 3709 17697 3743 17731
rect 3893 17697 3927 17731
rect 4353 17697 4387 17731
rect 4813 17697 4847 17731
rect 4905 17697 4939 17731
rect 5089 17697 5123 17731
rect 5181 17697 5215 17731
rect 5273 17697 5307 17731
rect 5457 17697 5491 17731
rect 6009 17697 6043 17731
rect 6101 17697 6135 17731
rect 6193 17697 6227 17731
rect 6331 17697 6365 17731
rect 6745 17697 6779 17731
rect 7021 17697 7055 17731
rect 7205 17697 7239 17731
rect 8585 17697 8619 17731
rect 8677 17697 8711 17731
rect 8944 17697 8978 17731
rect 11345 17697 11379 17731
rect 11989 17697 12023 17731
rect 12245 17697 12279 17731
rect 13461 17697 13495 17731
rect 14381 17697 14415 17731
rect 14473 17697 14507 17731
rect 14657 17697 14691 17731
rect 14933 17697 14967 17731
rect 15393 17697 15427 17731
rect 15577 17697 15611 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 15945 17697 15979 17731
rect 16129 17697 16163 17731
rect 16313 17697 16347 17731
rect 16589 17697 16623 17731
rect 18889 17697 18923 17731
rect 19073 17697 19107 17731
rect 19165 17697 19199 17731
rect 19257 17697 19291 17731
rect 19809 17697 19843 17731
rect 20729 17697 20763 17731
rect 20913 17697 20947 17731
rect 22201 17697 22235 17731
rect 22661 17697 22695 17731
rect 23121 17697 23155 17731
rect 23305 17697 23339 17731
rect 23397 17697 23431 17731
rect 23489 17697 23523 17731
rect 24317 17697 24351 17731
rect 24409 17697 24443 17731
rect 24501 17697 24535 17731
rect 24685 17697 24719 17731
rect 25145 17697 25179 17731
rect 25881 17697 25915 17731
rect 25973 17697 26007 17731
rect 26157 17697 26191 17731
rect 26249 17697 26283 17731
rect 27629 17697 27663 17731
rect 27721 17697 27755 17731
rect 27905 17697 27939 17731
rect 27997 17697 28031 17731
rect 28365 17697 28399 17731
rect 28549 17697 28583 17731
rect 28641 17697 28675 17731
rect 28733 17697 28767 17731
rect 30113 17697 30147 17731
rect 30297 17697 30331 17731
rect 30389 17697 30423 17731
rect 30481 17697 30515 17731
rect 3157 17629 3191 17663
rect 3617 17629 3651 17663
rect 4169 17629 4203 17663
rect 4261 17629 4295 17663
rect 4445 17629 4479 17663
rect 4629 17629 4663 17663
rect 6469 17629 6503 17663
rect 10241 17629 10275 17663
rect 11621 17629 11655 17663
rect 16405 17629 16439 17663
rect 16681 17629 16715 17663
rect 22477 17629 22511 17663
rect 24961 17629 24995 17663
rect 29469 17629 29503 17663
rect 3433 17561 3467 17595
rect 3893 17561 3927 17595
rect 7113 17561 7147 17595
rect 13369 17561 13403 17595
rect 25697 17561 25731 17595
rect 2421 17493 2455 17527
rect 5825 17493 5859 17527
rect 10977 17493 11011 17527
rect 14841 17493 14875 17527
rect 15025 17493 15059 17527
rect 15209 17493 15243 17527
rect 23029 17493 23063 17527
rect 23765 17493 23799 17527
rect 30021 17493 30055 17527
rect 30757 17493 30791 17527
rect 3709 17289 3743 17323
rect 3801 17289 3835 17323
rect 4721 17289 4755 17323
rect 5917 17289 5951 17323
rect 10885 17289 10919 17323
rect 11805 17289 11839 17323
rect 14013 17289 14047 17323
rect 16313 17289 16347 17323
rect 25697 17289 25731 17323
rect 27261 17289 27295 17323
rect 28825 17289 28859 17323
rect 31033 17289 31067 17323
rect 2789 17221 2823 17255
rect 4537 17221 4571 17255
rect 6101 17221 6135 17255
rect 9781 17221 9815 17255
rect 9873 17221 9907 17255
rect 14841 17221 14875 17255
rect 20269 17221 20303 17255
rect 1225 17153 1259 17187
rect 1409 17153 1443 17187
rect 3617 17153 3651 17187
rect 4629 17153 4663 17187
rect 5089 17153 5123 17187
rect 5733 17153 5767 17187
rect 6469 17153 6503 17187
rect 10701 17153 10735 17187
rect 15209 17153 15243 17187
rect 20913 17153 20947 17187
rect 21072 17153 21106 17187
rect 21465 17153 21499 17187
rect 21925 17153 21959 17187
rect 23581 17153 23615 17187
rect 23949 17153 23983 17187
rect 25145 17153 25179 17187
rect 30389 17153 30423 17187
rect 1317 17085 1351 17119
rect 1676 17085 1710 17119
rect 4077 17085 4111 17119
rect 4813 17085 4847 17119
rect 4997 17085 5031 17119
rect 5273 17085 5307 17119
rect 5457 17085 5491 17119
rect 5825 17085 5859 17119
rect 6009 17085 6043 17119
rect 6101 17085 6135 17119
rect 6285 17085 6319 17119
rect 6377 17085 6411 17119
rect 6561 17085 6595 17119
rect 8033 17085 8067 17119
rect 8125 17085 8159 17119
rect 8401 17085 8435 17119
rect 8668 17085 8702 17119
rect 10149 17085 10183 17119
rect 10241 17085 10275 17119
rect 10333 17085 10367 17119
rect 10517 17085 10551 17119
rect 10609 17085 10643 17119
rect 10885 17085 10919 17119
rect 11161 17085 11195 17119
rect 12918 17085 12952 17119
rect 13185 17085 13219 17119
rect 13645 17085 13679 17119
rect 13737 17085 13771 17119
rect 13829 17085 13863 17119
rect 14197 17085 14231 17119
rect 14381 17085 14415 17119
rect 14473 17085 14507 17119
rect 14565 17085 14599 17119
rect 14933 17085 14967 17119
rect 16681 17085 16715 17119
rect 18061 17085 18095 17119
rect 18245 17085 18279 17119
rect 18705 17085 18739 17119
rect 18797 17085 18831 17119
rect 18981 17085 19015 17119
rect 19073 17085 19107 17119
rect 19625 17085 19659 17119
rect 19993 17085 20027 17119
rect 21189 17085 21223 17119
rect 22109 17085 22143 17119
rect 23314 17085 23348 17119
rect 23857 17085 23891 17119
rect 24225 17085 24259 17119
rect 24409 17085 24443 17119
rect 24501 17085 24535 17119
rect 24593 17085 24627 17119
rect 25329 17085 25363 17119
rect 27169 17085 27203 17119
rect 27537 17085 27571 17119
rect 27629 17085 27663 17119
rect 27721 17085 27755 17119
rect 27905 17085 27939 17119
rect 28365 17085 28399 17119
rect 29009 17085 29043 17119
rect 29193 17085 29227 17119
rect 29285 17085 29319 17119
rect 29377 17085 29411 17119
rect 29745 17085 29779 17119
rect 30481 17085 30515 17119
rect 30573 17085 30607 17119
rect 30757 17085 30791 17119
rect 30849 17085 30883 17119
rect 31125 17085 31159 17119
rect 4261 17017 4295 17051
rect 5365 17017 5399 17051
rect 5595 17017 5629 17051
rect 19257 17017 19291 17051
rect 20085 17017 20119 17051
rect 27997 17017 28031 17051
rect 28181 17017 28215 17051
rect 28457 17017 28491 17051
rect 28641 17017 28675 17051
rect 3341 16949 3375 16983
rect 3985 16949 4019 16983
rect 11069 16949 11103 16983
rect 16865 16949 16899 16983
rect 18245 16949 18279 16983
rect 19441 16949 19475 16983
rect 22201 16949 22235 16983
rect 24869 16949 24903 16983
rect 25237 16949 25271 16983
rect 29653 16949 29687 16983
rect 31217 16949 31251 16983
rect 4169 16745 4203 16779
rect 4997 16745 5031 16779
rect 6193 16745 6227 16779
rect 6469 16745 6503 16779
rect 8953 16745 8987 16779
rect 14565 16745 14599 16779
rect 18521 16745 18555 16779
rect 18981 16745 19015 16779
rect 19165 16745 19199 16779
rect 22661 16745 22695 16779
rect 24501 16745 24535 16779
rect 28181 16745 28215 16779
rect 2881 16677 2915 16711
rect 3617 16677 3651 16711
rect 4537 16677 4571 16711
rect 6837 16677 6871 16711
rect 11345 16677 11379 16711
rect 13645 16677 13679 16711
rect 15678 16677 15712 16711
rect 23397 16677 23431 16711
rect 25706 16677 25740 16711
rect 30214 16677 30248 16711
rect 2421 16609 2455 16643
rect 2513 16609 2547 16643
rect 2605 16609 2639 16643
rect 2789 16609 2823 16643
rect 3525 16609 3559 16643
rect 3801 16609 3835 16643
rect 4077 16609 4111 16643
rect 4261 16609 4295 16643
rect 5181 16609 5215 16643
rect 5365 16609 5399 16643
rect 5549 16609 5583 16643
rect 5641 16609 5675 16643
rect 5825 16609 5859 16643
rect 6193 16609 6227 16643
rect 6653 16609 6687 16643
rect 9597 16609 9631 16643
rect 10793 16609 10827 16643
rect 10977 16609 11011 16643
rect 11161 16609 11195 16643
rect 11437 16609 11471 16643
rect 11621 16609 11655 16643
rect 12725 16609 12759 16643
rect 12817 16609 12851 16643
rect 15945 16609 15979 16643
rect 16221 16609 16255 16643
rect 16313 16609 16347 16643
rect 17785 16609 17819 16643
rect 17877 16609 17911 16643
rect 17969 16609 18003 16643
rect 18153 16609 18187 16643
rect 18613 16609 18647 16643
rect 19625 16609 19659 16643
rect 20085 16609 20119 16643
rect 21281 16609 21315 16643
rect 21537 16609 21571 16643
rect 22937 16609 22971 16643
rect 23029 16609 23063 16643
rect 23213 16609 23247 16643
rect 23305 16609 23339 16643
rect 23581 16609 23615 16643
rect 23765 16609 23799 16643
rect 23857 16609 23891 16643
rect 24041 16609 24075 16643
rect 24133 16609 24167 16643
rect 24225 16609 24259 16643
rect 25973 16609 26007 16643
rect 26157 16609 26191 16643
rect 26249 16609 26283 16643
rect 26709 16609 26743 16643
rect 27813 16609 27847 16643
rect 27997 16609 28031 16643
rect 28641 16609 28675 16643
rect 28733 16609 28767 16643
rect 28825 16609 28859 16643
rect 29009 16609 29043 16643
rect 30481 16609 30515 16643
rect 6377 16541 6411 16575
rect 9756 16541 9790 16575
rect 9873 16541 9907 16575
rect 10149 16541 10183 16575
rect 10609 16541 10643 16575
rect 11989 16541 12023 16575
rect 18337 16541 18371 16575
rect 22753 16541 22787 16575
rect 3985 16473 4019 16507
rect 4905 16473 4939 16507
rect 11437 16473 11471 16507
rect 19257 16473 19291 16507
rect 24593 16473 24627 16507
rect 28365 16473 28399 16507
rect 2145 16405 2179 16439
rect 17509 16405 17543 16439
rect 29101 16405 29135 16439
rect 4997 16201 5031 16235
rect 5549 16201 5583 16235
rect 8953 16201 8987 16235
rect 17509 16201 17543 16235
rect 18429 16201 18463 16235
rect 19073 16201 19107 16235
rect 25329 16201 25363 16235
rect 27077 16201 27111 16235
rect 28089 16201 28123 16235
rect 3065 16133 3099 16167
rect 4629 16133 4663 16167
rect 21649 16133 21683 16167
rect 22569 16133 22603 16167
rect 29009 16133 29043 16167
rect 4261 16065 4295 16099
rect 19533 16065 19567 16099
rect 19625 16065 19659 16099
rect 21005 16065 21039 16099
rect 21189 16065 21223 16099
rect 24685 16065 24719 16099
rect 29469 16065 29503 16099
rect 29561 16065 29595 16099
rect 1409 15997 1443 16031
rect 1501 15997 1535 16031
rect 1685 15997 1719 16031
rect 1952 15997 1986 16031
rect 5365 15997 5399 16031
rect 5641 15997 5675 16031
rect 6745 15997 6779 16031
rect 8033 15997 8067 16031
rect 8585 15997 8619 16031
rect 9321 15997 9355 16031
rect 9413 15997 9447 16031
rect 9505 15997 9539 16031
rect 9689 15997 9723 16031
rect 10609 15997 10643 16031
rect 11069 15997 11103 16031
rect 11989 15997 12023 16031
rect 13001 15997 13035 16031
rect 13829 15997 13863 16031
rect 13921 15997 13955 16031
rect 14013 15997 14047 16031
rect 14197 15997 14231 16031
rect 17141 15997 17175 16031
rect 17647 15997 17681 16031
rect 17785 15997 17819 16031
rect 18337 15997 18371 16031
rect 19441 15997 19475 16031
rect 19901 15997 19935 16031
rect 21281 15997 21315 16031
rect 21925 15997 21959 16031
rect 22017 15997 22051 16031
rect 22201 15997 22235 16031
rect 22293 15997 22327 16031
rect 22385 15997 22419 16031
rect 22753 15997 22787 16031
rect 24041 15997 24075 16031
rect 24225 15997 24259 16031
rect 24869 15997 24903 16031
rect 25513 15997 25547 16031
rect 25605 15997 25639 16031
rect 25789 15997 25823 16031
rect 25881 15997 25915 16031
rect 26065 15997 26099 16031
rect 27261 15997 27295 16031
rect 27537 15997 27571 16031
rect 27629 15997 27663 16031
rect 27813 15997 27847 16031
rect 27905 15997 27939 16031
rect 28825 15997 28859 16031
rect 30021 15997 30055 16031
rect 4997 15929 5031 15963
rect 5825 15929 5859 15963
rect 6653 15929 6687 15963
rect 8769 15929 8803 15963
rect 10057 15929 10091 15963
rect 18061 15929 18095 15963
rect 18153 15929 18187 15963
rect 20729 15929 20763 15963
rect 24409 15929 24443 15963
rect 26801 15929 26835 15963
rect 27445 15929 27479 15963
rect 4721 15861 4755 15895
rect 4813 15861 4847 15895
rect 7389 15861 7423 15895
rect 8125 15861 8159 15895
rect 9045 15861 9079 15895
rect 11713 15861 11747 15895
rect 13093 15861 13127 15895
rect 13553 15861 13587 15895
rect 17233 15861 17267 15895
rect 21741 15861 21775 15895
rect 22937 15861 22971 15895
rect 24777 15861 24811 15895
rect 25237 15861 25271 15895
rect 28181 15861 28215 15895
rect 29377 15861 29411 15895
rect 29929 15861 29963 15895
rect 2697 15657 2731 15691
rect 7205 15657 7239 15691
rect 7297 15657 7331 15691
rect 10149 15657 10183 15691
rect 11621 15657 11655 15691
rect 12173 15657 12207 15691
rect 18613 15657 18647 15691
rect 18981 15657 19015 15691
rect 19073 15657 19107 15691
rect 21097 15657 21131 15691
rect 21925 15657 21959 15691
rect 22201 15657 22235 15691
rect 24501 15657 24535 15691
rect 28457 15657 28491 15691
rect 29929 15657 29963 15691
rect 30389 15657 30423 15691
rect 5825 15589 5859 15623
rect 16497 15589 16531 15623
rect 17500 15589 17534 15623
rect 19441 15589 19475 15623
rect 19809 15589 19843 15623
rect 20177 15589 20211 15623
rect 28365 15589 28399 15623
rect 29570 15589 29604 15623
rect 1317 15521 1351 15555
rect 2789 15521 2823 15555
rect 3157 15521 3191 15555
rect 4445 15521 4479 15555
rect 5457 15521 5491 15555
rect 6561 15521 6595 15555
rect 8769 15521 8803 15555
rect 9036 15521 9070 15555
rect 10425 15521 10459 15555
rect 10701 15521 10735 15555
rect 11805 15521 11839 15555
rect 11989 15521 12023 15555
rect 13389 15521 13423 15555
rect 13645 15521 13679 15555
rect 13829 15521 13863 15555
rect 14013 15521 14047 15555
rect 14105 15521 14139 15555
rect 14197 15521 14231 15555
rect 14841 15521 14875 15555
rect 14933 15521 14967 15555
rect 16772 15521 16806 15555
rect 16865 15521 16899 15555
rect 16957 15521 16991 15555
rect 17141 15521 17175 15555
rect 17233 15521 17267 15555
rect 18889 15521 18923 15555
rect 19717 15521 19751 15555
rect 19993 15521 20027 15555
rect 20453 15521 20487 15555
rect 20637 15521 20671 15555
rect 20729 15521 20763 15555
rect 20867 15521 20901 15555
rect 21281 15521 21315 15555
rect 21465 15521 21499 15555
rect 21557 15521 21591 15555
rect 21649 15521 21683 15555
rect 22017 15521 22051 15555
rect 23949 15521 23983 15555
rect 24317 15521 24351 15555
rect 25145 15521 25179 15555
rect 27721 15521 27755 15555
rect 27905 15521 27939 15555
rect 27997 15521 28031 15555
rect 28089 15521 28123 15555
rect 29837 15521 29871 15555
rect 30297 15521 30331 15555
rect 2237 15453 2271 15487
rect 2973 15453 3007 15487
rect 3801 15453 3835 15487
rect 7389 15453 7423 15487
rect 10517 15453 10551 15487
rect 10977 15453 11011 15487
rect 19625 15453 19659 15487
rect 30481 15453 30515 15487
rect 2329 15385 2363 15419
rect 10241 15385 10275 15419
rect 15025 15385 15059 15419
rect 1409 15317 1443 15351
rect 1593 15317 1627 15351
rect 6837 15317 6871 15351
rect 10425 15317 10459 15351
rect 12265 15317 12299 15351
rect 14473 15317 14507 15351
rect 14657 15317 14691 15351
rect 24133 15317 24167 15351
rect 25053 15317 25087 15351
rect 9781 15113 9815 15147
rect 12081 15113 12115 15147
rect 14013 15113 14047 15147
rect 16681 15113 16715 15147
rect 17049 15113 17083 15147
rect 17785 15113 17819 15147
rect 17969 15113 18003 15147
rect 19349 15113 19383 15147
rect 19901 15113 19935 15147
rect 21373 15113 21407 15147
rect 21741 15113 21775 15147
rect 26157 15113 26191 15147
rect 28273 15113 28307 15147
rect 30389 15113 30423 15147
rect 4353 15045 4387 15079
rect 20085 15045 20119 15079
rect 1593 14977 1627 15011
rect 3709 14977 3743 15011
rect 4077 14977 4111 15011
rect 7113 14977 7147 15011
rect 7297 14977 7331 15011
rect 11161 14977 11195 15011
rect 14105 14977 14139 15011
rect 19809 14977 19843 15011
rect 1317 14909 1351 14943
rect 3433 14909 3467 14943
rect 3617 14909 3651 14943
rect 3801 14909 3835 14943
rect 3985 14909 4019 14943
rect 4261 14909 4295 14943
rect 4445 14909 4479 14943
rect 4537 14909 4571 14943
rect 4721 14909 4755 14943
rect 7205 14909 7239 14943
rect 8953 14909 8987 14943
rect 9321 14909 9355 14943
rect 9413 14909 9447 14943
rect 9505 14909 9539 14943
rect 9689 14909 9723 14943
rect 11529 14909 11563 14943
rect 11621 14909 11655 14943
rect 11713 14909 11747 14943
rect 11897 14909 11931 14943
rect 12173 14909 12207 14943
rect 12725 14909 12759 14943
rect 12909 14909 12943 14943
rect 13001 14909 13035 14943
rect 13093 14909 13127 14943
rect 13645 14909 13679 14943
rect 14372 14909 14406 14943
rect 15577 14909 15611 14943
rect 16313 14909 16347 14943
rect 16681 14909 16715 14943
rect 16865 14909 16899 14943
rect 17325 14909 17359 14943
rect 17417 14909 17451 14943
rect 17785 14909 17819 14943
rect 18049 14909 18083 14943
rect 18245 14909 18279 14943
rect 18705 14909 18739 14943
rect 18798 14909 18832 14943
rect 18935 14909 18969 14943
rect 19073 14909 19107 14943
rect 19170 14909 19204 14943
rect 19912 14909 19946 14943
rect 20821 14909 20855 14943
rect 20913 14909 20947 14943
rect 21097 14909 21131 14943
rect 21373 14909 21407 14943
rect 21557 14909 21591 14943
rect 23673 14909 23707 14943
rect 24041 14909 24075 14943
rect 24133 14909 24167 14943
rect 24317 14909 24351 14943
rect 24409 14909 24443 14943
rect 24685 14909 24719 14943
rect 24869 14909 24903 14943
rect 24961 14909 24995 14943
rect 25053 14909 25087 14943
rect 25651 14909 25685 14943
rect 25789 14909 25823 14943
rect 25881 14909 25915 14943
rect 26065 14909 26099 14943
rect 26709 14909 26743 14943
rect 27169 14909 27203 14943
rect 27261 14909 27295 14943
rect 27353 14909 27387 14943
rect 27537 14909 27571 14943
rect 28457 14909 28491 14943
rect 28549 14909 28583 14943
rect 28733 14909 28767 14943
rect 28825 14909 28859 14943
rect 29009 14909 29043 14943
rect 29193 14909 29227 14943
rect 29285 14909 29319 14943
rect 29377 14909 29411 14943
rect 29745 14909 29779 14943
rect 29929 14909 29963 14943
rect 30021 14909 30055 14943
rect 30113 14909 30147 14943
rect 1860 14841 1894 14875
rect 3249 14841 3283 14875
rect 6846 14841 6880 14875
rect 10916 14841 10950 14875
rect 11253 14841 11287 14875
rect 13829 14841 13863 14875
rect 19625 14841 19659 14875
rect 20361 14841 20395 14875
rect 21281 14841 21315 14875
rect 23489 14841 23523 14875
rect 27813 14841 27847 14875
rect 27997 14841 28031 14875
rect 28181 14841 28215 14875
rect 1409 14773 1443 14807
rect 2973 14773 3007 14807
rect 5365 14773 5399 14807
rect 5733 14773 5767 14807
rect 8861 14773 8895 14807
rect 9045 14773 9079 14807
rect 13369 14773 13403 14807
rect 15485 14773 15519 14807
rect 15761 14773 15795 14807
rect 16497 14773 16531 14807
rect 18153 14773 18187 14807
rect 23305 14773 23339 14807
rect 23857 14773 23891 14807
rect 25329 14773 25363 14807
rect 25421 14773 25455 14807
rect 26893 14773 26927 14807
rect 29653 14773 29687 14807
rect 2881 14569 2915 14603
rect 5089 14569 5123 14603
rect 6285 14569 6319 14603
rect 7021 14569 7055 14603
rect 13277 14569 13311 14603
rect 15117 14569 15151 14603
rect 17509 14569 17543 14603
rect 18797 14569 18831 14603
rect 21005 14569 21039 14603
rect 23765 14569 23799 14603
rect 24225 14569 24259 14603
rect 26249 14569 26283 14603
rect 26893 14569 26927 14603
rect 27353 14569 27387 14603
rect 29469 14569 29503 14603
rect 29561 14569 29595 14603
rect 29929 14569 29963 14603
rect 1746 14501 1780 14535
rect 9474 14501 9508 14535
rect 12081 14501 12115 14535
rect 12265 14501 12299 14535
rect 13982 14501 14016 14535
rect 19809 14501 19843 14535
rect 22569 14501 22603 14535
rect 22753 14501 22787 14535
rect 23857 14501 23891 14535
rect 25136 14501 25170 14535
rect 1501 14433 1535 14467
rect 3065 14433 3099 14467
rect 3157 14433 3191 14467
rect 7389 14433 7423 14467
rect 8401 14433 8435 14467
rect 9229 14433 9263 14467
rect 12449 14433 12483 14467
rect 12541 14433 12575 14467
rect 12725 14433 12759 14467
rect 13461 14433 13495 14467
rect 13645 14433 13679 14467
rect 15209 14433 15243 14467
rect 15363 14433 15397 14467
rect 16773 14433 16807 14467
rect 17141 14433 17175 14467
rect 17693 14433 17727 14467
rect 18153 14433 18187 14467
rect 18429 14433 18463 14467
rect 18613 14433 18647 14467
rect 19993 14433 20027 14467
rect 20085 14433 20119 14467
rect 20269 14433 20303 14467
rect 20729 14433 20763 14467
rect 21833 14433 21867 14467
rect 21925 14433 21959 14467
rect 22017 14433 22051 14467
rect 22201 14433 22235 14467
rect 22385 14433 22419 14467
rect 22477 14433 22511 14467
rect 22661 14433 22695 14467
rect 23029 14433 23063 14467
rect 23121 14433 23155 14467
rect 23213 14433 23247 14467
rect 23397 14433 23431 14467
rect 24409 14433 24443 14467
rect 24869 14433 24903 14467
rect 26985 14433 27019 14467
rect 27537 14433 27571 14467
rect 27721 14433 27755 14467
rect 27997 14433 28031 14467
rect 28181 14433 28215 14467
rect 28365 14433 28399 14467
rect 28457 14433 28491 14467
rect 28549 14433 28583 14467
rect 30205 14433 30239 14467
rect 30297 14433 30331 14467
rect 30481 14433 30515 14467
rect 30573 14433 30607 14467
rect 30665 14433 30699 14467
rect 30757 14433 30791 14467
rect 30941 14433 30975 14467
rect 31033 14433 31067 14467
rect 6377 14365 6411 14399
rect 6469 14365 6503 14399
rect 6837 14365 6871 14399
rect 7297 14365 7331 14399
rect 7849 14365 7883 14399
rect 7941 14365 7975 14399
rect 8217 14365 8251 14399
rect 11529 14365 11563 14399
rect 13737 14365 13771 14399
rect 15577 14365 15611 14399
rect 17785 14365 17819 14399
rect 20545 14365 20579 14399
rect 21097 14365 21131 14399
rect 21557 14365 21591 14399
rect 23673 14365 23707 14399
rect 27077 14365 27111 14399
rect 29285 14365 29319 14399
rect 3065 14297 3099 14331
rect 4905 14297 4939 14331
rect 5457 14297 5491 14331
rect 10609 14297 10643 14331
rect 12541 14297 12575 14331
rect 16957 14297 16991 14331
rect 31217 14297 31251 14331
rect 5089 14229 5123 14263
rect 5917 14229 5951 14263
rect 10977 14229 11011 14263
rect 17325 14229 17359 14263
rect 17693 14229 17727 14263
rect 20453 14229 20487 14263
rect 21281 14229 21315 14263
rect 21741 14229 21775 14263
rect 24685 14229 24719 14263
rect 26525 14229 26559 14263
rect 27905 14229 27939 14263
rect 28825 14229 28859 14263
rect 30021 14229 30055 14263
rect 7021 14025 7055 14059
rect 9965 14025 9999 14059
rect 13921 14025 13955 14059
rect 15025 14025 15059 14059
rect 15209 14025 15243 14059
rect 18153 14025 18187 14059
rect 20085 14025 20119 14059
rect 25237 14025 25271 14059
rect 27997 14025 28031 14059
rect 29837 14025 29871 14059
rect 30573 14025 30607 14059
rect 17509 13957 17543 13991
rect 17601 13957 17635 13991
rect 20361 13957 20395 13991
rect 20545 13957 20579 13991
rect 20913 13957 20947 13991
rect 4813 13889 4847 13923
rect 5641 13889 5675 13923
rect 7757 13889 7791 13923
rect 15393 13889 15427 13923
rect 16405 13889 16439 13923
rect 20821 13889 20855 13923
rect 22293 13889 22327 13923
rect 22477 13889 22511 13923
rect 23029 13889 23063 13923
rect 25973 13889 26007 13923
rect 27353 13889 27387 13923
rect 27905 13889 27939 13923
rect 29285 13889 29319 13923
rect 2605 13821 2639 13855
rect 2881 13821 2915 13855
rect 3065 13821 3099 13855
rect 3709 13821 3743 13855
rect 3893 13821 3927 13855
rect 4169 13821 4203 13855
rect 4353 13821 4387 13855
rect 4721 13821 4755 13855
rect 5211 13821 5245 13855
rect 5365 13821 5399 13855
rect 5908 13821 5942 13855
rect 9689 13821 9723 13855
rect 10149 13821 10183 13855
rect 10333 13821 10367 13855
rect 10701 13821 10735 13855
rect 11253 13821 11287 13855
rect 14013 13821 14047 13855
rect 15209 13821 15243 13855
rect 16313 13821 16347 13855
rect 16497 13821 16531 13855
rect 17693 13821 17727 13855
rect 18061 13821 18095 13855
rect 18153 13821 18187 13855
rect 22026 13821 22060 13855
rect 22385 13821 22419 13855
rect 23305 13821 23339 13855
rect 23397 13821 23431 13855
rect 23489 13821 23523 13855
rect 23673 13821 23707 13855
rect 23857 13821 23891 13855
rect 24113 13821 24147 13855
rect 25697 13821 25731 13855
rect 26709 13821 26743 13855
rect 26893 13821 26927 13855
rect 26985 13821 27019 13855
rect 27077 13821 27111 13855
rect 28549 13821 28583 13855
rect 29929 13821 29963 13855
rect 30113 13821 30147 13855
rect 30205 13821 30239 13855
rect 30297 13821 30331 13855
rect 7573 13753 7607 13787
rect 9505 13753 9539 13787
rect 9873 13753 9907 13787
rect 15485 13753 15519 13787
rect 17141 13753 17175 13787
rect 19901 13753 19935 13787
rect 20117 13753 20151 13787
rect 27537 13753 27571 13787
rect 27721 13753 27755 13787
rect 29469 13753 29503 13787
rect 2513 13685 2547 13719
rect 2973 13685 3007 13719
rect 4997 13685 5031 13719
rect 7205 13685 7239 13719
rect 7665 13685 7699 13719
rect 10517 13685 10551 13719
rect 11161 13685 11195 13719
rect 18337 13685 18371 13719
rect 20269 13685 20303 13719
rect 25329 13685 25363 13719
rect 25789 13685 25823 13719
rect 29377 13685 29411 13719
rect 3801 13481 3835 13515
rect 4077 13481 4111 13515
rect 7481 13481 7515 13515
rect 12357 13481 12391 13515
rect 12909 13481 12943 13515
rect 14473 13481 14507 13515
rect 18153 13481 18187 13515
rect 24133 13481 24167 13515
rect 28733 13481 28767 13515
rect 29745 13481 29779 13515
rect 2596 13413 2630 13447
rect 3985 13413 4019 13447
rect 4353 13413 4387 13447
rect 10609 13413 10643 13447
rect 11222 13413 11256 13447
rect 13185 13413 13219 13447
rect 24317 13413 24351 13447
rect 25053 13413 25087 13447
rect 25697 13413 25731 13447
rect 25881 13413 25915 13447
rect 26065 13413 26099 13447
rect 27077 13413 27111 13447
rect 2329 13345 2363 13379
rect 4169 13345 4203 13379
rect 5457 13345 5491 13379
rect 6092 13345 6126 13379
rect 8309 13343 8343 13377
rect 9321 13345 9355 13379
rect 9505 13345 9539 13379
rect 9965 13345 9999 13379
rect 10149 13345 10183 13379
rect 10241 13345 10275 13379
rect 10333 13345 10367 13379
rect 10977 13345 11011 13379
rect 12725 13345 12759 13379
rect 13369 13345 13403 13379
rect 13645 13345 13679 13379
rect 13829 13345 13863 13379
rect 13921 13345 13955 13379
rect 14013 13345 14047 13379
rect 14657 13345 14691 13379
rect 15209 13345 15243 13379
rect 15393 13345 15427 13379
rect 16681 13345 16715 13379
rect 17049 13345 17083 13379
rect 17693 13345 17727 13379
rect 18613 13345 18647 13379
rect 21465 13345 21499 13379
rect 23949 13345 23983 13379
rect 24225 13345 24259 13379
rect 24961 13345 24995 13379
rect 25237 13345 25271 13379
rect 25329 13345 25363 13379
rect 25513 13345 25547 13379
rect 25605 13345 25639 13379
rect 26525 13345 26559 13379
rect 26617 13345 26651 13379
rect 26801 13345 26835 13379
rect 26893 13345 26927 13379
rect 27353 13345 27387 13379
rect 27620 13345 27654 13379
rect 28917 13345 28951 13379
rect 29101 13345 29135 13379
rect 29193 13345 29227 13379
rect 29285 13345 29319 13379
rect 30481 13345 30515 13379
rect 5549 13277 5583 13311
rect 5825 13277 5859 13311
rect 8033 13277 8067 13311
rect 13093 13277 13127 13311
rect 13553 13277 13587 13311
rect 17785 13277 17819 13311
rect 18889 13277 18923 13311
rect 21741 13277 21775 13311
rect 21833 13277 21867 13311
rect 30389 13277 30423 13311
rect 31033 13277 31067 13311
rect 18337 13209 18371 13243
rect 18797 13209 18831 13243
rect 23765 13209 23799 13243
rect 3709 13141 3743 13175
rect 7205 13141 7239 13175
rect 8401 13141 8435 13175
rect 9137 13141 9171 13175
rect 12725 13141 12759 13175
rect 14289 13141 14323 13175
rect 15301 13141 15335 13175
rect 16589 13141 16623 13175
rect 17141 13141 17175 13175
rect 17509 13141 17543 13175
rect 18153 13141 18187 13175
rect 18429 13141 18463 13175
rect 29561 13141 29595 13175
rect 9505 12937 9539 12971
rect 12909 12937 12943 12971
rect 15577 12937 15611 12971
rect 18061 12937 18095 12971
rect 18889 12937 18923 12971
rect 19073 12937 19107 12971
rect 30665 12937 30699 12971
rect 3065 12869 3099 12903
rect 15485 12869 15519 12903
rect 16313 12869 16347 12903
rect 17463 12869 17497 12903
rect 17601 12869 17635 12903
rect 17877 12869 17911 12903
rect 26065 12869 26099 12903
rect 13737 12801 13771 12835
rect 28733 12801 28767 12835
rect 29285 12801 29319 12835
rect 1409 12733 1443 12767
rect 1501 12733 1535 12767
rect 1685 12733 1719 12767
rect 3341 12733 3375 12767
rect 4537 12733 4571 12767
rect 7021 12733 7055 12767
rect 7113 12733 7147 12767
rect 8125 12733 8159 12767
rect 8677 12733 8711 12767
rect 8769 12733 8803 12767
rect 8861 12733 8895 12767
rect 9045 12733 9079 12767
rect 10057 12733 10091 12767
rect 11375 12733 11409 12767
rect 11529 12733 11563 12767
rect 12081 12733 12115 12767
rect 12265 12733 12299 12767
rect 12541 12733 12575 12767
rect 12633 12733 12667 12767
rect 12725 12733 12759 12767
rect 13645 12733 13679 12767
rect 13921 12733 13955 12767
rect 14105 12733 14139 12767
rect 14372 12733 14406 12767
rect 15577 12733 15611 12767
rect 15761 12733 15795 12767
rect 15853 12733 15887 12767
rect 16129 12733 16163 12767
rect 17233 12733 17267 12767
rect 17325 12733 17359 12767
rect 17785 12733 17819 12767
rect 18061 12733 18095 12767
rect 18153 12733 18187 12767
rect 25973 12733 26007 12767
rect 26157 12733 26191 12767
rect 26433 12733 26467 12767
rect 26709 12733 26743 12767
rect 28641 12733 28675 12767
rect 29009 12733 29043 12767
rect 29552 12733 29586 12767
rect 1952 12665 1986 12699
rect 3985 12665 4019 12699
rect 7297 12665 7331 12699
rect 7573 12665 7607 12699
rect 13553 12665 13587 12699
rect 17693 12665 17727 12699
rect 18521 12665 18555 12699
rect 18705 12665 18739 12699
rect 3893 12597 3927 12631
rect 6929 12597 6963 12631
rect 7481 12597 7515 12631
rect 8401 12597 8435 12631
rect 11161 12597 11195 12631
rect 12265 12597 12299 12631
rect 13829 12597 13863 12631
rect 16037 12597 16071 12631
rect 16589 12597 16623 12631
rect 18905 12597 18939 12631
rect 26341 12597 26375 12631
rect 26617 12597 26651 12631
rect 29101 12597 29135 12631
rect 4077 12393 4111 12427
rect 8125 12393 8159 12427
rect 9781 12393 9815 12427
rect 13645 12393 13679 12427
rect 14289 12393 14323 12427
rect 14473 12393 14507 12427
rect 17509 12393 17543 12427
rect 19165 12393 19199 12427
rect 19809 12393 19843 12427
rect 25605 12393 25639 12427
rect 27905 12393 27939 12427
rect 30757 12393 30791 12427
rect 2865 12325 2899 12359
rect 3065 12325 3099 12359
rect 8484 12325 8518 12359
rect 11989 12325 12023 12359
rect 18052 12325 18086 12359
rect 22063 12325 22097 12359
rect 22201 12325 22235 12359
rect 22819 12325 22853 12359
rect 26091 12325 26125 12359
rect 29622 12325 29656 12359
rect 2329 12257 2363 12291
rect 3801 12257 3835 12291
rect 3893 12257 3927 12291
rect 4169 12257 4203 12291
rect 5089 12257 5123 12291
rect 5243 12257 5277 12291
rect 6039 12257 6073 12291
rect 6193 12257 6227 12291
rect 6745 12257 6779 12291
rect 7012 12257 7046 12291
rect 8217 12257 8251 12291
rect 9873 12257 9907 12291
rect 10609 12257 10643 12291
rect 10793 12257 10827 12291
rect 11161 12257 11195 12291
rect 11345 12257 11379 12291
rect 11713 12257 11747 12291
rect 12081 12257 12115 12291
rect 12449 12257 12483 12291
rect 12725 12257 12759 12291
rect 12909 12257 12943 12291
rect 13461 12257 13495 12291
rect 14381 12257 14415 12291
rect 14687 12257 14721 12291
rect 14841 12257 14875 12291
rect 15577 12257 15611 12291
rect 16129 12257 16163 12291
rect 16385 12257 16419 12291
rect 17785 12257 17819 12291
rect 19441 12257 19475 12291
rect 19717 12257 19751 12291
rect 19993 12257 20027 12291
rect 20177 12257 20211 12291
rect 22293 12257 22327 12291
rect 22384 12247 22418 12281
rect 22661 12257 22695 12291
rect 22937 12257 22971 12291
rect 23029 12257 23063 12291
rect 23121 12257 23155 12291
rect 25237 12257 25271 12291
rect 25789 12257 25823 12291
rect 25881 12257 25915 12291
rect 25973 12257 26007 12291
rect 26249 12257 26283 12291
rect 26433 12257 26467 12291
rect 26617 12257 26651 12291
rect 26709 12257 26743 12291
rect 26801 12257 26835 12291
rect 27261 12257 27295 12291
rect 27813 12257 27847 12291
rect 29377 12257 29411 12291
rect 1961 12189 1995 12223
rect 2237 12189 2271 12223
rect 3249 12189 3283 12223
rect 19625 12189 19659 12223
rect 21925 12189 21959 12223
rect 25421 12189 25455 12223
rect 27537 12189 27571 12223
rect 5825 12121 5859 12155
rect 15761 12121 15795 12155
rect 19257 12121 19291 12155
rect 20361 12121 20395 12155
rect 27077 12121 27111 12155
rect 2697 12053 2731 12087
rect 2881 12053 2915 12087
rect 3893 12053 3927 12087
rect 5273 12053 5307 12087
rect 9597 12053 9631 12087
rect 10793 12053 10827 12087
rect 11437 12053 11471 12087
rect 22569 12053 22603 12087
rect 23305 12053 23339 12087
rect 25053 12053 25087 12087
rect 3065 11849 3099 11883
rect 4169 11849 4203 11883
rect 4629 11849 4663 11883
rect 7573 11849 7607 11883
rect 16589 11849 16623 11883
rect 23121 11849 23155 11883
rect 26617 11849 26651 11883
rect 28273 11849 28307 11883
rect 4997 11781 5031 11815
rect 16037 11781 16071 11815
rect 20545 11781 20579 11815
rect 3985 11713 4019 11747
rect 4721 11713 4755 11747
rect 5181 11713 5215 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 21281 11713 21315 11747
rect 23581 11713 23615 11747
rect 1317 11645 1351 11679
rect 1409 11645 1443 11679
rect 1501 11645 1535 11679
rect 1685 11645 1719 11679
rect 3249 11645 3283 11679
rect 3433 11645 3467 11679
rect 3893 11645 3927 11679
rect 4169 11645 4203 11679
rect 4445 11645 4479 11679
rect 4629 11645 4663 11679
rect 5273 11645 5307 11679
rect 5421 11645 5455 11679
rect 5549 11645 5583 11679
rect 5738 11645 5772 11679
rect 7849 11645 7883 11679
rect 7941 11645 7975 11679
rect 8033 11645 8067 11679
rect 8217 11645 8251 11679
rect 9965 11645 9999 11679
rect 10149 11645 10183 11679
rect 10241 11645 10275 11679
rect 11253 11645 11287 11679
rect 11437 11645 11471 11679
rect 11713 11645 11747 11679
rect 12633 11645 12667 11679
rect 13093 11645 13127 11679
rect 13369 11645 13403 11679
rect 18337 11645 18371 11679
rect 18429 11645 18463 11679
rect 18889 11645 18923 11679
rect 19145 11645 19179 11679
rect 20361 11645 20395 11679
rect 21465 11645 21499 11679
rect 21741 11645 21775 11679
rect 23397 11645 23431 11679
rect 23857 11645 23891 11679
rect 24685 11645 24719 11679
rect 24777 11645 24811 11679
rect 24961 11645 24995 11679
rect 25217 11645 25251 11679
rect 27730 11645 27764 11679
rect 27997 11645 28031 11679
rect 28549 11645 28583 11679
rect 28641 11645 28675 11679
rect 29653 11645 29687 11679
rect 30573 11645 30607 11679
rect 1952 11577 1986 11611
rect 3341 11577 3375 11611
rect 5641 11577 5675 11611
rect 9698 11577 9732 11611
rect 17877 11577 17911 11611
rect 21649 11577 21683 11611
rect 21986 11577 22020 11611
rect 28181 11577 28215 11611
rect 1225 11509 1259 11543
rect 4353 11509 4387 11543
rect 5917 11509 5951 11543
rect 8585 11509 8619 11543
rect 11897 11509 11931 11543
rect 15669 11509 15703 11543
rect 20269 11509 20303 11543
rect 23213 11509 23247 11543
rect 23949 11509 23983 11543
rect 26341 11509 26375 11543
rect 29561 11509 29595 11543
rect 29929 11509 29963 11543
rect 5549 11305 5583 11339
rect 8769 11305 8803 11339
rect 15577 11305 15611 11339
rect 19165 11305 19199 11339
rect 21925 11305 21959 11339
rect 25329 11305 25363 11339
rect 26249 11305 26283 11339
rect 27813 11305 27847 11339
rect 9689 11237 9723 11271
rect 19671 11237 19705 11271
rect 23222 11237 23256 11271
rect 25697 11237 25731 11271
rect 26700 11237 26734 11271
rect 29285 11237 29319 11271
rect 29622 11237 29656 11271
rect 1869 11169 1903 11203
rect 2136 11169 2170 11203
rect 4261 11169 4295 11203
rect 4721 11169 4755 11203
rect 5365 11169 5399 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 6009 11169 6043 11203
rect 6101 11169 6135 11203
rect 6377 11169 6411 11203
rect 9045 11169 9079 11203
rect 9137 11169 9171 11203
rect 9229 11169 9263 11203
rect 9413 11169 9447 11203
rect 9873 11169 9907 11203
rect 15853 11169 15887 11203
rect 16405 11169 16439 11203
rect 19349 11169 19383 11203
rect 19441 11169 19475 11203
rect 19533 11169 19567 11203
rect 19809 11169 19843 11203
rect 20085 11169 20119 11203
rect 20177 11169 20211 11203
rect 20269 11169 20303 11203
rect 20387 11169 20421 11203
rect 22017 11169 22051 11203
rect 23489 11169 23523 11203
rect 25513 11169 25547 11203
rect 25605 11169 25639 11203
rect 25815 11169 25849 11203
rect 25973 11169 26007 11203
rect 26065 11169 26099 11203
rect 26249 11169 26283 11203
rect 26433 11169 26467 11203
rect 28641 11169 28675 11203
rect 28825 11169 28859 11203
rect 28917 11169 28951 11203
rect 29009 11169 29043 11203
rect 29377 11169 29411 11203
rect 3893 11101 3927 11135
rect 4445 11101 4479 11135
rect 4813 11101 4847 11135
rect 6285 11101 6319 11135
rect 9505 11101 9539 11135
rect 16221 11101 16255 11135
rect 20545 11101 20579 11135
rect 3341 11033 3375 11067
rect 5181 11033 5215 11067
rect 22109 11033 22143 11067
rect 30757 11033 30791 11067
rect 3249 10965 3283 10999
rect 4077 10965 4111 10999
rect 16589 10965 16623 10999
rect 19901 10965 19935 10999
rect 2421 10761 2455 10795
rect 5641 10761 5675 10795
rect 16037 10761 16071 10795
rect 20913 10761 20947 10795
rect 26893 10761 26927 10795
rect 29193 10761 29227 10795
rect 26433 10693 26467 10727
rect 2697 10625 2731 10659
rect 4537 10625 4571 10659
rect 18889 10625 18923 10659
rect 19533 10625 19567 10659
rect 24501 10625 24535 10659
rect 2237 10557 2271 10591
rect 2421 10557 2455 10591
rect 2605 10557 2639 10591
rect 2789 10557 2823 10591
rect 3433 10557 3467 10591
rect 4445 10557 4479 10591
rect 5825 10557 5859 10591
rect 6009 10557 6043 10591
rect 6193 10557 6227 10591
rect 8033 10557 8067 10591
rect 8677 10557 8711 10591
rect 8769 10557 8803 10591
rect 8861 10557 8895 10591
rect 9045 10557 9079 10591
rect 9321 10557 9355 10591
rect 10241 10557 10275 10591
rect 10885 10557 10919 10591
rect 12725 10557 12759 10591
rect 12909 10557 12943 10591
rect 13001 10557 13035 10591
rect 13737 10557 13771 10591
rect 14289 10557 14323 10591
rect 14381 10557 14415 10591
rect 14657 10557 14691 10591
rect 16129 10557 16163 10591
rect 18797 10557 18831 10591
rect 19073 10557 19107 10591
rect 19257 10557 19291 10591
rect 21189 10557 21223 10591
rect 24041 10557 24075 10591
rect 25237 10557 25271 10591
rect 25605 10557 25639 10591
rect 26985 10557 27019 10591
rect 29101 10557 29135 10591
rect 29285 10557 29319 10591
rect 29745 10557 29779 10591
rect 29837 10557 29871 10591
rect 29929 10557 29963 10591
rect 30113 10557 30147 10591
rect 30757 10557 30791 10591
rect 5917 10489 5951 10523
rect 7849 10489 7883 10523
rect 8217 10489 8251 10523
rect 10425 10489 10459 10523
rect 11069 10489 11103 10523
rect 12458 10489 12492 10523
rect 14924 10489 14958 10523
rect 16396 10489 16430 10523
rect 19441 10489 19475 10523
rect 19778 10489 19812 10523
rect 24133 10489 24167 10523
rect 24225 10489 24259 10523
rect 24363 10489 24397 10523
rect 26617 10489 26651 10523
rect 3341 10421 3375 10455
rect 8401 10421 8435 10455
rect 9229 10421 9263 10455
rect 10609 10421 10643 10455
rect 11253 10421 11287 10455
rect 11345 10421 11379 10455
rect 13645 10421 13679 10455
rect 14565 10421 14599 10455
rect 17509 10421 17543 10455
rect 21097 10421 21131 10455
rect 23857 10421 23891 10455
rect 24685 10421 24719 10455
rect 25513 10421 25547 10455
rect 30021 10421 30055 10455
rect 30849 10421 30883 10455
rect 3157 10217 3191 10251
rect 5089 10217 5123 10251
rect 7389 10217 7423 10251
rect 11989 10217 12023 10251
rect 14841 10217 14875 10251
rect 15853 10217 15887 10251
rect 16313 10217 16347 10251
rect 16497 10217 16531 10251
rect 17233 10217 17267 10251
rect 29285 10217 29319 10251
rect 5365 10149 5399 10183
rect 8502 10149 8536 10183
rect 16773 10149 16807 10183
rect 16865 10149 16899 10183
rect 16983 10149 17017 10183
rect 17385 10149 17419 10183
rect 17601 10149 17635 10183
rect 26157 10149 26191 10183
rect 26591 10149 26625 10183
rect 27077 10149 27111 10183
rect 28917 10149 28951 10183
rect 29009 10149 29043 10183
rect 30490 10149 30524 10183
rect 2145 10081 2179 10115
rect 2605 10081 2639 10115
rect 2697 10081 2731 10115
rect 2881 10081 2915 10115
rect 3893 10081 3927 10115
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 5641 10081 5675 10115
rect 6009 10081 6043 10115
rect 6101 10081 6135 10115
rect 6377 10081 6411 10115
rect 8769 10081 8803 10115
rect 9137 10081 9171 10115
rect 9229 10081 9263 10115
rect 9321 10081 9355 10115
rect 9505 10081 9539 10115
rect 10425 10081 10459 10115
rect 10517 10081 10551 10115
rect 10609 10081 10643 10115
rect 10793 10081 10827 10115
rect 11345 10081 11379 10115
rect 11529 10081 11563 10115
rect 11621 10081 11655 10115
rect 11713 10081 11747 10115
rect 13185 10081 13219 10115
rect 13452 10081 13486 10115
rect 14933 10081 14967 10115
rect 15025 10081 15059 10115
rect 15209 10081 15243 10115
rect 15669 10081 15703 10115
rect 15945 10081 15979 10115
rect 16221 10081 16255 10115
rect 16681 10081 16715 10115
rect 17141 10081 17175 10115
rect 19717 10081 19751 10115
rect 19984 10081 20018 10115
rect 22385 10081 22419 10115
rect 23673 10081 23707 10115
rect 23940 10081 23974 10115
rect 26709 10081 26743 10115
rect 26801 10081 26835 10115
rect 26893 10081 26927 10115
rect 27307 10081 27341 10115
rect 27445 10081 27479 10115
rect 27537 10081 27571 10115
rect 27629 10081 27663 10115
rect 28089 10081 28123 10115
rect 28273 10081 28307 10115
rect 28779 10081 28813 10115
rect 29101 10081 29135 10115
rect 30757 10081 30791 10115
rect 2237 10013 2271 10047
rect 3709 10013 3743 10047
rect 4445 10013 4479 10047
rect 21833 10013 21867 10047
rect 22201 10013 22235 10047
rect 26433 10013 26467 10047
rect 27169 10013 27203 10047
rect 28641 10013 28675 10047
rect 15301 9945 15335 9979
rect 15485 9945 15519 9979
rect 21281 9945 21315 9979
rect 27813 9945 27847 9979
rect 1869 9877 1903 9911
rect 2881 9877 2915 9911
rect 4721 9877 4755 9911
rect 5825 9877 5859 9911
rect 6285 9877 6319 9911
rect 8861 9877 8895 9911
rect 10149 9877 10183 9911
rect 14565 9877 14599 9911
rect 17417 9877 17451 9911
rect 21097 9877 21131 9911
rect 22569 9877 22603 9911
rect 25053 9877 25087 9911
rect 26065 9877 26099 9911
rect 27905 9877 27939 9911
rect 29377 9877 29411 9911
rect 3065 9673 3099 9707
rect 4261 9673 4295 9707
rect 4537 9673 4571 9707
rect 5457 9673 5491 9707
rect 6285 9673 6319 9707
rect 13645 9673 13679 9707
rect 14657 9673 14691 9707
rect 14933 9673 14967 9707
rect 20085 9673 20119 9707
rect 26433 9673 26467 9707
rect 30021 9673 30055 9707
rect 4445 9605 4479 9639
rect 5181 9605 5215 9639
rect 6745 9605 6779 9639
rect 11529 9605 11563 9639
rect 12265 9605 12299 9639
rect 12449 9605 12483 9639
rect 14749 9605 14783 9639
rect 16497 9605 16531 9639
rect 3801 9537 3835 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 16313 9537 16347 9571
rect 27813 9537 27847 9571
rect 28457 9537 28491 9571
rect 1317 9469 1351 9503
rect 1409 9469 1443 9503
rect 1501 9469 1535 9503
rect 1685 9469 1719 9503
rect 1952 9469 1986 9503
rect 3985 9469 4019 9503
rect 4169 9469 4203 9503
rect 4261 9469 4295 9503
rect 4721 9469 4755 9503
rect 4905 9469 4939 9503
rect 4997 9469 5031 9503
rect 5089 9469 5123 9503
rect 5549 9469 5583 9503
rect 5825 9469 5859 9503
rect 6009 9469 6043 9503
rect 6193 9469 6227 9503
rect 6469 9469 6503 9503
rect 6561 9469 6595 9503
rect 6837 9469 6871 9503
rect 7113 9469 7147 9503
rect 7573 9469 7607 9503
rect 7757 9469 7791 9503
rect 7849 9469 7883 9503
rect 7941 9469 7975 9503
rect 8401 9469 8435 9503
rect 10057 9469 10091 9503
rect 11805 9469 11839 9503
rect 12081 9469 12115 9503
rect 12357 9469 12391 9503
rect 12633 9469 12667 9503
rect 12725 9469 12759 9503
rect 13829 9469 13863 9503
rect 14013 9469 14047 9503
rect 14105 9469 14139 9503
rect 14289 9469 14323 9503
rect 14473 9469 14507 9503
rect 16037 9469 16071 9503
rect 16129 9469 16163 9503
rect 16405 9469 16439 9503
rect 19257 9469 19291 9503
rect 19441 9469 19475 9503
rect 20269 9469 20303 9503
rect 20361 9469 20395 9503
rect 20453 9469 20487 9503
rect 20729 9469 20763 9503
rect 22017 9469 22051 9503
rect 22109 9469 22143 9503
rect 22293 9469 22327 9503
rect 22560 9469 22594 9503
rect 23857 9469 23891 9503
rect 25881 9469 25915 9503
rect 27557 9469 27591 9503
rect 28089 9469 28123 9503
rect 28273 9469 28307 9503
rect 28549 9469 28583 9503
rect 28825 9469 28859 9503
rect 29561 9469 29595 9503
rect 29929 9469 29963 9503
rect 3249 9401 3283 9435
rect 5917 9401 5951 9435
rect 7297 9401 7331 9435
rect 7481 9401 7515 9435
rect 8668 9401 8702 9435
rect 10394 9401 10428 9435
rect 15117 9401 15151 9435
rect 20571 9401 20605 9435
rect 24124 9401 24158 9435
rect 1225 9333 1259 9367
rect 5641 9333 5675 9367
rect 8217 9333 8251 9367
rect 9781 9333 9815 9367
rect 11713 9333 11747 9367
rect 11897 9333 11931 9367
rect 14907 9333 14941 9367
rect 19533 9333 19567 9367
rect 23673 9333 23707 9367
rect 25237 9333 25271 9367
rect 25329 9333 25363 9367
rect 27905 9333 27939 9367
rect 28733 9333 28767 9367
rect 29469 9333 29503 9367
rect 6193 9129 6227 9163
rect 9045 9129 9079 9163
rect 9505 9129 9539 9163
rect 13001 9129 13035 9163
rect 13169 9129 13203 9163
rect 16957 9129 16991 9163
rect 22293 9129 22327 9163
rect 9137 9061 9171 9095
rect 11796 9061 11830 9095
rect 13369 9061 13403 9095
rect 22109 9061 22143 9095
rect 23831 9061 23865 9095
rect 23949 9061 23983 9095
rect 27660 9061 27694 9095
rect 29193 9061 29227 9095
rect 29530 9061 29564 9095
rect 1961 8993 1995 9027
rect 2228 8993 2262 9027
rect 3617 8993 3651 9027
rect 6009 8993 6043 9027
rect 6101 8993 6135 9027
rect 7389 8993 7423 9027
rect 7932 8993 7966 9027
rect 9321 8993 9355 9027
rect 11529 8993 11563 9027
rect 15025 8993 15059 9027
rect 15577 8993 15611 9027
rect 17141 8993 17175 9027
rect 17325 8993 17359 9027
rect 18521 8993 18555 9027
rect 19165 8993 19199 9027
rect 20085 8993 20119 9027
rect 21005 8993 21039 9027
rect 21281 8993 21315 9027
rect 22477 8993 22511 9027
rect 22569 8993 22603 9027
rect 22661 8993 22695 9027
rect 22799 8993 22833 9027
rect 24041 8993 24075 9027
rect 24133 8993 24167 9027
rect 24593 8993 24627 9027
rect 27905 8993 27939 9027
rect 29009 8993 29043 9027
rect 29285 8993 29319 9027
rect 3525 8925 3559 8959
rect 4261 8925 4295 8959
rect 4997 8925 5031 8959
rect 5549 8925 5583 8959
rect 7481 8925 7515 8959
rect 7665 8925 7699 8959
rect 15209 8925 15243 8959
rect 18337 8925 18371 8959
rect 19073 8925 19107 8959
rect 19901 8925 19935 8959
rect 22937 8925 22971 8959
rect 23673 8925 23707 8959
rect 24317 8925 24351 8959
rect 28825 8925 28859 8959
rect 3985 8857 4019 8891
rect 12909 8857 12943 8891
rect 15393 8857 15427 8891
rect 26525 8857 26559 8891
rect 3341 8789 3375 8823
rect 4813 8789 4847 8823
rect 5917 8789 5951 8823
rect 13185 8789 13219 8823
rect 14841 8789 14875 8823
rect 18705 8789 18739 8823
rect 18797 8789 18831 8823
rect 19165 8789 19199 8823
rect 20269 8789 20303 8823
rect 24501 8789 24535 8823
rect 30665 8789 30699 8823
rect 2605 8585 2639 8619
rect 3249 8585 3283 8619
rect 3433 8585 3467 8619
rect 8585 8585 8619 8619
rect 13645 8585 13679 8619
rect 20085 8585 20119 8619
rect 25605 8585 25639 8619
rect 25973 8585 26007 8619
rect 29653 8585 29687 8619
rect 4353 8517 4387 8551
rect 4077 8449 4111 8483
rect 5825 8449 5859 8483
rect 16313 8449 16347 8483
rect 28365 8449 28399 8483
rect 28733 8449 28767 8483
rect 2605 8381 2639 8415
rect 2789 8381 2823 8415
rect 2881 8381 2915 8415
rect 3985 8381 4019 8415
rect 5558 8381 5592 8415
rect 6469 8381 6503 8415
rect 8677 8381 8711 8415
rect 13553 8381 13587 8415
rect 14473 8381 14507 8415
rect 14565 8381 14599 8415
rect 14749 8381 14783 8415
rect 15005 8381 15039 8415
rect 16497 8381 16531 8415
rect 16773 8381 16807 8415
rect 18337 8381 18371 8415
rect 18429 8381 18463 8415
rect 18705 8381 18739 8415
rect 18961 8381 18995 8415
rect 20361 8381 20395 8415
rect 20453 8381 20487 8415
rect 20637 8381 20671 8415
rect 20904 8381 20938 8415
rect 22293 8381 22327 8415
rect 22569 8381 22603 8415
rect 22661 8381 22695 8415
rect 22753 8381 22787 8415
rect 22937 8381 22971 8415
rect 23213 8381 23247 8415
rect 23397 8381 23431 8415
rect 23673 8381 23707 8415
rect 25789 8381 25823 8415
rect 25881 8381 25915 8415
rect 26525 8381 26559 8415
rect 27629 8381 27663 8415
rect 28089 8381 28123 8415
rect 28549 8381 28583 8415
rect 29009 8381 29043 8415
rect 29469 8381 29503 8415
rect 3417 8313 3451 8347
rect 3617 8313 3651 8347
rect 5917 8313 5951 8347
rect 16681 8313 16715 8347
rect 17018 8313 17052 8347
rect 22431 8313 22465 8347
rect 26065 8313 26099 8347
rect 27261 8313 27295 8347
rect 29167 8313 29201 8347
rect 29285 8313 29319 8347
rect 29377 8313 29411 8347
rect 2973 8245 3007 8279
rect 4445 8245 4479 8279
rect 16129 8245 16163 8279
rect 18153 8245 18187 8279
rect 22017 8245 22051 8279
rect 23029 8245 23063 8279
rect 23581 8245 23615 8279
rect 28181 8245 28215 8279
rect 4997 8041 5031 8075
rect 15209 8041 15243 8075
rect 16405 8041 16439 8075
rect 16957 8041 16991 8075
rect 18705 8041 18739 8075
rect 20361 8041 20395 8075
rect 24317 8041 24351 8075
rect 28641 8041 28675 8075
rect 3884 7973 3918 8007
rect 12233 7973 12267 8007
rect 12449 7973 12483 8007
rect 14657 7973 14691 8007
rect 14749 7973 14783 8007
rect 14887 7973 14921 8007
rect 15485 7973 15519 8007
rect 16497 7973 16531 8007
rect 17509 7973 17543 8007
rect 17627 7973 17661 8007
rect 18153 7973 18187 8007
rect 18337 7973 18371 8007
rect 18981 7973 19015 8007
rect 19073 7973 19107 8007
rect 20729 7973 20763 8007
rect 20847 7973 20881 8007
rect 22845 7973 22879 8007
rect 26433 7973 26467 8007
rect 28135 7973 28169 8007
rect 28273 7973 28307 8007
rect 28365 7973 28399 8007
rect 28978 7973 29012 8007
rect 30573 7973 30607 8007
rect 30711 7973 30745 8007
rect 3617 7905 3651 7939
rect 7757 7905 7791 7939
rect 8033 7905 8067 7939
rect 9873 7905 9907 7939
rect 10057 7905 10091 7939
rect 10609 7905 10643 7939
rect 11253 7905 11287 7939
rect 11805 7905 11839 7939
rect 12633 7905 12667 7939
rect 13369 7905 13403 7939
rect 13645 7905 13679 7939
rect 14105 7905 14139 7939
rect 14381 7905 14415 7939
rect 14565 7905 14599 7939
rect 15025 7905 15059 7939
rect 15393 7905 15427 7939
rect 15577 7905 15611 7939
rect 15695 7905 15729 7939
rect 15853 7905 15887 7939
rect 17049 7905 17083 7939
rect 17325 7905 17359 7939
rect 17417 7905 17451 7939
rect 17785 7905 17819 7939
rect 17877 7905 17911 7939
rect 18889 7905 18923 7939
rect 19191 7905 19225 7939
rect 20545 7905 20579 7939
rect 20637 7905 20671 7939
rect 21005 7905 21039 7939
rect 21465 7905 21499 7939
rect 21741 7905 21775 7939
rect 22017 7905 22051 7939
rect 22569 7905 22603 7939
rect 22661 7905 22695 7939
rect 22937 7905 22971 7939
rect 23193 7905 23227 7939
rect 26249 7905 26283 7939
rect 27169 7905 27203 7939
rect 28457 7905 28491 7939
rect 28733 7905 28767 7939
rect 30389 7905 30423 7939
rect 30481 7905 30515 7939
rect 30849 7905 30883 7939
rect 7941 7837 7975 7871
rect 11529 7837 11563 7871
rect 11989 7837 12023 7871
rect 14289 7837 14323 7871
rect 17141 7837 17175 7871
rect 19349 7837 19383 7871
rect 21557 7837 21591 7871
rect 27997 7837 28031 7871
rect 9873 7769 9907 7803
rect 12081 7769 12115 7803
rect 22109 7769 22143 7803
rect 30205 7769 30239 7803
rect 7573 7701 7607 7735
rect 8125 7701 8159 7735
rect 10701 7701 10735 7735
rect 11069 7701 11103 7735
rect 11437 7701 11471 7735
rect 11621 7701 11655 7735
rect 12265 7701 12299 7735
rect 13461 7701 13495 7735
rect 13737 7701 13771 7735
rect 13921 7701 13955 7735
rect 18153 7701 18187 7735
rect 21649 7701 21683 7735
rect 21925 7701 21959 7735
rect 22385 7701 22419 7735
rect 22569 7701 22603 7735
rect 30113 7701 30147 7735
rect 8401 7497 8435 7531
rect 10425 7497 10459 7531
rect 12173 7497 12207 7531
rect 15117 7497 15151 7531
rect 17693 7497 17727 7531
rect 18889 7497 18923 7531
rect 28825 7497 28859 7531
rect 8217 7429 8251 7463
rect 11989 7429 12023 7463
rect 18705 7429 18739 7463
rect 26525 7429 26559 7463
rect 9045 7361 9079 7395
rect 9873 7361 9907 7395
rect 10609 7361 10643 7395
rect 13185 7361 13219 7395
rect 13737 7361 13771 7395
rect 17509 7361 17543 7395
rect 19073 7361 19107 7395
rect 20453 7361 20487 7395
rect 20729 7361 20763 7395
rect 24317 7361 24351 7395
rect 24777 7361 24811 7395
rect 28273 7361 28307 7395
rect 29009 7361 29043 7395
rect 6561 7293 6595 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 7104 7293 7138 7327
rect 8585 7293 8619 7327
rect 8677 7293 8711 7327
rect 9321 7293 9355 7327
rect 9965 7293 9999 7327
rect 10241 7293 10275 7327
rect 10517 7293 10551 7327
rect 10876 7293 10910 7327
rect 12449 7293 12483 7327
rect 14004 7293 14038 7327
rect 15393 7293 15427 7327
rect 15577 7293 15611 7327
rect 15715 7293 15749 7327
rect 15853 7293 15887 7327
rect 17417 7293 17451 7327
rect 17693 7293 17727 7327
rect 18889 7293 18923 7327
rect 20361 7293 20395 7327
rect 20821 7293 20855 7327
rect 24685 7293 24719 7327
rect 25145 7293 25179 7327
rect 25973 7293 26007 7327
rect 26157 7293 26191 7327
rect 27169 7293 27203 7327
rect 28181 7293 28215 7327
rect 28457 7293 28491 7327
rect 28641 7293 28675 7327
rect 29265 7293 29299 7327
rect 8769 7225 8803 7259
rect 8907 7225 8941 7259
rect 12265 7225 12299 7259
rect 15209 7225 15243 7259
rect 15485 7225 15519 7259
rect 19165 7225 19199 7259
rect 26249 7225 26283 7259
rect 26985 7225 27019 7259
rect 9137 7157 9171 7191
rect 10057 7157 10091 7191
rect 17877 7157 17911 7191
rect 25053 7157 25087 7191
rect 25973 7157 26007 7191
rect 26709 7157 26743 7191
rect 26801 7157 26835 7191
rect 30389 7157 30423 7191
rect 17785 6953 17819 6987
rect 20913 6953 20947 6987
rect 7021 6885 7055 6919
rect 9137 6885 9171 6919
rect 22017 6885 22051 6919
rect 23581 6885 23615 6919
rect 24317 6885 24351 6919
rect 26893 6885 26927 6919
rect 3617 6817 3651 6851
rect 3801 6817 3835 6851
rect 3893 6817 3927 6851
rect 4169 6817 4203 6851
rect 6285 6817 6319 6851
rect 8410 6817 8444 6851
rect 8677 6817 8711 6851
rect 8953 6817 8987 6851
rect 9045 6817 9079 6851
rect 9255 6817 9289 6851
rect 10425 6817 10459 6851
rect 10609 6817 10643 6851
rect 10977 6817 11011 6851
rect 11233 6817 11267 6851
rect 12541 6817 12575 6851
rect 12725 6817 12759 6851
rect 12817 6817 12851 6851
rect 13093 6817 13127 6851
rect 13185 6817 13219 6851
rect 13461 6817 13495 6851
rect 13717 6817 13751 6851
rect 15577 6817 15611 6851
rect 18061 6817 18095 6851
rect 19073 6817 19107 6851
rect 19257 6817 19291 6851
rect 19349 6817 19383 6851
rect 21097 6817 21131 6851
rect 21281 6817 21315 6851
rect 22477 6817 22511 6851
rect 22753 6817 22787 6851
rect 23213 6817 23247 6851
rect 23305 6817 23339 6851
rect 23489 6817 23523 6851
rect 23949 6817 23983 6851
rect 24041 6817 24075 6851
rect 24134 6817 24168 6851
rect 24409 6817 24443 6851
rect 24547 6817 24581 6851
rect 24961 6817 24995 6851
rect 25053 6817 25087 6851
rect 25237 6817 25271 6851
rect 25329 6817 25363 6851
rect 29101 6817 29135 6851
rect 29561 6817 29595 6851
rect 29654 6817 29688 6851
rect 29837 6817 29871 6851
rect 29929 6817 29963 6851
rect 30067 6817 30101 6851
rect 30481 6817 30515 6851
rect 30665 6817 30699 6851
rect 4353 6749 4387 6783
rect 4905 6749 4939 6783
rect 9413 6749 9447 6783
rect 13369 6749 13403 6783
rect 15485 6749 15519 6783
rect 17509 6749 17543 6783
rect 18153 6749 18187 6783
rect 18797 6749 18831 6783
rect 19441 6749 19475 6783
rect 22661 6749 22695 6783
rect 23765 6749 23799 6783
rect 25789 6749 25823 6783
rect 26985 6749 27019 6783
rect 29193 6749 29227 6783
rect 29469 6749 29503 6783
rect 30297 6749 30331 6783
rect 7297 6681 7331 6715
rect 14841 6681 14875 6715
rect 18521 6681 18555 6715
rect 19717 6681 19751 6715
rect 19901 6681 19935 6715
rect 22937 6681 22971 6715
rect 24685 6681 24719 6715
rect 26065 6681 26099 6715
rect 26617 6681 26651 6715
rect 27353 6681 27387 6715
rect 30205 6681 30239 6715
rect 3617 6613 3651 6647
rect 4077 6613 4111 6647
rect 8769 6613 8803 6647
rect 10793 6613 10827 6647
rect 12357 6613 12391 6647
rect 15945 6613 15979 6647
rect 18981 6613 19015 6647
rect 22477 6613 22511 6647
rect 23029 6613 23063 6647
rect 23489 6613 23523 6647
rect 23765 6613 23799 6647
rect 23857 6613 23891 6647
rect 25513 6613 25547 6647
rect 26249 6613 26283 6647
rect 26433 6613 26467 6647
rect 27445 6613 27479 6647
rect 8217 6409 8251 6443
rect 11529 6409 11563 6443
rect 11713 6409 11747 6443
rect 19441 6409 19475 6443
rect 20545 6409 20579 6443
rect 22109 6409 22143 6443
rect 22385 6409 22419 6443
rect 22569 6409 22603 6443
rect 22937 6409 22971 6443
rect 26157 6409 26191 6443
rect 26617 6409 26651 6443
rect 26893 6409 26927 6443
rect 29653 6409 29687 6443
rect 29837 6409 29871 6443
rect 30113 6409 30147 6443
rect 18429 6341 18463 6375
rect 23029 6341 23063 6375
rect 23949 6341 23983 6375
rect 9873 6273 9907 6307
rect 10057 6273 10091 6307
rect 13553 6273 13587 6307
rect 16221 6273 16255 6307
rect 16497 6273 16531 6307
rect 17233 6273 17267 6307
rect 17509 6273 17543 6307
rect 22753 6273 22787 6307
rect 26525 6273 26559 6307
rect 3249 6205 3283 6239
rect 3341 6205 3375 6239
rect 3525 6205 3559 6239
rect 3781 6205 3815 6239
rect 7297 6205 7331 6239
rect 7941 6205 7975 6239
rect 8033 6205 8067 6239
rect 9965 6205 9999 6239
rect 12173 6205 12207 6239
rect 13369 6205 13403 6239
rect 13737 6205 13771 6239
rect 16129 6205 16163 6239
rect 17141 6205 17175 6239
rect 17877 6205 17911 6239
rect 18245 6205 18279 6239
rect 18694 6205 18728 6239
rect 18798 6205 18832 6239
rect 19170 6205 19204 6239
rect 19625 6205 19659 6239
rect 19717 6205 19751 6239
rect 19901 6205 19935 6239
rect 19993 6205 20027 6239
rect 20269 6205 20303 6239
rect 20361 6205 20395 6239
rect 20637 6205 20671 6239
rect 22017 6205 22051 6239
rect 22109 6205 22143 6239
rect 22569 6205 22603 6239
rect 24041 6205 24075 6239
rect 26341 6205 26375 6239
rect 26893 6205 26927 6239
rect 27077 6205 27111 6239
rect 29285 6205 29319 6239
rect 29469 6205 29503 6239
rect 29745 6205 29779 6239
rect 29929 6205 29963 6239
rect 30021 6205 30055 6239
rect 30205 6205 30239 6239
rect 6377 6137 6411 6171
rect 7113 6137 7147 6171
rect 9606 6137 9640 6171
rect 11697 6137 11731 6171
rect 11897 6137 11931 6171
rect 12633 6137 12667 6171
rect 18061 6137 18095 6171
rect 18153 6137 18187 6171
rect 18981 6137 19015 6171
rect 19073 6137 19107 6171
rect 21833 6137 21867 6171
rect 22845 6137 22879 6171
rect 23397 6137 23431 6171
rect 26617 6137 26651 6171
rect 4905 6069 4939 6103
rect 8493 6069 8527 6103
rect 12265 6069 12299 6103
rect 13921 6069 13955 6103
rect 19349 6069 19383 6103
rect 20085 6069 20119 6103
rect 22293 6069 22327 6103
rect 26709 6069 26743 6103
rect 2697 5865 2731 5899
rect 8217 5865 8251 5899
rect 21373 5865 21407 5899
rect 21925 5865 21959 5899
rect 23857 5865 23891 5899
rect 6713 5797 6747 5831
rect 6929 5797 6963 5831
rect 8861 5797 8895 5831
rect 21833 5797 21867 5831
rect 22385 5797 22419 5831
rect 24317 5797 24351 5831
rect 28917 5797 28951 5831
rect 29377 5797 29411 5831
rect 2881 5729 2915 5763
rect 2973 5729 3007 5763
rect 3341 5729 3375 5763
rect 3709 5729 3743 5763
rect 3965 5729 3999 5763
rect 5365 5729 5399 5763
rect 7941 5729 7975 5763
rect 8033 5729 8067 5763
rect 8493 5729 8527 5763
rect 8677 5729 8711 5763
rect 8769 5729 8803 5763
rect 8979 5729 9013 5763
rect 9137 5729 9171 5763
rect 9413 5729 9447 5763
rect 9505 5729 9539 5763
rect 9597 5729 9631 5763
rect 9715 5729 9749 5763
rect 9873 5729 9907 5763
rect 11161 5729 11195 5763
rect 11345 5729 11379 5763
rect 12909 5729 12943 5763
rect 13277 5729 13311 5763
rect 13737 5729 13771 5763
rect 18889 5729 18923 5763
rect 19257 5729 19291 5763
rect 19441 5729 19475 5763
rect 19533 5729 19567 5763
rect 19717 5729 19751 5763
rect 21557 5729 21591 5763
rect 22109 5729 22143 5763
rect 22477 5729 22511 5763
rect 22661 5729 22695 5763
rect 23305 5729 23339 5763
rect 23489 5729 23523 5763
rect 23581 5729 23615 5763
rect 24041 5729 24075 5763
rect 24409 5729 24443 5763
rect 24593 5729 24627 5763
rect 25421 5729 25455 5763
rect 25513 5729 25547 5763
rect 28089 5729 28123 5763
rect 28273 5729 28307 5763
rect 29193 5729 29227 5763
rect 2697 5661 2731 5695
rect 3157 5661 3191 5695
rect 3249 5661 3283 5695
rect 3433 5661 3467 5695
rect 5641 5661 5675 5695
rect 5825 5661 5859 5695
rect 6377 5661 6411 5695
rect 13461 5661 13495 5695
rect 19073 5661 19107 5695
rect 19165 5661 19199 5695
rect 21741 5661 21775 5695
rect 22293 5661 22327 5695
rect 22937 5661 22971 5695
rect 24225 5661 24259 5695
rect 5181 5593 5215 5627
rect 13645 5593 13679 5627
rect 19717 5593 19751 5627
rect 28549 5593 28583 5627
rect 3617 5525 3651 5559
rect 5089 5525 5123 5559
rect 5549 5525 5583 5559
rect 6561 5525 6595 5559
rect 6745 5525 6779 5559
rect 9229 5525 9263 5559
rect 11529 5525 11563 5559
rect 13093 5525 13127 5559
rect 18705 5525 18739 5559
rect 21557 5525 21591 5559
rect 22109 5525 22143 5559
rect 22753 5525 22787 5559
rect 22845 5525 22879 5559
rect 23213 5525 23247 5559
rect 23305 5525 23339 5559
rect 23765 5525 23799 5559
rect 24041 5525 24075 5559
rect 24409 5525 24443 5559
rect 28457 5525 28491 5559
rect 28917 5525 28951 5559
rect 29101 5525 29135 5559
rect 29561 5525 29595 5559
rect 11621 5321 11655 5355
rect 12173 5321 12207 5355
rect 12550 5321 12584 5355
rect 13277 5321 13311 5355
rect 13921 5321 13955 5355
rect 14289 5321 14323 5355
rect 21465 5321 21499 5355
rect 22569 5321 22603 5355
rect 23397 5321 23431 5355
rect 24593 5321 24627 5355
rect 24869 5321 24903 5355
rect 28181 5321 28215 5355
rect 28641 5321 28675 5355
rect 12357 5253 12391 5287
rect 14105 5253 14139 5287
rect 21281 5253 21315 5287
rect 21833 5253 21867 5287
rect 22017 5253 22051 5287
rect 23489 5253 23523 5287
rect 23673 5253 23707 5287
rect 24133 5253 24167 5287
rect 25145 5253 25179 5287
rect 25329 5253 25363 5287
rect 25881 5253 25915 5287
rect 28273 5253 28307 5287
rect 28825 5253 28859 5287
rect 29101 5253 29135 5287
rect 4905 5185 4939 5219
rect 5549 5185 5583 5219
rect 5825 5185 5859 5219
rect 6745 5185 6779 5219
rect 9321 5185 9355 5219
rect 11713 5185 11747 5219
rect 13369 5185 13403 5219
rect 15853 5185 15887 5219
rect 21005 5185 21039 5219
rect 23305 5185 23339 5219
rect 24225 5185 24259 5219
rect 24317 5185 24351 5219
rect 24961 5185 24995 5219
rect 25697 5185 25731 5219
rect 26157 5185 26191 5219
rect 1409 5117 1443 5151
rect 1501 5117 1535 5151
rect 1685 5117 1719 5151
rect 3433 5117 3467 5151
rect 3700 5117 3734 5151
rect 5089 5117 5123 5151
rect 5942 5117 5976 5151
rect 6101 5117 6135 5151
rect 8125 5117 8159 5151
rect 8401 5117 8435 5151
rect 8861 5117 8895 5151
rect 9137 5117 9171 5151
rect 11161 5117 11195 5151
rect 11437 5117 11471 5151
rect 11989 5117 12023 5151
rect 12265 5117 12299 5151
rect 13093 5117 13127 5151
rect 13737 5117 13771 5151
rect 14013 5117 14047 5151
rect 15945 5117 15979 5151
rect 18705 5117 18739 5151
rect 18797 5117 18831 5151
rect 22753 5117 22787 5151
rect 22845 5117 22879 5151
rect 23857 5117 23891 5151
rect 24041 5117 24075 5151
rect 25053 5117 25087 5151
rect 27813 5117 27847 5151
rect 27997 5117 28031 5151
rect 30214 5117 30248 5151
rect 30481 5117 30515 5151
rect 30665 5117 30699 5151
rect 30757 5117 30791 5151
rect 30849 5117 30883 5151
rect 1952 5049 1986 5083
rect 8493 5049 8527 5083
rect 12725 5049 12759 5083
rect 14473 5049 14507 5083
rect 21557 5049 21591 5083
rect 23121 5049 23155 5083
rect 23213 5049 23247 5083
rect 23673 5049 23707 5083
rect 25605 5049 25639 5083
rect 3065 4981 3099 5015
rect 4813 4981 4847 5015
rect 8033 4981 8067 5015
rect 8585 4981 8619 5015
rect 8953 4981 8987 5015
rect 11069 4981 11103 5015
rect 11253 4981 11287 5015
rect 11805 4981 11839 5015
rect 12515 4981 12549 5015
rect 12909 4981 12943 5015
rect 13553 4981 13587 5015
rect 14273 4981 14307 5015
rect 16313 4981 16347 5015
rect 24685 4981 24719 5015
rect 28641 4981 28675 5015
rect 30941 4981 30975 5015
rect 1869 4777 1903 4811
rect 2145 4777 2179 4811
rect 3893 4777 3927 4811
rect 4077 4777 4111 4811
rect 9229 4777 9263 4811
rect 12449 4777 12483 4811
rect 14381 4777 14415 4811
rect 18245 4777 18279 4811
rect 18521 4777 18555 4811
rect 22569 4777 22603 4811
rect 23213 4777 23247 4811
rect 23397 4777 23431 4811
rect 24317 4777 24351 4811
rect 26433 4777 26467 4811
rect 27153 4777 27187 4811
rect 28089 4777 28123 4811
rect 28825 4777 28859 4811
rect 2329 4709 2363 4743
rect 3157 4709 3191 4743
rect 4689 4709 4723 4743
rect 4905 4709 4939 4743
rect 8116 4709 8150 4743
rect 11244 4709 11278 4743
rect 12601 4709 12635 4743
rect 12817 4709 12851 4743
rect 14533 4709 14567 4743
rect 14749 4709 14783 4743
rect 18981 4709 19015 4743
rect 19533 4709 19567 4743
rect 23857 4709 23891 4743
rect 24041 4709 24075 4743
rect 25513 4709 25547 4743
rect 27353 4709 27387 4743
rect 27997 4709 28031 4743
rect 28257 4709 28291 4743
rect 28457 4709 28491 4743
rect 29938 4709 29972 4743
rect 1777 4641 1811 4675
rect 1961 4641 1995 4675
rect 2053 4641 2087 4675
rect 2605 4641 2639 4675
rect 2881 4641 2915 4675
rect 3065 4641 3099 4675
rect 3801 4641 3835 4675
rect 5181 4641 5215 4675
rect 7849 4641 7883 4675
rect 10977 4641 11011 4675
rect 12909 4641 12943 4675
rect 13165 4641 13199 4675
rect 14933 4641 14967 4675
rect 15117 4641 15151 4675
rect 16129 4641 16163 4675
rect 16221 4641 16255 4675
rect 16405 4641 16439 4675
rect 16497 4641 16531 4675
rect 16681 4641 16715 4675
rect 17325 4641 17359 4675
rect 17509 4641 17543 4675
rect 17693 4641 17727 4675
rect 17877 4641 17911 4675
rect 19165 4641 19199 4675
rect 19258 4641 19292 4675
rect 19441 4641 19475 4675
rect 19671 4641 19705 4675
rect 19993 4641 20027 4675
rect 20085 4641 20119 4675
rect 22661 4641 22695 4675
rect 22845 4641 22879 4675
rect 22937 4641 22971 4675
rect 23029 4641 23063 4675
rect 23581 4641 23615 4675
rect 23949 4641 23983 4675
rect 24133 4641 24167 4675
rect 24685 4641 24719 4675
rect 25237 4641 25271 4675
rect 26893 4641 26927 4675
rect 27813 4641 27847 4675
rect 30205 4641 30239 4675
rect 2329 4573 2363 4607
rect 4445 4573 4479 4607
rect 17601 4573 17635 4607
rect 18061 4573 18095 4607
rect 18429 4573 18463 4607
rect 22109 4573 22143 4607
rect 23765 4573 23799 4607
rect 24593 4573 24627 4607
rect 25329 4573 25363 4607
rect 25605 4573 25639 4607
rect 26065 4573 26099 4607
rect 2513 4505 2547 4539
rect 12357 4505 12391 4539
rect 14289 4505 14323 4539
rect 18981 4505 19015 4539
rect 19809 4505 19843 4539
rect 22385 4505 22419 4539
rect 25053 4505 25087 4539
rect 25789 4505 25823 4539
rect 26617 4505 26651 4539
rect 2697 4437 2731 4471
rect 4077 4437 4111 4471
rect 4537 4437 4571 4471
rect 4721 4437 4755 4471
rect 5089 4437 5123 4471
rect 12633 4437 12667 4471
rect 14565 4437 14599 4471
rect 15025 4437 15059 4471
rect 16405 4437 16439 4471
rect 16681 4437 16715 4471
rect 23581 4437 23615 4471
rect 24685 4437 24719 4471
rect 25237 4437 25271 4471
rect 26985 4437 27019 4471
rect 27169 4437 27203 4471
rect 27629 4437 27663 4471
rect 28273 4437 28307 4471
rect 4169 4233 4203 4267
rect 9045 4233 9079 4267
rect 14933 4233 14967 4267
rect 18153 4233 18187 4267
rect 18337 4233 18371 4267
rect 19349 4233 19383 4267
rect 23949 4233 23983 4267
rect 28641 4233 28675 4267
rect 2697 4165 2731 4199
rect 2973 4165 3007 4199
rect 4537 4165 4571 4199
rect 7849 4165 7883 4199
rect 16681 4165 16715 4199
rect 23213 4165 23247 4199
rect 2789 4097 2823 4131
rect 5181 4097 5215 4131
rect 5641 4097 5675 4131
rect 5917 4097 5951 4131
rect 6193 4097 6227 4131
rect 9781 4097 9815 4131
rect 10333 4097 10367 4131
rect 10517 4097 10551 4131
rect 17325 4097 17359 4131
rect 17509 4097 17543 4131
rect 17969 4097 18003 4131
rect 22937 4097 22971 4131
rect 23397 4097 23431 4131
rect 2053 4029 2087 4063
rect 2145 4029 2179 4063
rect 2329 4029 2363 4063
rect 2421 4029 2455 4063
rect 3065 4029 3099 4063
rect 3249 4029 3283 4063
rect 3893 4029 3927 4063
rect 4997 4029 5031 4063
rect 6034 4029 6068 4063
rect 6837 4029 6871 4063
rect 8063 4029 8097 4063
rect 8217 4029 8251 4063
rect 8615 4029 8649 4063
rect 9137 4029 9171 4063
rect 9689 4029 9723 4063
rect 10425 4029 10459 4063
rect 13185 4029 13219 4063
rect 13277 4029 13311 4063
rect 13553 4029 13587 4063
rect 13820 4029 13854 4063
rect 15025 4029 15059 4063
rect 15117 4029 15151 4063
rect 15301 4029 15335 4063
rect 17876 4029 17910 4063
rect 18245 4029 18279 4063
rect 18429 4029 18463 4063
rect 18705 4029 18739 4063
rect 18798 4029 18832 4063
rect 19170 4029 19204 4063
rect 21925 4029 21959 4063
rect 24041 4029 24075 4063
rect 27261 4029 27295 4063
rect 27445 4029 27479 4063
rect 27629 4029 27663 4063
rect 28273 4029 28307 4063
rect 29009 4029 29043 4063
rect 2697 3961 2731 3995
rect 2789 3961 2823 3995
rect 10784 3961 10818 3995
rect 15568 3961 15602 3995
rect 17601 3961 17635 3995
rect 18981 3961 19015 3995
rect 19073 3961 19107 3995
rect 28641 3961 28675 3995
rect 29254 3961 29288 3995
rect 1961 3893 1995 3927
rect 2237 3893 2271 3927
rect 2513 3893 2547 3927
rect 3985 3893 4019 3927
rect 4169 3893 4203 3927
rect 8493 3893 8527 3927
rect 8677 3893 8711 3927
rect 9229 3893 9263 3927
rect 9597 3893 9631 3927
rect 11897 3893 11931 3927
rect 16773 3893 16807 3927
rect 21833 3893 21867 3927
rect 28825 3893 28859 3927
rect 30389 3893 30423 3927
rect 3157 3689 3191 3723
rect 3433 3689 3467 3723
rect 16129 3689 16163 3723
rect 18337 3689 18371 3723
rect 21833 3689 21867 3723
rect 25145 3689 25179 3723
rect 25237 3689 25271 3723
rect 25329 3689 25363 3723
rect 29193 3689 29227 3723
rect 2044 3621 2078 3655
rect 9965 3621 9999 3655
rect 17969 3621 18003 3655
rect 18153 3621 18187 3655
rect 22109 3621 22143 3655
rect 25605 3621 25639 3655
rect 25881 3621 25915 3655
rect 26769 3621 26803 3655
rect 26985 3621 27019 3655
rect 27997 3621 28031 3655
rect 28181 3621 28215 3655
rect 1777 3553 1811 3587
rect 3617 3553 3651 3587
rect 4077 3553 4111 3587
rect 4333 3553 4367 3587
rect 14105 3553 14139 3587
rect 14289 3553 14323 3587
rect 16313 3553 16347 3587
rect 16497 3553 16531 3587
rect 16589 3553 16623 3587
rect 18521 3553 18555 3587
rect 18613 3553 18647 3587
rect 21741 3553 21775 3587
rect 21925 3553 21959 3587
rect 22201 3553 22235 3587
rect 22293 3553 22327 3587
rect 22477 3553 22511 3587
rect 22661 3553 22695 3587
rect 22753 3553 22787 3587
rect 22937 3553 22971 3587
rect 25513 3553 25547 3587
rect 25789 3553 25823 3587
rect 25973 3553 26007 3587
rect 26157 3553 26191 3587
rect 29285 3553 29319 3587
rect 3801 3485 3835 3519
rect 9597 3417 9631 3451
rect 24961 3417 24995 3451
rect 5457 3349 5491 3383
rect 9965 3349 9999 3383
rect 10149 3349 10183 3383
rect 14289 3349 14323 3383
rect 21557 3349 21591 3383
rect 22661 3349 22695 3383
rect 22845 3349 22879 3383
rect 26617 3349 26651 3383
rect 26801 3349 26835 3383
rect 28365 3349 28399 3383
rect 4077 3145 4111 3179
rect 6009 3145 6043 3179
rect 9321 3145 9355 3179
rect 18797 3145 18831 3179
rect 22201 3145 22235 3179
rect 22293 3145 22327 3179
rect 26525 3145 26559 3179
rect 28365 3145 28399 3179
rect 30389 3145 30423 3179
rect 3065 3077 3099 3111
rect 7113 3077 7147 3111
rect 9229 3077 9263 3111
rect 10517 3077 10551 3111
rect 26709 3077 26743 3111
rect 4261 3009 4295 3043
rect 4445 3009 4479 3043
rect 4537 3009 4571 3043
rect 6285 3009 6319 3043
rect 9965 3009 9999 3043
rect 27997 3009 28031 3043
rect 1409 2941 1443 2975
rect 1501 2941 1535 2975
rect 1685 2941 1719 2975
rect 1952 2941 1986 2975
rect 3985 2941 4019 2975
rect 4353 2941 4387 2975
rect 5181 2941 5215 2975
rect 5365 2941 5399 2975
rect 6469 2941 6503 2975
rect 6561 2941 6595 2975
rect 6745 2941 6779 2975
rect 6929 2941 6963 2975
rect 7205 2941 7239 2975
rect 8953 2941 8987 2975
rect 9229 2941 9263 2975
rect 10124 2941 10158 2975
rect 10241 2941 10275 2975
rect 10977 2941 11011 2975
rect 11161 2941 11195 2975
rect 12817 2941 12851 2975
rect 13369 2941 13403 2975
rect 14105 2941 14139 2975
rect 14381 2941 14415 2975
rect 18705 2941 18739 2975
rect 20545 2941 20579 2975
rect 20637 2941 20671 2975
rect 20821 2941 20855 2975
rect 23673 2941 23707 2975
rect 23857 2941 23891 2975
rect 26985 2941 27019 2975
rect 27077 2941 27111 2975
rect 28641 2941 28675 2975
rect 28733 2941 28767 2975
rect 29009 2941 29043 2975
rect 26571 2907 26605 2941
rect 6193 2873 6227 2907
rect 6285 2873 6319 2907
rect 8493 2873 8527 2907
rect 12909 2873 12943 2907
rect 13093 2873 13127 2907
rect 21088 2873 21122 2907
rect 23406 2873 23440 2907
rect 26341 2873 26375 2907
rect 26801 2873 26835 2907
rect 27261 2873 27295 2907
rect 27445 2873 27479 2907
rect 28365 2873 28399 2907
rect 29254 2873 29288 2907
rect 3341 2805 3375 2839
rect 5273 2805 5307 2839
rect 5825 2805 5859 2839
rect 5993 2805 6027 2839
rect 6837 2805 6871 2839
rect 8585 2805 8619 2839
rect 9045 2805 9079 2839
rect 12817 2805 12851 2839
rect 13277 2805 13311 2839
rect 24041 2805 24075 2839
rect 27629 2805 27663 2839
rect 28549 2805 28583 2839
rect 3249 2601 3283 2635
rect 5917 2601 5951 2635
rect 7021 2601 7055 2635
rect 9137 2601 9171 2635
rect 10057 2601 10091 2635
rect 10977 2601 11011 2635
rect 12817 2601 12851 2635
rect 14289 2601 14323 2635
rect 18337 2601 18371 2635
rect 19533 2601 19567 2635
rect 21281 2601 21315 2635
rect 9965 2533 9999 2567
rect 12449 2533 12483 2567
rect 12649 2533 12683 2567
rect 13154 2533 13188 2567
rect 18245 2533 18279 2567
rect 23121 2533 23155 2567
rect 24317 2533 24351 2567
rect 24777 2533 24811 2567
rect 26065 2533 26099 2567
rect 27169 2533 27203 2567
rect 27813 2533 27847 2567
rect 3433 2465 3467 2499
rect 3525 2465 3559 2499
rect 5457 2465 5491 2499
rect 5641 2465 5675 2499
rect 6101 2465 6135 2499
rect 6377 2465 6411 2499
rect 9597 2465 9631 2499
rect 9689 2465 9723 2499
rect 9781 2465 9815 2499
rect 11253 2465 11287 2499
rect 11345 2465 11379 2499
rect 11437 2465 11471 2499
rect 12909 2465 12943 2499
rect 14565 2465 14599 2499
rect 15025 2465 15059 2499
rect 15577 2465 15611 2499
rect 16221 2465 16255 2499
rect 16773 2465 16807 2499
rect 16865 2465 16899 2499
rect 16957 2465 16991 2499
rect 17141 2465 17175 2499
rect 17233 2465 17267 2499
rect 17417 2465 17451 2499
rect 17693 2465 17727 2499
rect 17785 2465 17819 2499
rect 18061 2465 18095 2499
rect 18429 2465 18463 2499
rect 19349 2465 19383 2499
rect 19625 2465 19659 2499
rect 20913 2465 20947 2499
rect 21557 2465 21591 2499
rect 21649 2465 21683 2499
rect 21741 2465 21775 2499
rect 21925 2465 21959 2499
rect 22017 2465 22051 2499
rect 22569 2465 22603 2499
rect 22753 2465 22787 2499
rect 23673 2465 23707 2499
rect 23949 2465 23983 2499
rect 24133 2465 24167 2499
rect 24409 2465 24443 2499
rect 24685 2465 24719 2499
rect 24869 2465 24903 2499
rect 24961 2465 24995 2499
rect 25237 2465 25271 2499
rect 25881 2465 25915 2499
rect 26709 2465 26743 2499
rect 27629 2465 27663 2499
rect 3249 2397 3283 2431
rect 6285 2397 6319 2431
rect 7297 2397 7331 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 8334 2397 8368 2431
rect 8493 2397 8527 2431
rect 10609 2397 10643 2431
rect 11161 2397 11195 2431
rect 15669 2397 15703 2431
rect 17325 2397 17359 2431
rect 23489 2397 23523 2431
rect 23857 2397 23891 2431
rect 14473 2329 14507 2363
rect 17601 2329 17635 2363
rect 18613 2329 18647 2363
rect 21005 2329 21039 2363
rect 23305 2329 23339 2363
rect 24501 2329 24535 2363
rect 25329 2329 25363 2363
rect 26801 2329 26835 2363
rect 5457 2261 5491 2295
rect 9413 2261 9447 2295
rect 12633 2261 12667 2295
rect 15117 2261 15151 2295
rect 15853 2261 15887 2295
rect 16313 2261 16347 2295
rect 16497 2261 16531 2295
rect 17877 2261 17911 2295
rect 19165 2261 19199 2295
rect 23121 2261 23155 2295
rect 25053 2261 25087 2295
rect 25697 2261 25731 2295
rect 26617 2261 26651 2295
rect 27169 2261 27203 2295
rect 27353 2261 27387 2295
rect 27445 2261 27479 2295
rect 6285 2057 6319 2091
rect 8401 2057 8435 2091
rect 9965 2057 9999 2091
rect 11621 2057 11655 2091
rect 13553 2057 13587 2091
rect 16681 2057 16715 2091
rect 18521 2057 18555 2091
rect 25697 2057 25731 2091
rect 26157 2057 26191 2091
rect 27813 2057 27847 2091
rect 12633 1989 12667 2023
rect 14933 1989 14967 2023
rect 25329 1989 25363 2023
rect 25973 1989 26007 2023
rect 6929 1921 6963 1955
rect 8033 1921 8067 1955
rect 11713 1921 11747 1955
rect 11897 1921 11931 1955
rect 12725 1921 12759 1955
rect 14841 1921 14875 1955
rect 15301 1921 15335 1955
rect 16773 1921 16807 1955
rect 17141 1921 17175 1955
rect 19257 1921 19291 1955
rect 25237 1921 25271 1955
rect 26433 1921 26467 1955
rect 4537 1853 4571 1887
rect 4629 1853 4663 1887
rect 4721 1853 4755 1887
rect 4905 1853 4939 1887
rect 5172 1853 5206 1887
rect 9781 1853 9815 1887
rect 11078 1853 11112 1887
rect 11345 1853 11379 1887
rect 11437 1853 11471 1887
rect 11529 1853 11563 1887
rect 11989 1853 12023 1887
rect 12081 1853 12115 1887
rect 12357 1853 12391 1887
rect 12633 1853 12667 1887
rect 13737 1853 13771 1887
rect 14013 1853 14047 1887
rect 14657 1853 14691 1887
rect 15025 1853 15059 1887
rect 15117 1853 15151 1887
rect 16957 1853 16991 1887
rect 19717 1853 19751 1887
rect 19809 1853 19843 1887
rect 19901 1853 19935 1887
rect 20085 1853 20119 1887
rect 20361 1853 20395 1887
rect 20453 1853 20487 1887
rect 20637 1853 20671 1887
rect 20821 1853 20855 1887
rect 21373 1853 21407 1887
rect 22753 1853 22787 1887
rect 22845 1853 22879 1887
rect 23029 1853 23063 1887
rect 23121 1853 23155 1887
rect 23213 1853 23247 1887
rect 28089 1853 28123 1887
rect 6377 1785 6411 1819
rect 9514 1785 9548 1819
rect 14105 1785 14139 1819
rect 15568 1785 15602 1819
rect 17408 1785 17442 1819
rect 18705 1785 18739 1819
rect 20545 1785 20579 1819
rect 23489 1785 23523 1819
rect 24970 1785 25004 1819
rect 25697 1785 25731 1819
rect 26341 1785 26375 1819
rect 26700 1785 26734 1819
rect 4445 1717 4479 1751
rect 7389 1717 7423 1751
rect 12173 1717 12207 1751
rect 12449 1717 12483 1751
rect 13369 1717 13403 1751
rect 13921 1717 13955 1751
rect 19441 1717 19475 1751
rect 20269 1717 20303 1751
rect 22661 1717 22695 1751
rect 23857 1717 23891 1751
rect 25881 1717 25915 1751
rect 26141 1717 26175 1751
rect 27997 1717 28031 1751
rect 5641 1513 5675 1547
rect 7573 1513 7607 1547
rect 7941 1513 7975 1547
rect 8861 1513 8895 1547
rect 10701 1513 10735 1547
rect 12541 1513 12575 1547
rect 14013 1513 14047 1547
rect 15485 1513 15519 1547
rect 15577 1513 15611 1547
rect 17601 1513 17635 1547
rect 17693 1513 17727 1547
rect 19165 1513 19199 1547
rect 21005 1513 21039 1547
rect 23029 1513 23063 1547
rect 23213 1513 23247 1547
rect 24685 1513 24719 1547
rect 24869 1513 24903 1547
rect 26801 1513 26835 1547
rect 26985 1513 27019 1547
rect 28917 1513 28951 1547
rect 4528 1445 4562 1479
rect 6460 1445 6494 1479
rect 8033 1445 8067 1479
rect 8677 1445 8711 1479
rect 9566 1445 9600 1479
rect 12081 1445 12115 1479
rect 12900 1445 12934 1479
rect 14350 1445 14384 1479
rect 16488 1445 16522 1479
rect 19870 1445 19904 1479
rect 23550 1445 23584 1479
rect 25982 1445 26016 1479
rect 4261 1377 4295 1411
rect 6101 1377 6135 1411
rect 7849 1377 7883 1411
rect 9045 1377 9079 1411
rect 14105 1377 14139 1411
rect 15761 1377 15795 1411
rect 16221 1377 16255 1411
rect 17969 1377 18003 1411
rect 18061 1377 18095 1411
rect 18153 1377 18187 1411
rect 18337 1377 18371 1411
rect 19625 1377 19659 1411
rect 23305 1377 23339 1411
rect 27804 1377 27838 1411
rect 5825 1309 5859 1343
rect 6193 1309 6227 1343
rect 8309 1309 8343 1343
rect 9137 1309 9171 1343
rect 9321 1309 9355 1343
rect 12633 1309 12667 1343
rect 15945 1309 15979 1343
rect 18797 1309 18831 1343
rect 26249 1309 26283 1343
rect 26433 1309 26467 1343
rect 27537 1309 27571 1343
rect 5917 1241 5951 1275
rect 8217 1241 8251 1275
rect 12357 1241 12391 1275
rect 22661 1241 22695 1275
rect 6009 1173 6043 1207
rect 7665 1173 7699 1207
rect 8677 1173 8711 1207
rect 19165 1173 19199 1207
rect 19349 1173 19383 1207
rect 23029 1173 23063 1207
rect 26801 1173 26835 1207
rect 6929 969 6963 1003
rect 7021 969 7055 1003
rect 7205 969 7239 1003
rect 7389 969 7423 1003
rect 8861 969 8895 1003
rect 9045 969 9079 1003
rect 18705 969 18739 1003
rect 18889 969 18923 1003
rect 6837 833 6871 867
rect 7113 765 7147 799
rect 8401 765 8435 799
rect 8677 765 8711 799
rect 8953 765 8987 799
rect 18337 765 18371 799
rect 18429 765 18463 799
rect 19349 765 19383 799
rect 19616 765 19650 799
rect 7373 697 7407 731
rect 7573 697 7607 731
rect 8493 697 8527 731
rect 18873 697 18907 731
rect 19073 697 19107 731
rect 20729 629 20763 663
<< metal1 >>
rect 552 21786 31648 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 11436 21786
rect 11488 21734 11500 21786
rect 11552 21734 11564 21786
rect 11616 21734 11628 21786
rect 11680 21734 11692 21786
rect 11744 21734 19210 21786
rect 19262 21734 19274 21786
rect 19326 21734 19338 21786
rect 19390 21734 19402 21786
rect 19454 21734 19466 21786
rect 19518 21734 26984 21786
rect 27036 21734 27048 21786
rect 27100 21734 27112 21786
rect 27164 21734 27176 21786
rect 27228 21734 27240 21786
rect 27292 21734 31648 21786
rect 552 21712 31648 21734
rect 6086 21632 6092 21684
rect 6144 21632 6150 21684
rect 8018 21632 8024 21684
rect 8076 21632 8082 21684
rect 8386 21632 8392 21684
rect 8444 21632 8450 21684
rect 8662 21632 8668 21684
rect 8720 21632 8726 21684
rect 11701 21675 11759 21681
rect 11701 21641 11713 21675
rect 11747 21672 11759 21675
rect 11790 21672 11796 21684
rect 11747 21644 11796 21672
rect 11747 21641 11759 21644
rect 11701 21635 11759 21641
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12250 21632 12256 21684
rect 12308 21632 12314 21684
rect 12986 21632 12992 21684
rect 13044 21632 13050 21684
rect 18049 21675 18107 21681
rect 18049 21641 18061 21675
rect 18095 21672 18107 21675
rect 18782 21672 18788 21684
rect 18095 21644 18788 21672
rect 18095 21641 18107 21644
rect 18049 21635 18107 21641
rect 18782 21632 18788 21644
rect 18840 21632 18846 21684
rect 27893 21675 27951 21681
rect 27893 21641 27905 21675
rect 27939 21672 27951 21675
rect 29270 21672 29276 21684
rect 27939 21644 29276 21672
rect 27939 21641 27951 21644
rect 27893 21635 27951 21641
rect 29270 21632 29276 21644
rect 29328 21632 29334 21684
rect 7190 21536 7196 21548
rect 6288 21508 7196 21536
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 2225 21471 2283 21477
rect 2225 21468 2237 21471
rect 1452 21440 2237 21468
rect 1452 21428 1458 21440
rect 2225 21437 2237 21440
rect 2271 21437 2283 21471
rect 2225 21431 2283 21437
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21437 2835 21471
rect 2777 21431 2835 21437
rect 2792 21400 2820 21431
rect 2958 21428 2964 21480
rect 3016 21428 3022 21480
rect 4154 21428 4160 21480
rect 4212 21468 4218 21480
rect 5169 21471 5227 21477
rect 5169 21468 5181 21471
rect 4212 21440 5181 21468
rect 4212 21428 4218 21440
rect 5169 21437 5181 21440
rect 5215 21468 5227 21471
rect 5350 21468 5356 21480
rect 5215 21440 5356 21468
rect 5215 21437 5227 21440
rect 5169 21431 5227 21437
rect 5350 21428 5356 21440
rect 5408 21468 5414 21480
rect 6288 21477 6316 21508
rect 7190 21496 7196 21508
rect 7248 21536 7254 21548
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 7248 21508 7849 21536
rect 7248 21496 7254 21508
rect 7837 21505 7849 21508
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 13906 21496 13912 21548
rect 13964 21536 13970 21548
rect 14093 21539 14151 21545
rect 14093 21536 14105 21539
rect 13964 21508 14105 21536
rect 13964 21496 13970 21508
rect 14093 21505 14105 21508
rect 14139 21505 14151 21539
rect 14093 21499 14151 21505
rect 23658 21496 23664 21548
rect 23716 21536 23722 21548
rect 24673 21539 24731 21545
rect 24673 21536 24685 21539
rect 23716 21508 24685 21536
rect 23716 21496 23722 21508
rect 24673 21505 24685 21508
rect 24719 21505 24731 21539
rect 24673 21499 24731 21505
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 5408 21440 5457 21468
rect 5408 21428 5414 21440
rect 5445 21437 5457 21440
rect 5491 21437 5503 21471
rect 5445 21431 5503 21437
rect 6273 21471 6331 21477
rect 6273 21437 6285 21471
rect 6319 21437 6331 21471
rect 6273 21431 6331 21437
rect 6457 21471 6515 21477
rect 6457 21437 6469 21471
rect 6503 21437 6515 21471
rect 6457 21431 6515 21437
rect 6733 21471 6791 21477
rect 6733 21437 6745 21471
rect 6779 21468 6791 21471
rect 6914 21468 6920 21480
rect 6779 21440 6920 21468
rect 6779 21437 6791 21440
rect 6733 21431 6791 21437
rect 3142 21400 3148 21412
rect 2792 21372 3148 21400
rect 3142 21360 3148 21372
rect 3200 21360 3206 21412
rect 5537 21403 5595 21409
rect 5537 21369 5549 21403
rect 5583 21400 5595 21403
rect 6472 21400 6500 21431
rect 6914 21428 6920 21440
rect 6972 21428 6978 21480
rect 12802 21428 12808 21480
rect 12860 21468 12866 21480
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12860 21440 12909 21468
rect 12860 21428 12866 21440
rect 12897 21437 12909 21440
rect 12943 21437 12955 21471
rect 12897 21431 12955 21437
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21468 17187 21471
rect 19610 21468 19616 21480
rect 17175 21440 19616 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 19610 21428 19616 21440
rect 19668 21468 19674 21480
rect 20622 21468 20628 21480
rect 19668 21440 20628 21468
rect 19668 21428 19674 21440
rect 20622 21428 20628 21440
rect 20680 21468 20686 21480
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 20680 21440 21557 21468
rect 20680 21428 20686 21440
rect 21545 21437 21557 21440
rect 21591 21437 21603 21471
rect 21545 21431 21603 21437
rect 22097 21471 22155 21477
rect 22097 21437 22109 21471
rect 22143 21437 22155 21471
rect 22097 21431 22155 21437
rect 5583 21372 6500 21400
rect 5583 21369 5595 21372
rect 5537 21363 5595 21369
rect 7006 21360 7012 21412
rect 7064 21360 7070 21412
rect 7193 21403 7251 21409
rect 7193 21369 7205 21403
rect 7239 21400 7251 21403
rect 7285 21403 7343 21409
rect 7285 21400 7297 21403
rect 7239 21372 7297 21400
rect 7239 21369 7251 21372
rect 7193 21363 7251 21369
rect 7285 21369 7297 21372
rect 7331 21369 7343 21403
rect 7285 21363 7343 21369
rect 13909 21403 13967 21409
rect 13909 21369 13921 21403
rect 13955 21400 13967 21403
rect 14642 21400 14648 21412
rect 13955 21372 14648 21400
rect 13955 21369 13967 21372
rect 13909 21363 13967 21369
rect 14642 21360 14648 21372
rect 14700 21360 14706 21412
rect 17862 21360 17868 21412
rect 17920 21360 17926 21412
rect 18046 21360 18052 21412
rect 18104 21409 18110 21412
rect 18104 21403 18123 21409
rect 18111 21369 18123 21403
rect 22112 21400 22140 21431
rect 22186 21428 22192 21480
rect 22244 21428 22250 21480
rect 23842 21428 23848 21480
rect 23900 21428 23906 21480
rect 24394 21428 24400 21480
rect 24452 21428 24458 21480
rect 26418 21428 26424 21480
rect 26476 21428 26482 21480
rect 26694 21428 26700 21480
rect 26752 21428 26758 21480
rect 27157 21471 27215 21477
rect 27157 21437 27169 21471
rect 27203 21468 27215 21471
rect 27338 21468 27344 21480
rect 27203 21440 27344 21468
rect 27203 21437 27215 21440
rect 27157 21431 27215 21437
rect 27338 21428 27344 21440
rect 27396 21428 27402 21480
rect 27706 21428 27712 21480
rect 27764 21428 27770 21480
rect 28258 21428 28264 21480
rect 28316 21428 28322 21480
rect 28994 21428 29000 21480
rect 29052 21428 29058 21480
rect 24670 21400 24676 21412
rect 22112 21372 24676 21400
rect 18104 21363 18123 21369
rect 18104 21360 18110 21363
rect 24670 21360 24676 21372
rect 24728 21360 24734 21412
rect 24940 21403 24998 21409
rect 24940 21369 24952 21403
rect 24986 21400 24998 21403
rect 25130 21400 25136 21412
rect 24986 21372 25136 21400
rect 24986 21369 24998 21372
rect 24940 21363 24998 21369
rect 25130 21360 25136 21372
rect 25188 21360 25194 21412
rect 29242 21403 29300 21409
rect 29242 21400 29254 21403
rect 26620 21372 29254 21400
rect 1946 21292 1952 21344
rect 2004 21332 2010 21344
rect 2133 21335 2191 21341
rect 2133 21332 2145 21335
rect 2004 21304 2145 21332
rect 2004 21292 2010 21304
rect 2133 21301 2145 21304
rect 2179 21301 2191 21335
rect 2133 21295 2191 21301
rect 2866 21292 2872 21344
rect 2924 21292 2930 21344
rect 5258 21292 5264 21344
rect 5316 21292 5322 21344
rect 6638 21292 6644 21344
rect 6696 21292 6702 21344
rect 6822 21292 6828 21344
rect 6880 21292 6886 21344
rect 12618 21292 12624 21344
rect 12676 21332 12682 21344
rect 12805 21335 12863 21341
rect 12805 21332 12817 21335
rect 12676 21304 12817 21332
rect 12676 21292 12682 21304
rect 12805 21301 12817 21304
rect 12851 21301 12863 21335
rect 12805 21295 12863 21301
rect 12986 21292 12992 21344
rect 13044 21332 13050 21344
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 13044 21304 13553 21332
rect 13044 21292 13050 21304
rect 13541 21301 13553 21304
rect 13587 21301 13599 21335
rect 13541 21295 13599 21301
rect 13998 21292 14004 21344
rect 14056 21292 14062 21344
rect 16850 21292 16856 21344
rect 16908 21332 16914 21344
rect 17037 21335 17095 21341
rect 17037 21332 17049 21335
rect 16908 21304 17049 21332
rect 16908 21292 16914 21304
rect 17037 21301 17049 21304
rect 17083 21301 17095 21335
rect 17037 21295 17095 21301
rect 18230 21292 18236 21344
rect 18288 21292 18294 21344
rect 21266 21292 21272 21344
rect 21324 21332 21330 21344
rect 21453 21335 21511 21341
rect 21453 21332 21465 21335
rect 21324 21304 21465 21332
rect 21324 21292 21330 21304
rect 21453 21301 21465 21304
rect 21499 21301 21511 21335
rect 21453 21295 21511 21301
rect 21818 21292 21824 21344
rect 21876 21332 21882 21344
rect 21913 21335 21971 21341
rect 21913 21332 21925 21335
rect 21876 21304 21925 21332
rect 21876 21292 21882 21304
rect 21913 21301 21925 21304
rect 21959 21301 21971 21335
rect 21913 21295 21971 21301
rect 22370 21292 22376 21344
rect 22428 21292 22434 21344
rect 24026 21292 24032 21344
rect 24084 21292 24090 21344
rect 24578 21292 24584 21344
rect 24636 21292 24642 21344
rect 26050 21292 26056 21344
rect 26108 21292 26114 21344
rect 26620 21341 26648 21372
rect 29242 21369 29254 21372
rect 29288 21369 29300 21403
rect 29242 21363 29300 21369
rect 26605 21335 26663 21341
rect 26605 21301 26617 21335
rect 26651 21301 26663 21335
rect 26605 21295 26663 21301
rect 26881 21335 26939 21341
rect 26881 21301 26893 21335
rect 26927 21332 26939 21335
rect 27062 21332 27068 21344
rect 26927 21304 27068 21332
rect 26927 21301 26939 21304
rect 26881 21295 26939 21301
rect 27062 21292 27068 21304
rect 27120 21292 27126 21344
rect 27338 21292 27344 21344
rect 27396 21292 27402 21344
rect 28445 21335 28503 21341
rect 28445 21301 28457 21335
rect 28491 21332 28503 21335
rect 30098 21332 30104 21344
rect 28491 21304 30104 21332
rect 28491 21301 28503 21304
rect 28445 21295 28503 21301
rect 30098 21292 30104 21304
rect 30156 21292 30162 21344
rect 30374 21292 30380 21344
rect 30432 21292 30438 21344
rect 552 21242 31648 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 12096 21242
rect 12148 21190 12160 21242
rect 12212 21190 12224 21242
rect 12276 21190 12288 21242
rect 12340 21190 12352 21242
rect 12404 21190 19870 21242
rect 19922 21190 19934 21242
rect 19986 21190 19998 21242
rect 20050 21190 20062 21242
rect 20114 21190 20126 21242
rect 20178 21190 27644 21242
rect 27696 21190 27708 21242
rect 27760 21190 27772 21242
rect 27824 21190 27836 21242
rect 27888 21190 27900 21242
rect 27952 21190 31648 21242
rect 552 21168 31648 21190
rect 2958 21088 2964 21140
rect 3016 21128 3022 21140
rect 3513 21131 3571 21137
rect 3513 21128 3525 21131
rect 3016 21100 3525 21128
rect 3016 21088 3022 21100
rect 3513 21097 3525 21100
rect 3559 21097 3571 21131
rect 6822 21128 6828 21140
rect 3513 21091 3571 21097
rect 6472 21100 6828 21128
rect 6080 21063 6138 21069
rect 6080 21029 6092 21063
rect 6126 21060 6138 21063
rect 6472 21060 6500 21100
rect 6822 21088 6828 21100
rect 6880 21088 6886 21140
rect 7190 21088 7196 21140
rect 7248 21128 7254 21140
rect 8110 21128 8116 21140
rect 7248 21100 8116 21128
rect 7248 21088 7254 21100
rect 8110 21088 8116 21100
rect 8168 21128 8174 21140
rect 8168 21100 8432 21128
rect 8168 21088 8174 21100
rect 6126 21032 6500 21060
rect 6126 21029 6138 21032
rect 6080 21023 6138 21029
rect 6638 21020 6644 21072
rect 6696 21060 6702 21072
rect 6696 21032 8064 21060
rect 6696 21020 6702 21032
rect 1946 20952 1952 21004
rect 2004 20952 2010 21004
rect 2216 20995 2274 21001
rect 2216 20961 2228 20995
rect 2262 20992 2274 20995
rect 2498 20992 2504 21004
rect 2262 20964 2504 20992
rect 2262 20961 2274 20964
rect 2216 20955 2274 20961
rect 2498 20952 2504 20964
rect 2556 20952 2562 21004
rect 3510 20952 3516 21004
rect 3568 20992 3574 21004
rect 3697 20995 3755 21001
rect 3697 20992 3709 20995
rect 3568 20964 3709 20992
rect 3568 20952 3574 20964
rect 3697 20961 3709 20964
rect 3743 20961 3755 20995
rect 3697 20955 3755 20961
rect 3881 20995 3939 21001
rect 3881 20961 3893 20995
rect 3927 20992 3939 20995
rect 4062 20992 4068 21004
rect 3927 20964 4068 20992
rect 3927 20961 3939 20964
rect 3881 20955 3939 20961
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 4154 20952 4160 21004
rect 4212 20952 4218 21004
rect 4706 20952 4712 21004
rect 4764 20952 4770 21004
rect 4890 20952 4896 21004
rect 4948 20952 4954 21004
rect 5258 20952 5264 21004
rect 5316 20992 5322 21004
rect 5813 20995 5871 21001
rect 5813 20992 5825 20995
rect 5316 20964 5825 20992
rect 5316 20952 5322 20964
rect 5813 20961 5825 20964
rect 5859 20961 5871 20995
rect 5813 20955 5871 20961
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 8036 21001 8064 21032
rect 8404 21001 8432 21100
rect 8570 21088 8576 21140
rect 8628 21088 8634 21140
rect 8938 21088 8944 21140
rect 8996 21088 9002 21140
rect 9766 21088 9772 21140
rect 9824 21088 9830 21140
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21128 14795 21131
rect 17862 21128 17868 21140
rect 14783 21100 17868 21128
rect 14783 21097 14795 21100
rect 14737 21091 14795 21097
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 18046 21088 18052 21140
rect 18104 21128 18110 21140
rect 18785 21131 18843 21137
rect 18785 21128 18797 21131
rect 18104 21100 18797 21128
rect 18104 21088 18110 21100
rect 18785 21097 18797 21100
rect 18831 21097 18843 21131
rect 18785 21091 18843 21097
rect 19518 21088 19524 21140
rect 19576 21128 19582 21140
rect 22186 21128 22192 21140
rect 19576 21100 22192 21128
rect 19576 21088 19582 21100
rect 22186 21088 22192 21100
rect 22244 21128 22250 21140
rect 22649 21131 22707 21137
rect 22649 21128 22661 21131
rect 22244 21100 22661 21128
rect 22244 21088 22250 21100
rect 22649 21097 22661 21100
rect 22695 21097 22707 21131
rect 22649 21091 22707 21097
rect 25130 21088 25136 21140
rect 25188 21088 25194 21140
rect 27338 21088 27344 21140
rect 27396 21128 27402 21140
rect 30127 21131 30185 21137
rect 27396 21100 28580 21128
rect 27396 21088 27402 21100
rect 8772 21032 9628 21060
rect 8772 21001 8800 21032
rect 7561 20995 7619 21001
rect 7561 20992 7573 20995
rect 6972 20964 7573 20992
rect 6972 20952 6978 20964
rect 7561 20961 7573 20964
rect 7607 20961 7619 20995
rect 7561 20955 7619 20961
rect 8021 20995 8079 21001
rect 8021 20961 8033 20995
rect 8067 20961 8079 20995
rect 8021 20955 8079 20961
rect 8389 20995 8447 21001
rect 8389 20961 8401 20995
rect 8435 20992 8447 20995
rect 8757 20995 8815 21001
rect 8757 20992 8769 20995
rect 8435 20964 8769 20992
rect 8435 20961 8447 20964
rect 8389 20955 8447 20961
rect 8757 20961 8769 20964
rect 8803 20961 8815 20995
rect 8757 20955 8815 20961
rect 9309 20995 9367 21001
rect 9309 20961 9321 20995
rect 9355 20992 9367 20995
rect 9398 20992 9404 21004
rect 9355 20964 9404 20992
rect 9355 20961 9367 20964
rect 9309 20955 9367 20961
rect 9398 20952 9404 20964
rect 9456 20952 9462 21004
rect 9490 20952 9496 21004
rect 9548 20952 9554 21004
rect 9600 21001 9628 21032
rect 18230 21020 18236 21072
rect 18288 21060 18294 21072
rect 23928 21063 23986 21069
rect 18288 21032 19932 21060
rect 18288 21020 18294 21032
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20961 9643 20995
rect 9585 20955 9643 20961
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 10413 20995 10471 21001
rect 10413 20992 10425 20995
rect 9732 20964 10425 20992
rect 9732 20952 9738 20964
rect 10413 20961 10425 20964
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 11238 20952 11244 21004
rect 11296 20952 11302 21004
rect 12618 20952 12624 21004
rect 12676 20952 12682 21004
rect 16850 20952 16856 21004
rect 16908 20952 16914 21004
rect 17126 21001 17132 21004
rect 17120 20955 17132 21001
rect 17126 20952 17132 20955
rect 17184 20952 17190 21004
rect 18322 20952 18328 21004
rect 18380 20992 18386 21004
rect 18877 20995 18935 21001
rect 18877 20992 18889 20995
rect 18380 20964 18889 20992
rect 18380 20952 18386 20964
rect 18877 20961 18889 20964
rect 18923 20992 18935 20995
rect 19058 20992 19064 21004
rect 18923 20964 19064 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 19424 20995 19482 21001
rect 19424 20961 19436 20995
rect 19470 20961 19482 20995
rect 19424 20955 19482 20961
rect 8846 20884 8852 20936
rect 8904 20924 8910 20936
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 8904 20896 9137 20924
rect 8904 20884 8910 20896
rect 9125 20893 9137 20896
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 12894 20884 12900 20936
rect 12952 20884 12958 20936
rect 14826 20884 14832 20936
rect 14884 20884 14890 20936
rect 14918 20884 14924 20936
rect 14976 20884 14982 20936
rect 18690 20884 18696 20936
rect 18748 20924 18754 20936
rect 18969 20927 19027 20933
rect 18969 20924 18981 20927
rect 18748 20896 18981 20924
rect 18748 20884 18754 20896
rect 18969 20893 18981 20896
rect 19015 20893 19027 20927
rect 18969 20887 19027 20893
rect 3234 20816 3240 20868
rect 3292 20856 3298 20868
rect 4065 20859 4123 20865
rect 4065 20856 4077 20859
rect 3292 20828 4077 20856
rect 3292 20816 3298 20828
rect 4065 20825 4077 20828
rect 4111 20825 4123 20859
rect 4065 20819 4123 20825
rect 13630 20816 13636 20868
rect 13688 20856 13694 20868
rect 14369 20859 14427 20865
rect 14369 20856 14381 20859
rect 13688 20828 14381 20856
rect 13688 20816 13694 20828
rect 14369 20825 14381 20828
rect 14415 20825 14427 20859
rect 14369 20819 14427 20825
rect 17862 20816 17868 20868
rect 17920 20856 17926 20868
rect 18417 20859 18475 20865
rect 18417 20856 18429 20859
rect 17920 20828 18429 20856
rect 17920 20816 17926 20828
rect 18417 20825 18429 20828
rect 18463 20825 18475 20859
rect 19444 20856 19472 20955
rect 19518 20952 19524 21004
rect 19576 20952 19582 21004
rect 19613 20995 19671 21001
rect 19613 20961 19625 20995
rect 19659 20961 19671 20995
rect 19613 20955 19671 20961
rect 19628 20924 19656 20955
rect 19702 20952 19708 21004
rect 19760 21001 19766 21004
rect 19904 21001 19932 21032
rect 23928 21029 23940 21063
rect 23974 21060 23986 21063
rect 24026 21060 24032 21072
rect 23974 21032 24032 21060
rect 23974 21029 23986 21032
rect 23928 21023 23986 21029
rect 24026 21020 24032 21032
rect 24084 21020 24090 21072
rect 28552 21060 28580 21100
rect 30127 21097 30139 21131
rect 30173 21128 30185 21131
rect 30374 21128 30380 21140
rect 30173 21100 30380 21128
rect 30173 21097 30185 21100
rect 30127 21091 30185 21097
rect 30374 21088 30380 21100
rect 30432 21088 30438 21140
rect 28690 21063 28748 21069
rect 28690 21060 28702 21063
rect 26988 21032 28488 21060
rect 28552 21032 28702 21060
rect 19760 20995 19799 21001
rect 19787 20961 19799 20995
rect 19760 20955 19799 20961
rect 19889 20995 19947 21001
rect 19889 20961 19901 20995
rect 19935 20961 19947 20995
rect 19889 20955 19947 20961
rect 19760 20952 19766 20955
rect 20622 20952 20628 21004
rect 20680 20992 20686 21004
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 20680 20964 20913 20992
rect 20680 20952 20686 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 21266 20952 21272 21004
rect 21324 20952 21330 21004
rect 21818 20992 21824 21004
rect 21376 20964 21824 20992
rect 19978 20924 19984 20936
rect 19628 20896 19984 20924
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 21376 20924 21404 20964
rect 21818 20952 21824 20964
rect 21876 20952 21882 21004
rect 25314 20952 25320 21004
rect 25372 20952 25378 21004
rect 25498 20952 25504 21004
rect 25556 20952 25562 21004
rect 20772 20896 21404 20924
rect 20772 20884 20778 20896
rect 21542 20884 21548 20936
rect 21600 20884 21606 20936
rect 23658 20884 23664 20936
rect 23716 20884 23722 20936
rect 25866 20884 25872 20936
rect 25924 20924 25930 20936
rect 26988 20933 27016 21032
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 28460 21001 28488 21032
rect 28690 21029 28702 21032
rect 28736 21029 28748 21063
rect 28690 21023 28748 21029
rect 29178 21020 29184 21072
rect 29236 21060 29242 21072
rect 29917 21063 29975 21069
rect 29917 21060 29929 21063
rect 29236 21032 29929 21060
rect 29236 21020 29242 21032
rect 29917 21029 29929 21032
rect 29963 21029 29975 21063
rect 29917 21023 29975 21029
rect 27229 20995 27287 21001
rect 27229 20992 27241 20995
rect 27120 20964 27241 20992
rect 27120 20952 27126 20964
rect 27229 20961 27241 20964
rect 27275 20961 27287 20995
rect 27229 20955 27287 20961
rect 28445 20995 28503 21001
rect 28445 20961 28457 20995
rect 28491 20961 28503 20995
rect 28445 20955 28503 20961
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 25924 20896 26985 20924
rect 25924 20884 25930 20896
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 19794 20856 19800 20868
rect 19444 20828 19800 20856
rect 18417 20819 18475 20825
rect 19794 20816 19800 20828
rect 19852 20816 19858 20868
rect 29454 20816 29460 20868
rect 29512 20856 29518 20868
rect 30285 20859 30343 20865
rect 30285 20856 30297 20859
rect 29512 20828 30297 20856
rect 29512 20816 29518 20828
rect 30285 20825 30297 20828
rect 30331 20825 30343 20859
rect 30285 20819 30343 20825
rect 3326 20748 3332 20800
rect 3384 20748 3390 20800
rect 4798 20748 4804 20800
rect 4856 20748 4862 20800
rect 7834 20748 7840 20800
rect 7892 20748 7898 20800
rect 8202 20748 8208 20800
rect 8260 20748 8266 20800
rect 10321 20791 10379 20797
rect 10321 20757 10333 20791
rect 10367 20788 10379 20791
rect 11054 20788 11060 20800
rect 10367 20760 11060 20788
rect 10367 20757 10379 20760
rect 10321 20751 10379 20757
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11517 20791 11575 20797
rect 11517 20757 11529 20791
rect 11563 20788 11575 20791
rect 13262 20788 13268 20800
rect 11563 20760 13268 20788
rect 11563 20757 11575 20760
rect 11517 20751 11575 20757
rect 13262 20748 13268 20760
rect 13320 20748 13326 20800
rect 14182 20748 14188 20800
rect 14240 20788 14246 20800
rect 15194 20788 15200 20800
rect 14240 20760 15200 20788
rect 14240 20748 14246 20760
rect 15194 20748 15200 20760
rect 15252 20748 15258 20800
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 18233 20791 18291 20797
rect 18233 20788 18245 20791
rect 18104 20760 18245 20788
rect 18104 20748 18110 20760
rect 18233 20757 18245 20760
rect 18279 20757 18291 20791
rect 18233 20751 18291 20757
rect 18506 20748 18512 20800
rect 18564 20788 18570 20800
rect 19245 20791 19303 20797
rect 19245 20788 19257 20791
rect 18564 20760 19257 20788
rect 18564 20748 18570 20760
rect 19245 20757 19257 20760
rect 19291 20757 19303 20791
rect 19245 20751 19303 20757
rect 20990 20748 20996 20800
rect 21048 20748 21054 20800
rect 25041 20791 25099 20797
rect 25041 20757 25053 20791
rect 25087 20788 25099 20791
rect 25314 20788 25320 20800
rect 25087 20760 25320 20788
rect 25087 20757 25099 20760
rect 25041 20751 25099 20757
rect 25314 20748 25320 20760
rect 25372 20748 25378 20800
rect 25685 20791 25743 20797
rect 25685 20757 25697 20791
rect 25731 20788 25743 20791
rect 25958 20788 25964 20800
rect 25731 20760 25964 20788
rect 25731 20757 25743 20760
rect 25685 20751 25743 20757
rect 25958 20748 25964 20760
rect 26016 20748 26022 20800
rect 28350 20748 28356 20800
rect 28408 20748 28414 20800
rect 29362 20748 29368 20800
rect 29420 20788 29426 20800
rect 29825 20791 29883 20797
rect 29825 20788 29837 20791
rect 29420 20760 29837 20788
rect 29420 20748 29426 20760
rect 29825 20757 29837 20760
rect 29871 20757 29883 20791
rect 29825 20751 29883 20757
rect 30006 20748 30012 20800
rect 30064 20788 30070 20800
rect 30101 20791 30159 20797
rect 30101 20788 30113 20791
rect 30064 20760 30113 20788
rect 30064 20748 30070 20760
rect 30101 20757 30113 20760
rect 30147 20757 30159 20791
rect 30101 20751 30159 20757
rect 552 20698 31648 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 11436 20698
rect 11488 20646 11500 20698
rect 11552 20646 11564 20698
rect 11616 20646 11628 20698
rect 11680 20646 11692 20698
rect 11744 20646 19210 20698
rect 19262 20646 19274 20698
rect 19326 20646 19338 20698
rect 19390 20646 19402 20698
rect 19454 20646 19466 20698
rect 19518 20646 26984 20698
rect 27036 20646 27048 20698
rect 27100 20646 27112 20698
rect 27164 20646 27176 20698
rect 27228 20646 27240 20698
rect 27292 20646 31648 20698
rect 552 20624 31648 20646
rect 1394 20544 1400 20596
rect 1452 20584 1458 20596
rect 4154 20584 4160 20596
rect 1452 20556 4160 20584
rect 1452 20544 1458 20556
rect 4154 20544 4160 20556
rect 4212 20544 4218 20596
rect 4801 20587 4859 20593
rect 4801 20553 4813 20587
rect 4847 20584 4859 20587
rect 4890 20584 4896 20596
rect 4847 20556 4896 20584
rect 4847 20553 4859 20556
rect 4801 20547 4859 20553
rect 4890 20544 4896 20556
rect 4948 20544 4954 20596
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7009 20587 7067 20593
rect 7009 20584 7021 20587
rect 6972 20556 7021 20584
rect 6972 20544 6978 20556
rect 7009 20553 7021 20556
rect 7055 20553 7067 20587
rect 7009 20547 7067 20553
rect 9585 20587 9643 20593
rect 9585 20553 9597 20587
rect 9631 20584 9643 20587
rect 9674 20584 9680 20596
rect 9631 20556 9680 20584
rect 9631 20553 9643 20556
rect 9585 20547 9643 20553
rect 4617 20519 4675 20525
rect 4617 20485 4629 20519
rect 4663 20485 4675 20519
rect 4617 20479 4675 20485
rect 3234 20408 3240 20460
rect 3292 20408 3298 20460
rect 4632 20448 4660 20479
rect 5353 20451 5411 20457
rect 5353 20448 5365 20451
rect 4632 20420 5365 20448
rect 1302 20340 1308 20392
rect 1360 20340 1366 20392
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1581 20383 1639 20389
rect 1581 20380 1593 20383
rect 1443 20352 1593 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1581 20349 1593 20352
rect 1627 20349 1639 20383
rect 1581 20343 1639 20349
rect 3878 20340 3884 20392
rect 3936 20380 3942 20392
rect 4632 20380 4660 20420
rect 5353 20417 5365 20420
rect 5399 20448 5411 20451
rect 7024 20448 7052 20547
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 12894 20544 12900 20596
rect 12952 20584 12958 20596
rect 13541 20587 13599 20593
rect 13541 20584 13553 20587
rect 12952 20556 13553 20584
rect 12952 20544 12958 20556
rect 13541 20553 13553 20556
rect 13587 20553 13599 20587
rect 14550 20584 14556 20596
rect 13541 20547 13599 20553
rect 13924 20556 14556 20584
rect 13924 20528 13952 20556
rect 14550 20544 14556 20556
rect 14608 20544 14614 20596
rect 14826 20544 14832 20596
rect 14884 20584 14890 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 14884 20556 15025 20584
rect 14884 20544 14890 20556
rect 15013 20553 15025 20556
rect 15059 20553 15071 20587
rect 16482 20584 16488 20596
rect 15013 20547 15071 20553
rect 15396 20556 16488 20584
rect 9309 20519 9367 20525
rect 9309 20485 9321 20519
rect 9355 20516 9367 20519
rect 9398 20516 9404 20528
rect 9355 20488 9404 20516
rect 9355 20485 9367 20488
rect 9309 20479 9367 20485
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 13357 20519 13415 20525
rect 13357 20516 13369 20519
rect 13280 20488 13369 20516
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 5399 20420 5764 20448
rect 7024 20420 7665 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 3936 20352 4660 20380
rect 3936 20340 3942 20352
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5500 20352 5641 20380
rect 5500 20340 5506 20352
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 5736 20380 5764 20420
rect 7653 20417 7665 20420
rect 7699 20417 7711 20451
rect 7653 20411 7711 20417
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 9950 20448 9956 20460
rect 9640 20420 9956 20448
rect 9640 20408 9646 20420
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 12161 20451 12219 20457
rect 10888 20420 11284 20448
rect 6914 20380 6920 20392
rect 5736 20352 6920 20380
rect 5629 20343 5687 20349
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 8110 20340 8116 20392
rect 8168 20340 8174 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 8665 20383 8723 20389
rect 8665 20380 8677 20383
rect 8352 20352 8677 20380
rect 8352 20340 8358 20352
rect 8665 20349 8677 20352
rect 8711 20380 8723 20383
rect 10888 20380 10916 20420
rect 11256 20389 11284 20420
rect 12161 20417 12173 20451
rect 12207 20448 12219 20451
rect 12618 20448 12624 20460
rect 12207 20420 12624 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20448 12863 20451
rect 13170 20448 13176 20460
rect 12851 20420 13176 20448
rect 12851 20417 12863 20420
rect 12805 20411 12863 20417
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 8711 20352 10916 20380
rect 10965 20383 11023 20389
rect 8711 20349 8723 20352
rect 8665 20343 8723 20349
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11149 20383 11207 20389
rect 11149 20380 11161 20383
rect 11011 20352 11161 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 11149 20349 11161 20352
rect 11195 20349 11207 20383
rect 11149 20343 11207 20349
rect 11241 20383 11299 20389
rect 11241 20349 11253 20383
rect 11287 20380 11299 20383
rect 11885 20383 11943 20389
rect 11885 20380 11897 20383
rect 11287 20352 11897 20380
rect 11287 20349 11299 20352
rect 11241 20343 11299 20349
rect 11885 20349 11897 20352
rect 11931 20349 11943 20383
rect 11885 20343 11943 20349
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20380 12403 20383
rect 12986 20380 12992 20392
rect 12391 20352 12992 20380
rect 12391 20349 12403 20352
rect 12345 20343 12403 20349
rect 1848 20315 1906 20321
rect 1848 20281 1860 20315
rect 1894 20312 1906 20315
rect 2314 20312 2320 20324
rect 1894 20284 2320 20312
rect 1894 20281 1906 20284
rect 1848 20275 1906 20281
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 3050 20272 3056 20324
rect 3108 20312 3114 20324
rect 5902 20321 5908 20324
rect 3482 20315 3540 20321
rect 3482 20312 3494 20315
rect 3108 20284 3494 20312
rect 3108 20272 3114 20284
rect 3482 20281 3494 20284
rect 3528 20281 3540 20315
rect 3482 20275 3540 20281
rect 5896 20275 5908 20321
rect 5902 20272 5908 20275
rect 5960 20272 5966 20324
rect 6730 20272 6736 20324
rect 6788 20312 6794 20324
rect 8941 20315 8999 20321
rect 6788 20284 7972 20312
rect 6788 20272 6794 20284
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 2961 20247 3019 20253
rect 2961 20244 2973 20247
rect 2832 20216 2973 20244
rect 2832 20204 2838 20216
rect 2961 20213 2973 20216
rect 3007 20244 3019 20247
rect 3602 20244 3608 20256
rect 3007 20216 3608 20244
rect 3007 20213 3019 20216
rect 2961 20207 3019 20213
rect 3602 20204 3608 20216
rect 3660 20244 3666 20256
rect 3970 20244 3976 20256
rect 3660 20216 3976 20244
rect 3660 20204 3666 20216
rect 3970 20204 3976 20216
rect 4028 20204 4034 20256
rect 6086 20204 6092 20256
rect 6144 20244 6150 20256
rect 7944 20253 7972 20284
rect 8941 20281 8953 20315
rect 8987 20312 8999 20315
rect 9490 20312 9496 20324
rect 8987 20284 9496 20312
rect 8987 20281 8999 20284
rect 8941 20275 8999 20281
rect 9490 20272 9496 20284
rect 9548 20312 9554 20324
rect 9548 20284 9904 20312
rect 9548 20272 9554 20284
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 6144 20216 7113 20244
rect 6144 20204 6150 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7101 20207 7159 20213
rect 7929 20247 7987 20253
rect 7929 20213 7941 20247
rect 7975 20213 7987 20247
rect 7929 20207 7987 20213
rect 8757 20247 8815 20253
rect 8757 20213 8769 20247
rect 8803 20244 8815 20247
rect 9122 20244 9128 20256
rect 8803 20216 9128 20244
rect 8803 20213 8815 20216
rect 8757 20207 8815 20213
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 9401 20247 9459 20253
rect 9401 20213 9413 20247
rect 9447 20244 9459 20247
rect 9582 20244 9588 20256
rect 9447 20216 9588 20244
rect 9447 20213 9459 20216
rect 9401 20207 9459 20213
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 9876 20244 9904 20284
rect 9950 20272 9956 20324
rect 10008 20312 10014 20324
rect 10698 20315 10756 20321
rect 10698 20312 10710 20315
rect 10008 20284 10710 20312
rect 10008 20272 10014 20284
rect 10698 20281 10710 20284
rect 10744 20281 10756 20315
rect 11900 20312 11928 20343
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 13280 20380 13308 20488
rect 13357 20485 13369 20488
rect 13403 20485 13415 20519
rect 13357 20479 13415 20485
rect 13446 20476 13452 20528
rect 13504 20516 13510 20528
rect 13906 20516 13912 20528
rect 13504 20488 13912 20516
rect 13504 20476 13510 20488
rect 13906 20476 13912 20488
rect 13964 20476 13970 20528
rect 14274 20516 14280 20528
rect 14016 20488 14280 20516
rect 14016 20389 14044 20488
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 14642 20476 14648 20528
rect 14700 20516 14706 20528
rect 15396 20516 15424 20556
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 17126 20544 17132 20596
rect 17184 20544 17190 20596
rect 17770 20544 17776 20596
rect 17828 20584 17834 20596
rect 17957 20587 18015 20593
rect 17957 20584 17969 20587
rect 17828 20556 17969 20584
rect 17828 20544 17834 20556
rect 17957 20553 17969 20556
rect 18003 20553 18015 20587
rect 17957 20547 18015 20553
rect 18049 20587 18107 20593
rect 18049 20553 18061 20587
rect 18095 20584 18107 20587
rect 18506 20584 18512 20596
rect 18095 20556 18512 20584
rect 18095 20553 18107 20556
rect 18049 20547 18107 20553
rect 18506 20544 18512 20556
rect 18564 20544 18570 20596
rect 18782 20544 18788 20596
rect 18840 20584 18846 20596
rect 18877 20587 18935 20593
rect 18877 20584 18889 20587
rect 18840 20556 18889 20584
rect 18840 20544 18846 20556
rect 18877 20553 18889 20556
rect 18923 20553 18935 20587
rect 18877 20547 18935 20553
rect 18966 20544 18972 20596
rect 19024 20584 19030 20596
rect 19978 20584 19984 20596
rect 19024 20556 19984 20584
rect 19024 20544 19030 20556
rect 19978 20544 19984 20556
rect 20036 20584 20042 20596
rect 20898 20584 20904 20596
rect 20036 20556 20904 20584
rect 20036 20544 20042 20556
rect 20898 20544 20904 20556
rect 20956 20544 20962 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 21542 20584 21548 20596
rect 21131 20556 21548 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 25866 20584 25872 20596
rect 24412 20556 25872 20584
rect 14700 20488 15424 20516
rect 14700 20476 14706 20488
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14369 20451 14427 20457
rect 14369 20448 14381 20451
rect 14139 20420 14381 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14369 20417 14381 20420
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 14553 20451 14611 20457
rect 14553 20417 14565 20451
rect 14599 20448 14611 20451
rect 15194 20448 15200 20460
rect 14599 20420 15200 20448
rect 14599 20417 14611 20420
rect 14553 20411 14611 20417
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15396 20457 15424 20488
rect 15470 20476 15476 20528
rect 15528 20516 15534 20528
rect 15528 20488 15976 20516
rect 15528 20476 15534 20488
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20417 15439 20451
rect 15381 20411 15439 20417
rect 15838 20408 15844 20460
rect 15896 20408 15902 20460
rect 15948 20448 15976 20488
rect 18690 20476 18696 20528
rect 18748 20476 18754 20528
rect 19702 20476 19708 20528
rect 19760 20516 19766 20528
rect 19760 20488 21220 20516
rect 19760 20476 19766 20488
rect 16114 20448 16120 20460
rect 15948 20420 16120 20448
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 16206 20408 16212 20460
rect 16264 20457 16270 20460
rect 16264 20451 16292 20457
rect 16280 20417 16292 20451
rect 17862 20448 17868 20460
rect 16264 20411 16292 20417
rect 17328 20420 17868 20448
rect 16264 20408 16270 20411
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 13280 20352 13737 20380
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 13909 20383 13967 20389
rect 13909 20349 13921 20383
rect 13955 20349 13967 20383
rect 13909 20343 13967 20349
rect 14001 20383 14059 20389
rect 14001 20349 14013 20383
rect 14047 20349 14059 20383
rect 14001 20343 14059 20349
rect 14185 20383 14243 20389
rect 14185 20349 14197 20383
rect 14231 20380 14243 20383
rect 14274 20380 14280 20392
rect 14231 20352 14280 20380
rect 14231 20349 14243 20352
rect 14185 20343 14243 20349
rect 12802 20312 12808 20324
rect 11900 20284 12808 20312
rect 10698 20275 10756 20281
rect 12802 20272 12808 20284
rect 12860 20272 12866 20324
rect 12897 20315 12955 20321
rect 12897 20281 12909 20315
rect 12943 20312 12955 20315
rect 13630 20312 13636 20324
rect 12943 20284 13636 20312
rect 12943 20281 12955 20284
rect 12897 20275 12955 20281
rect 13630 20272 13636 20284
rect 13688 20272 13694 20324
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 13924 20312 13952 20343
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 16390 20340 16396 20392
rect 16448 20340 16454 20392
rect 17328 20389 17356 20420
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20448 18015 20451
rect 18874 20448 18880 20460
rect 18003 20420 18880 20448
rect 18003 20417 18015 20420
rect 17957 20411 18015 20417
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 19058 20408 19064 20460
rect 19116 20448 19122 20460
rect 21082 20448 21088 20460
rect 19116 20420 21088 20448
rect 19116 20408 19122 20420
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20349 17371 20383
rect 17313 20343 17371 20349
rect 17494 20340 17500 20392
rect 17552 20340 17558 20392
rect 18138 20340 18144 20392
rect 18196 20340 18202 20392
rect 20346 20380 20352 20392
rect 19306 20352 20352 20380
rect 15286 20312 15292 20324
rect 13872 20284 15292 20312
rect 13872 20272 13878 20284
rect 15286 20272 15292 20284
rect 15344 20272 15350 20324
rect 17037 20315 17095 20321
rect 17037 20281 17049 20315
rect 17083 20312 17095 20315
rect 17773 20315 17831 20321
rect 17773 20312 17785 20315
rect 17083 20284 17785 20312
rect 17083 20281 17095 20284
rect 17037 20275 17095 20281
rect 17773 20281 17785 20284
rect 17819 20281 17831 20315
rect 17773 20275 17831 20281
rect 17954 20272 17960 20324
rect 18012 20312 18018 20324
rect 18506 20312 18512 20324
rect 18012 20284 18512 20312
rect 18012 20272 18018 20284
rect 18506 20272 18512 20284
rect 18564 20312 18570 20324
rect 19061 20315 19119 20321
rect 19061 20312 19073 20315
rect 18564 20284 19073 20312
rect 18564 20272 18570 20284
rect 19061 20281 19073 20284
rect 19107 20312 19119 20315
rect 19306 20312 19334 20352
rect 20346 20340 20352 20352
rect 20404 20340 20410 20392
rect 20441 20383 20499 20389
rect 20441 20349 20453 20383
rect 20487 20380 20499 20383
rect 20530 20380 20536 20392
rect 20487 20352 20536 20380
rect 20487 20349 20499 20352
rect 20441 20343 20499 20349
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 20625 20383 20683 20389
rect 20625 20349 20637 20383
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 19107 20284 19334 20312
rect 19107 20281 19119 20284
rect 19061 20275 19119 20281
rect 10134 20244 10140 20256
rect 9876 20216 10140 20244
rect 10134 20204 10140 20216
rect 10192 20204 10198 20256
rect 11974 20204 11980 20256
rect 12032 20204 12038 20256
rect 12526 20204 12532 20256
rect 12584 20204 12590 20256
rect 12989 20247 13047 20253
rect 12989 20213 13001 20247
rect 13035 20244 13047 20247
rect 14182 20244 14188 20256
rect 13035 20216 14188 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 14645 20247 14703 20253
rect 14645 20213 14657 20247
rect 14691 20244 14703 20247
rect 15194 20244 15200 20256
rect 14691 20216 15200 20244
rect 14691 20213 14703 20216
rect 14645 20207 14703 20213
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 18861 20247 18919 20253
rect 18861 20213 18873 20247
rect 18907 20244 18919 20247
rect 19150 20244 19156 20256
rect 18907 20216 19156 20244
rect 18907 20213 18919 20216
rect 18861 20207 18919 20213
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 20640 20244 20668 20343
rect 20714 20340 20720 20392
rect 20772 20340 20778 20392
rect 20824 20389 20852 20420
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 21192 20448 21220 20488
rect 22557 20451 22615 20457
rect 22557 20448 22569 20451
rect 21192 20420 22569 20448
rect 22557 20417 22569 20420
rect 22603 20448 22615 20451
rect 22603 20420 23152 20448
rect 22603 20417 22615 20420
rect 22557 20411 22615 20417
rect 20809 20383 20867 20389
rect 20809 20349 20821 20383
rect 20855 20349 20867 20383
rect 20809 20343 20867 20349
rect 20990 20340 20996 20392
rect 21048 20380 21054 20392
rect 21177 20383 21235 20389
rect 21177 20380 21189 20383
rect 21048 20352 21189 20380
rect 21048 20340 21054 20352
rect 21177 20349 21189 20352
rect 21223 20349 21235 20383
rect 21177 20343 21235 20349
rect 21266 20340 21272 20392
rect 21324 20380 21330 20392
rect 21453 20383 21511 20389
rect 21453 20380 21465 20383
rect 21324 20352 21465 20380
rect 21324 20340 21330 20352
rect 21453 20349 21465 20352
rect 21499 20349 21511 20383
rect 21453 20343 21511 20349
rect 21542 20340 21548 20392
rect 21600 20380 21606 20392
rect 23124 20389 23152 20420
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 24412 20457 24440 20556
rect 25866 20544 25872 20556
rect 25924 20544 25930 20596
rect 24397 20451 24455 20457
rect 24397 20448 24409 20451
rect 23716 20420 24409 20448
rect 23716 20408 23722 20420
rect 24397 20417 24409 20420
rect 24443 20417 24455 20451
rect 24397 20411 24455 20417
rect 23109 20383 23167 20389
rect 21600 20352 22140 20380
rect 21600 20340 21606 20352
rect 22112 20312 22140 20352
rect 23109 20349 23121 20383
rect 23155 20349 23167 20383
rect 23109 20343 23167 20349
rect 23382 20340 23388 20392
rect 23440 20340 23446 20392
rect 25884 20389 25912 20544
rect 24664 20383 24722 20389
rect 24664 20349 24676 20383
rect 24710 20349 24722 20383
rect 24664 20343 24722 20349
rect 25869 20383 25927 20389
rect 25869 20349 25881 20383
rect 25915 20349 25927 20383
rect 25869 20343 25927 20349
rect 22112 20284 23336 20312
rect 21910 20244 21916 20256
rect 20640 20216 21916 20244
rect 21910 20204 21916 20216
rect 21968 20204 21974 20256
rect 22922 20204 22928 20256
rect 22980 20204 22986 20256
rect 23308 20253 23336 20284
rect 24578 20272 24584 20324
rect 24636 20312 24642 20324
rect 24688 20312 24716 20343
rect 25958 20340 25964 20392
rect 26016 20380 26022 20392
rect 26125 20383 26183 20389
rect 26125 20380 26137 20383
rect 26016 20352 26137 20380
rect 26016 20340 26022 20352
rect 26125 20349 26137 20352
rect 26171 20349 26183 20383
rect 26125 20343 26183 20349
rect 28994 20340 29000 20392
rect 29052 20340 29058 20392
rect 29270 20389 29276 20392
rect 29264 20380 29276 20389
rect 29231 20352 29276 20380
rect 29264 20343 29276 20352
rect 29270 20340 29276 20343
rect 29328 20340 29334 20392
rect 24636 20284 24716 20312
rect 24636 20272 24642 20284
rect 23293 20247 23351 20253
rect 23293 20213 23305 20247
rect 23339 20244 23351 20247
rect 25406 20244 25412 20256
rect 23339 20216 25412 20244
rect 23339 20213 23351 20216
rect 23293 20207 23351 20213
rect 25406 20204 25412 20216
rect 25464 20204 25470 20256
rect 25777 20247 25835 20253
rect 25777 20213 25789 20247
rect 25823 20244 25835 20247
rect 26602 20244 26608 20256
rect 25823 20216 26608 20244
rect 25823 20213 25835 20216
rect 25777 20207 25835 20213
rect 26602 20204 26608 20216
rect 26660 20204 26666 20256
rect 26694 20204 26700 20256
rect 26752 20244 26758 20256
rect 27249 20247 27307 20253
rect 27249 20244 27261 20247
rect 26752 20216 27261 20244
rect 26752 20204 26758 20216
rect 27249 20213 27261 20216
rect 27295 20213 27307 20247
rect 27249 20207 27307 20213
rect 29086 20204 29092 20256
rect 29144 20244 29150 20256
rect 30377 20247 30435 20253
rect 30377 20244 30389 20247
rect 29144 20216 30389 20244
rect 29144 20204 29150 20216
rect 30377 20213 30389 20216
rect 30423 20213 30435 20247
rect 30377 20207 30435 20213
rect 552 20154 31648 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 12096 20154
rect 12148 20102 12160 20154
rect 12212 20102 12224 20154
rect 12276 20102 12288 20154
rect 12340 20102 12352 20154
rect 12404 20102 19870 20154
rect 19922 20102 19934 20154
rect 19986 20102 19998 20154
rect 20050 20102 20062 20154
rect 20114 20102 20126 20154
rect 20178 20102 27644 20154
rect 27696 20102 27708 20154
rect 27760 20102 27772 20154
rect 27824 20102 27836 20154
rect 27888 20102 27900 20154
rect 27952 20102 31648 20154
rect 552 20080 31648 20102
rect 2314 20000 2320 20052
rect 2372 20000 2378 20052
rect 2685 20043 2743 20049
rect 2685 20009 2697 20043
rect 2731 20040 2743 20043
rect 2774 20040 2780 20052
rect 2731 20012 2780 20040
rect 2731 20009 2743 20012
rect 2685 20003 2743 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 2961 20043 3019 20049
rect 2961 20009 2973 20043
rect 3007 20040 3019 20043
rect 3050 20040 3056 20052
rect 3007 20012 3056 20040
rect 3007 20009 3019 20012
rect 2961 20003 3019 20009
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3142 20000 3148 20052
rect 3200 20040 3206 20052
rect 3200 20012 5396 20040
rect 3200 20000 3206 20012
rect 2866 19972 2872 19984
rect 2516 19944 2872 19972
rect 2038 19864 2044 19916
rect 2096 19864 2102 19916
rect 2516 19913 2544 19944
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 4798 19972 4804 19984
rect 3068 19944 4804 19972
rect 3068 19913 3096 19944
rect 4798 19932 4804 19944
rect 4856 19932 4862 19984
rect 5368 19972 5396 20012
rect 5442 20000 5448 20052
rect 5500 20000 5506 20052
rect 5813 20043 5871 20049
rect 5813 20009 5825 20043
rect 5859 20040 5871 20043
rect 5902 20040 5908 20052
rect 5859 20012 5908 20040
rect 5859 20009 5871 20012
rect 5813 20003 5871 20009
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 6549 20043 6607 20049
rect 6042 20012 6500 20040
rect 6042 19972 6070 20012
rect 5368 19944 6070 19972
rect 2225 19907 2283 19913
rect 2225 19873 2237 19907
rect 2271 19904 2283 19907
rect 2501 19907 2559 19913
rect 2271 19876 2452 19904
rect 2271 19873 2283 19876
rect 2225 19867 2283 19873
rect 2130 19660 2136 19712
rect 2188 19660 2194 19712
rect 2424 19700 2452 19876
rect 2501 19873 2513 19907
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19873 2835 19907
rect 2777 19867 2835 19873
rect 3053 19907 3111 19913
rect 3053 19873 3065 19907
rect 3099 19873 3111 19907
rect 3053 19867 3111 19873
rect 3329 19907 3387 19913
rect 3329 19873 3341 19907
rect 3375 19904 3387 19907
rect 3510 19904 3516 19916
rect 3375 19876 3516 19904
rect 3375 19873 3387 19876
rect 3329 19867 3387 19873
rect 2792 19768 2820 19867
rect 3510 19864 3516 19876
rect 3568 19864 3574 19916
rect 3878 19864 3884 19916
rect 3936 19864 3942 19916
rect 3970 19864 3976 19916
rect 4028 19864 4034 19916
rect 4890 19864 4896 19916
rect 4948 19864 4954 19916
rect 5350 19864 5356 19916
rect 5408 19864 5414 19916
rect 5810 19864 5816 19916
rect 5868 19904 5874 19916
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5868 19876 6009 19904
rect 5868 19864 5874 19876
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 5997 19867 6055 19873
rect 6086 19864 6092 19916
rect 6144 19864 6150 19916
rect 6270 19864 6276 19916
rect 6328 19864 6334 19916
rect 6365 19907 6423 19913
rect 6365 19873 6377 19907
rect 6411 19873 6423 19907
rect 6472 19904 6500 20012
rect 6549 20009 6561 20043
rect 6595 20040 6607 20043
rect 7006 20040 7012 20052
rect 6595 20012 7012 20040
rect 6595 20009 6607 20012
rect 6549 20003 6607 20009
rect 7006 20000 7012 20012
rect 7064 20000 7070 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 10965 20043 11023 20049
rect 10965 20040 10977 20043
rect 9732 20012 10977 20040
rect 9732 20000 9738 20012
rect 10965 20009 10977 20012
rect 11011 20009 11023 20043
rect 10965 20003 11023 20009
rect 13817 20043 13875 20049
rect 13817 20009 13829 20043
rect 13863 20040 13875 20043
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 13863 20012 14565 20040
rect 13863 20009 13875 20012
rect 13817 20003 13875 20009
rect 14553 20009 14565 20012
rect 14599 20040 14611 20043
rect 14642 20040 14648 20052
rect 14599 20012 14648 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 18046 20040 18052 20052
rect 15396 20012 18052 20040
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 14461 19975 14519 19981
rect 8904 19944 12388 19972
rect 8904 19932 8910 19944
rect 6641 19907 6699 19913
rect 6641 19904 6653 19907
rect 6472 19876 6653 19904
rect 6365 19867 6423 19873
rect 6641 19873 6653 19876
rect 6687 19904 6699 19907
rect 6687 19876 9076 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 3142 19836 3148 19848
rect 3007 19808 3148 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 3988 19768 4016 19864
rect 6380 19836 6408 19867
rect 7006 19836 7012 19848
rect 6380 19808 7012 19836
rect 7006 19796 7012 19808
rect 7064 19796 7070 19848
rect 8018 19768 8024 19780
rect 2792 19740 3280 19768
rect 3988 19740 8024 19768
rect 3252 19712 3280 19740
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 3142 19700 3148 19712
rect 2424 19672 3148 19700
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 3234 19660 3240 19712
rect 3292 19660 3298 19712
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 3605 19703 3663 19709
rect 3605 19700 3617 19703
rect 3568 19672 3617 19700
rect 3568 19660 3574 19672
rect 3605 19669 3617 19672
rect 3651 19669 3663 19703
rect 3605 19663 3663 19669
rect 3973 19703 4031 19709
rect 3973 19669 3985 19703
rect 4019 19700 4031 19703
rect 4154 19700 4160 19712
rect 4019 19672 4160 19700
rect 4019 19669 4031 19672
rect 3973 19663 4031 19669
rect 4154 19660 4160 19672
rect 4212 19660 4218 19712
rect 4801 19703 4859 19709
rect 4801 19669 4813 19703
rect 4847 19700 4859 19703
rect 5074 19700 5080 19712
rect 4847 19672 5080 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 5074 19660 5080 19672
rect 5132 19660 5138 19712
rect 9048 19700 9076 19876
rect 9122 19864 9128 19916
rect 9180 19864 9186 19916
rect 9392 19907 9450 19913
rect 9392 19873 9404 19907
rect 9438 19904 9450 19907
rect 9858 19904 9864 19916
rect 9438 19876 9864 19904
rect 9438 19873 9450 19876
rect 9392 19867 9450 19873
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 11974 19864 11980 19916
rect 12032 19904 12038 19916
rect 12253 19907 12311 19913
rect 12253 19904 12265 19907
rect 12032 19876 12265 19904
rect 12032 19864 12038 19876
rect 12253 19873 12265 19876
rect 12299 19873 12311 19907
rect 12253 19867 12311 19873
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19805 11575 19839
rect 12360 19836 12388 19944
rect 14461 19941 14473 19975
rect 14507 19972 14519 19975
rect 15194 19972 15200 19984
rect 14507 19944 15200 19972
rect 14507 19941 14519 19944
rect 14461 19935 14519 19941
rect 15194 19932 15200 19944
rect 15252 19932 15258 19984
rect 12526 19864 12532 19916
rect 12584 19864 12590 19916
rect 14826 19904 14832 19916
rect 14660 19876 14832 19904
rect 14660 19836 14688 19876
rect 14826 19864 14832 19876
rect 14884 19904 14890 19916
rect 14921 19907 14979 19913
rect 14921 19904 14933 19907
rect 14884 19876 14933 19904
rect 14884 19864 14890 19876
rect 14921 19873 14933 19876
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 15105 19907 15163 19913
rect 15105 19873 15117 19907
rect 15151 19904 15163 19907
rect 15396 19904 15424 20012
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 19061 20043 19119 20049
rect 19061 20040 19073 20043
rect 18196 20012 19073 20040
rect 18196 20000 18202 20012
rect 19061 20009 19073 20012
rect 19107 20009 19119 20043
rect 19061 20003 19119 20009
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 20622 20040 20628 20052
rect 19392 20012 20628 20040
rect 19392 20000 19398 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 20714 20000 20720 20052
rect 20772 20040 20778 20052
rect 20901 20043 20959 20049
rect 20901 20040 20913 20043
rect 20772 20012 20913 20040
rect 20772 20000 20778 20012
rect 20901 20009 20913 20012
rect 20947 20009 20959 20043
rect 20901 20003 20959 20009
rect 21266 20000 21272 20052
rect 21324 20000 21330 20052
rect 21910 20000 21916 20052
rect 21968 20040 21974 20052
rect 22005 20043 22063 20049
rect 22005 20040 22017 20043
rect 21968 20012 22017 20040
rect 21968 20000 21974 20012
rect 22005 20009 22017 20012
rect 22051 20009 22063 20043
rect 22005 20003 22063 20009
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22373 20043 22431 20049
rect 22373 20040 22385 20043
rect 22152 20012 22385 20040
rect 22152 20000 22158 20012
rect 22373 20009 22385 20012
rect 22419 20040 22431 20043
rect 22462 20040 22468 20052
rect 22419 20012 22468 20040
rect 22419 20009 22431 20012
rect 22373 20003 22431 20009
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 26326 20040 26332 20052
rect 25148 20012 26332 20040
rect 19429 19975 19487 19981
rect 19429 19972 19441 19975
rect 16132 19944 16896 19972
rect 15151 19876 15424 19904
rect 15151 19873 15163 19876
rect 15105 19867 15163 19873
rect 15470 19864 15476 19916
rect 15528 19864 15534 19916
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 16132 19913 16160 19944
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15620 19876 15853 19904
rect 15620 19864 15626 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 16117 19907 16175 19913
rect 16117 19873 16129 19907
rect 16163 19873 16175 19907
rect 16117 19867 16175 19873
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19873 16267 19907
rect 16209 19867 16267 19873
rect 12360 19808 14688 19836
rect 14737 19839 14795 19845
rect 11517 19799 11575 19805
rect 14737 19805 14749 19839
rect 14783 19836 14795 19839
rect 15013 19839 15071 19845
rect 15013 19836 15025 19839
rect 14783 19808 15025 19836
rect 14783 19805 14795 19808
rect 14737 19799 14795 19805
rect 15013 19805 15025 19808
rect 15059 19805 15071 19839
rect 16224 19836 16252 19867
rect 16298 19864 16304 19916
rect 16356 19904 16362 19916
rect 16868 19913 16896 19944
rect 18800 19944 19441 19972
rect 18800 19916 18828 19944
rect 19429 19941 19441 19944
rect 19475 19941 19487 19975
rect 22922 19972 22928 19984
rect 19429 19935 19487 19941
rect 21744 19944 22928 19972
rect 16393 19907 16451 19913
rect 16393 19904 16405 19907
rect 16356 19876 16405 19904
rect 16356 19864 16362 19876
rect 16393 19873 16405 19876
rect 16439 19873 16451 19907
rect 16393 19867 16451 19873
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 16853 19907 16911 19913
rect 16853 19873 16865 19907
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 16684 19836 16712 19867
rect 16868 19836 16896 19867
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 18012 19876 18705 19904
rect 18012 19864 18018 19876
rect 18693 19873 18705 19876
rect 18739 19904 18751 19907
rect 18782 19904 18788 19916
rect 18739 19876 18788 19904
rect 18739 19873 18751 19876
rect 18693 19867 18751 19873
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 18969 19907 19027 19913
rect 18969 19873 18981 19907
rect 19015 19904 19027 19907
rect 19058 19904 19064 19916
rect 19015 19876 19064 19904
rect 19015 19873 19027 19876
rect 18969 19867 19027 19873
rect 18892 19836 18920 19867
rect 19058 19864 19064 19876
rect 19116 19864 19122 19916
rect 19245 19907 19303 19913
rect 19245 19873 19257 19907
rect 19291 19904 19303 19907
rect 19334 19904 19340 19916
rect 19291 19876 19340 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19873 19579 19907
rect 19521 19867 19579 19873
rect 19536 19836 19564 19867
rect 19610 19864 19616 19916
rect 19668 19864 19674 19916
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 20438 19836 20444 19848
rect 15013 19799 15071 19805
rect 15212 19808 16804 19836
rect 16868 19808 20444 19836
rect 10505 19771 10563 19777
rect 10505 19737 10517 19771
rect 10551 19768 10563 19771
rect 11238 19768 11244 19780
rect 10551 19740 11244 19768
rect 10551 19737 10563 19740
rect 10505 19731 10563 19737
rect 11238 19728 11244 19740
rect 11296 19768 11302 19780
rect 11532 19768 11560 19799
rect 11296 19740 11560 19768
rect 11296 19728 11302 19740
rect 14274 19728 14280 19780
rect 14332 19768 14338 19780
rect 15212 19768 15240 19808
rect 14332 19740 15240 19768
rect 14332 19728 14338 19740
rect 15286 19728 15292 19780
rect 15344 19768 15350 19780
rect 16022 19768 16028 19780
rect 15344 19740 16028 19768
rect 15344 19728 15350 19740
rect 16022 19728 16028 19740
rect 16080 19728 16086 19780
rect 16776 19768 16804 19808
rect 18708 19780 18736 19808
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 20916 19836 20944 19867
rect 21082 19864 21088 19916
rect 21140 19864 21146 19916
rect 21174 19864 21180 19916
rect 21232 19904 21238 19916
rect 21545 19907 21603 19913
rect 21545 19904 21557 19907
rect 21232 19876 21557 19904
rect 21232 19864 21238 19876
rect 21545 19873 21557 19876
rect 21591 19873 21603 19907
rect 21545 19867 21603 19873
rect 21634 19864 21640 19916
rect 21692 19864 21698 19916
rect 21744 19913 21772 19944
rect 22922 19932 22928 19944
rect 22980 19932 22986 19984
rect 21729 19907 21787 19913
rect 21729 19873 21741 19907
rect 21775 19873 21787 19907
rect 21729 19867 21787 19873
rect 21818 19864 21824 19916
rect 21876 19904 21882 19916
rect 21913 19907 21971 19913
rect 21913 19904 21925 19907
rect 21876 19876 21925 19904
rect 21876 19864 21882 19876
rect 21913 19873 21925 19876
rect 21959 19873 21971 19907
rect 21913 19867 21971 19873
rect 22186 19864 22192 19916
rect 22244 19864 22250 19916
rect 22465 19907 22523 19913
rect 22465 19873 22477 19907
rect 22511 19904 22523 19907
rect 23382 19904 23388 19916
rect 22511 19876 23388 19904
rect 22511 19873 22523 19876
rect 22465 19867 22523 19873
rect 22094 19836 22100 19848
rect 20916 19808 22100 19836
rect 16850 19768 16856 19780
rect 16776 19740 16856 19768
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 18690 19728 18696 19780
rect 18748 19728 18754 19780
rect 18874 19728 18880 19780
rect 18932 19768 18938 19780
rect 19794 19768 19800 19780
rect 18932 19740 19800 19768
rect 18932 19728 18938 19740
rect 19794 19728 19800 19740
rect 19852 19768 19858 19780
rect 20916 19768 20944 19808
rect 22094 19796 22100 19808
rect 22152 19796 22158 19848
rect 19852 19740 20944 19768
rect 19852 19728 19858 19740
rect 21082 19728 21088 19780
rect 21140 19768 21146 19780
rect 22480 19768 22508 19867
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 24854 19864 24860 19916
rect 24912 19864 24918 19916
rect 24946 19864 24952 19916
rect 25004 19864 25010 19916
rect 25148 19913 25176 20012
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 26421 20043 26479 20049
rect 26421 20009 26433 20043
rect 26467 20009 26479 20043
rect 26421 20003 26479 20009
rect 25498 19932 25504 19984
rect 25556 19972 25562 19984
rect 25556 19944 26096 19972
rect 25556 19932 25562 19944
rect 25133 19907 25191 19913
rect 25133 19873 25145 19907
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 21140 19740 22508 19768
rect 21140 19728 21146 19740
rect 10870 19700 10876 19712
rect 9048 19672 10876 19700
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 14090 19660 14096 19712
rect 14148 19660 14154 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 15749 19703 15807 19709
rect 15749 19700 15761 19703
rect 15528 19672 15761 19700
rect 15528 19660 15534 19672
rect 15749 19669 15761 19672
rect 15795 19700 15807 19703
rect 16482 19700 16488 19712
rect 15795 19672 16488 19700
rect 15795 19669 15807 19672
rect 15749 19663 15807 19669
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 16574 19660 16580 19712
rect 16632 19660 16638 19712
rect 16758 19660 16764 19712
rect 16816 19660 16822 19712
rect 18046 19660 18052 19712
rect 18104 19700 18110 19712
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 18104 19672 18521 19700
rect 18104 19660 18110 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 18509 19663 18567 19669
rect 19702 19660 19708 19712
rect 19760 19660 19766 19712
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 25148 19700 25176 19867
rect 25222 19864 25228 19916
rect 25280 19864 25286 19916
rect 25314 19864 25320 19916
rect 25372 19864 25378 19916
rect 25406 19864 25412 19916
rect 25464 19904 25470 19916
rect 25777 19907 25835 19913
rect 25777 19904 25789 19907
rect 25464 19876 25789 19904
rect 25464 19864 25470 19876
rect 25777 19873 25789 19876
rect 25823 19873 25835 19907
rect 25777 19867 25835 19873
rect 25869 19907 25927 19913
rect 25869 19873 25881 19907
rect 25915 19904 25927 19907
rect 25958 19904 25964 19916
rect 25915 19876 25964 19904
rect 25915 19873 25927 19876
rect 25869 19867 25927 19873
rect 25792 19836 25820 19867
rect 25958 19864 25964 19876
rect 26016 19864 26022 19916
rect 26068 19913 26096 19944
rect 26053 19907 26111 19913
rect 26053 19873 26065 19907
rect 26099 19873 26111 19907
rect 26053 19867 26111 19873
rect 26145 19907 26203 19913
rect 26145 19873 26157 19907
rect 26191 19904 26203 19907
rect 26436 19904 26464 20003
rect 26602 20000 26608 20052
rect 26660 20040 26666 20052
rect 28077 20043 28135 20049
rect 26660 20012 27016 20040
rect 26660 20000 26666 20012
rect 26694 19932 26700 19984
rect 26752 19932 26758 19984
rect 26191 19876 26464 19904
rect 26191 19873 26203 19876
rect 26145 19867 26203 19873
rect 26510 19864 26516 19916
rect 26568 19904 26574 19916
rect 26605 19907 26663 19913
rect 26605 19904 26617 19907
rect 26568 19876 26617 19904
rect 26568 19864 26574 19876
rect 26605 19873 26617 19876
rect 26651 19873 26663 19907
rect 26605 19867 26663 19873
rect 26620 19836 26648 19867
rect 26786 19864 26792 19916
rect 26844 19864 26850 19916
rect 26988 19913 27016 20012
rect 28077 20009 28089 20043
rect 28123 20040 28135 20043
rect 28350 20040 28356 20052
rect 28123 20012 28356 20040
rect 28123 20009 28135 20012
rect 28077 20003 28135 20009
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 29086 19932 29092 19984
rect 29144 19932 29150 19984
rect 30098 19932 30104 19984
rect 30156 19932 30162 19984
rect 26973 19907 27031 19913
rect 26973 19873 26985 19907
rect 27019 19873 27031 19907
rect 26973 19867 27031 19873
rect 27801 19907 27859 19913
rect 27801 19873 27813 19907
rect 27847 19904 27859 19907
rect 27982 19904 27988 19916
rect 27847 19876 27988 19904
rect 27847 19873 27859 19876
rect 27801 19867 27859 19873
rect 27982 19864 27988 19876
rect 28040 19864 28046 19916
rect 28166 19864 28172 19916
rect 28224 19864 28230 19916
rect 28951 19907 29009 19913
rect 28951 19873 28963 19907
rect 28997 19873 29009 19907
rect 28951 19867 29009 19873
rect 29181 19907 29239 19913
rect 29181 19873 29193 19907
rect 29227 19873 29239 19907
rect 29362 19904 29368 19916
rect 29323 19876 29368 19904
rect 29181 19867 29239 19873
rect 28966 19836 28994 19867
rect 25792 19808 25896 19836
rect 26620 19808 28994 19836
rect 25498 19728 25504 19780
rect 25556 19728 25562 19780
rect 25868 19768 25896 19808
rect 29196 19768 29224 19867
rect 29362 19864 29368 19876
rect 29420 19864 29426 19916
rect 29454 19864 29460 19916
rect 29512 19864 29518 19916
rect 29730 19864 29736 19916
rect 29788 19904 29794 19916
rect 29917 19907 29975 19913
rect 29917 19904 29929 19907
rect 29788 19876 29929 19904
rect 29788 19864 29794 19876
rect 29917 19873 29929 19876
rect 29963 19873 29975 19907
rect 29917 19867 29975 19873
rect 25868 19740 29224 19768
rect 20404 19672 25176 19700
rect 20404 19660 20410 19672
rect 25590 19660 25596 19712
rect 25648 19660 25654 19712
rect 26234 19660 26240 19712
rect 26292 19700 26298 19712
rect 27433 19703 27491 19709
rect 27433 19700 27445 19703
rect 26292 19672 27445 19700
rect 26292 19660 26298 19672
rect 27433 19669 27445 19672
rect 27479 19669 27491 19703
rect 27433 19663 27491 19669
rect 27706 19660 27712 19712
rect 27764 19660 27770 19712
rect 27893 19703 27951 19709
rect 27893 19669 27905 19703
rect 27939 19700 27951 19703
rect 28813 19703 28871 19709
rect 28813 19700 28825 19703
rect 27939 19672 28825 19700
rect 27939 19669 27951 19672
rect 27893 19663 27951 19669
rect 28813 19669 28825 19672
rect 28859 19669 28871 19703
rect 28813 19663 28871 19669
rect 29086 19660 29092 19712
rect 29144 19700 29150 19712
rect 29641 19703 29699 19709
rect 29641 19700 29653 19703
rect 29144 19672 29653 19700
rect 29144 19660 29150 19672
rect 29641 19669 29653 19672
rect 29687 19700 29699 19703
rect 30190 19700 30196 19712
rect 29687 19672 30196 19700
rect 29687 19669 29699 19672
rect 29641 19663 29699 19669
rect 30190 19660 30196 19672
rect 30248 19660 30254 19712
rect 552 19610 31648 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 11436 19610
rect 11488 19558 11500 19610
rect 11552 19558 11564 19610
rect 11616 19558 11628 19610
rect 11680 19558 11692 19610
rect 11744 19558 19210 19610
rect 19262 19558 19274 19610
rect 19326 19558 19338 19610
rect 19390 19558 19402 19610
rect 19454 19558 19466 19610
rect 19518 19558 26984 19610
rect 27036 19558 27048 19610
rect 27100 19558 27112 19610
rect 27164 19558 27176 19610
rect 27228 19558 27240 19610
rect 27292 19558 31648 19610
rect 552 19536 31648 19558
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 4062 19496 4068 19508
rect 3292 19468 4068 19496
rect 3292 19456 3298 19468
rect 4062 19456 4068 19468
rect 4120 19496 4126 19508
rect 4617 19499 4675 19505
rect 4617 19496 4629 19499
rect 4120 19468 4629 19496
rect 4120 19456 4126 19468
rect 4617 19465 4629 19468
rect 4663 19465 4675 19499
rect 4617 19459 4675 19465
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 9582 19496 9588 19508
rect 7616 19468 9588 19496
rect 7616 19456 7622 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 9950 19456 9956 19508
rect 10008 19456 10014 19508
rect 11974 19456 11980 19508
rect 12032 19496 12038 19508
rect 14274 19496 14280 19508
rect 12032 19468 14280 19496
rect 12032 19456 12038 19468
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 16298 19456 16304 19508
rect 16356 19456 16362 19508
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 17034 19496 17040 19508
rect 16632 19468 17040 19496
rect 16632 19456 16638 19468
rect 17034 19456 17040 19468
rect 17092 19456 17098 19508
rect 18782 19456 18788 19508
rect 18840 19456 18846 19508
rect 20530 19496 20536 19508
rect 18892 19468 20536 19496
rect 2038 19388 2044 19440
rect 2096 19428 2102 19440
rect 4341 19431 4399 19437
rect 4341 19428 4353 19431
rect 2096 19400 4353 19428
rect 2096 19388 2102 19400
rect 4341 19397 4353 19400
rect 4387 19428 4399 19431
rect 4706 19428 4712 19440
rect 4387 19400 4712 19428
rect 4387 19397 4399 19400
rect 4341 19391 4399 19397
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 7837 19431 7895 19437
rect 7837 19397 7849 19431
rect 7883 19428 7895 19431
rect 7926 19428 7932 19440
rect 7883 19400 7932 19428
rect 7883 19397 7895 19400
rect 7837 19391 7895 19397
rect 7926 19388 7932 19400
rect 7984 19388 7990 19440
rect 8404 19400 9536 19428
rect 3326 19360 3332 19372
rect 2884 19332 3332 19360
rect 1394 19252 1400 19304
rect 1452 19292 1458 19304
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 1452 19264 1869 19292
rect 1452 19252 1458 19264
rect 1857 19261 1869 19264
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 2130 19252 2136 19304
rect 2188 19292 2194 19304
rect 2884 19301 2912 19332
rect 3326 19320 3332 19332
rect 3384 19360 3390 19372
rect 4062 19360 4068 19372
rect 3384 19332 4068 19360
rect 3384 19320 3390 19332
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 5074 19360 5080 19372
rect 4448 19332 5080 19360
rect 2685 19295 2743 19301
rect 2685 19292 2697 19295
rect 2188 19264 2697 19292
rect 2188 19252 2194 19264
rect 2685 19261 2697 19264
rect 2731 19261 2743 19295
rect 2685 19255 2743 19261
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19261 2927 19295
rect 2869 19255 2927 19261
rect 2958 19252 2964 19304
rect 3016 19252 3022 19304
rect 3234 19252 3240 19304
rect 3292 19252 3298 19304
rect 4448 19301 4476 19332
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 7576 19332 7788 19360
rect 4439 19295 4497 19301
rect 4439 19261 4451 19295
rect 4485 19261 4497 19295
rect 4439 19255 4497 19261
rect 4617 19295 4675 19301
rect 4617 19261 4629 19295
rect 4663 19292 4675 19295
rect 5718 19292 5724 19304
rect 4663 19264 5724 19292
rect 4663 19261 4675 19264
rect 4617 19255 4675 19261
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 7576 19292 7604 19332
rect 6840 19264 7604 19292
rect 7653 19295 7711 19301
rect 2498 19184 2504 19236
rect 2556 19184 2562 19236
rect 2976 19224 3004 19252
rect 3973 19227 4031 19233
rect 3973 19224 3985 19227
rect 2976 19196 3985 19224
rect 3973 19193 3985 19196
rect 4019 19193 4031 19227
rect 3973 19187 4031 19193
rect 4062 19184 4068 19236
rect 4120 19224 4126 19236
rect 4157 19227 4215 19233
rect 4157 19224 4169 19227
rect 4120 19196 4169 19224
rect 4120 19184 4126 19196
rect 4157 19193 4169 19196
rect 4203 19224 4215 19227
rect 6840 19224 6868 19264
rect 7653 19261 7665 19295
rect 7699 19261 7711 19295
rect 7653 19255 7711 19261
rect 4203 19196 6868 19224
rect 4203 19193 4215 19196
rect 4157 19187 4215 19193
rect 6914 19184 6920 19236
rect 6972 19224 6978 19236
rect 7668 19224 7696 19255
rect 7760 19236 7788 19332
rect 8404 19304 8432 19400
rect 9508 19369 9536 19400
rect 15838 19388 15844 19440
rect 15896 19428 15902 19440
rect 16316 19428 16344 19456
rect 15896 19400 16252 19428
rect 16316 19400 17080 19428
rect 15896 19388 15902 19400
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 8527 19332 9413 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 10244 19332 10548 19360
rect 8018 19292 8024 19304
rect 7944 19264 8024 19292
rect 6972 19196 7696 19224
rect 6972 19184 6978 19196
rect 1578 19116 1584 19168
rect 1636 19156 1642 19168
rect 1765 19159 1823 19165
rect 1765 19156 1777 19159
rect 1636 19128 1777 19156
rect 1636 19116 1642 19128
rect 1765 19125 1777 19128
rect 1811 19125 1823 19159
rect 1765 19119 1823 19125
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 3881 19159 3939 19165
rect 3881 19156 3893 19159
rect 3384 19128 3893 19156
rect 3384 19116 3390 19128
rect 3881 19125 3893 19128
rect 3927 19125 3939 19159
rect 3881 19119 3939 19125
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 7558 19156 7564 19168
rect 4856 19128 7564 19156
rect 4856 19116 4862 19128
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 7668 19156 7696 19196
rect 7742 19184 7748 19236
rect 7800 19184 7806 19236
rect 7944 19233 7972 19264
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 8386 19252 8392 19304
rect 8444 19252 8450 19304
rect 8570 19252 8576 19304
rect 8628 19252 8634 19304
rect 8662 19252 8668 19304
rect 8720 19292 8726 19304
rect 9033 19295 9091 19301
rect 9033 19294 9045 19295
rect 8864 19292 9045 19294
rect 8720 19266 9045 19292
rect 8720 19264 8892 19266
rect 8720 19252 8726 19264
rect 9033 19261 9045 19266
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9214 19292 9220 19304
rect 9171 19264 9220 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 9306 19252 9312 19304
rect 9364 19252 9370 19304
rect 9674 19252 9680 19304
rect 9732 19252 9738 19304
rect 9858 19252 9864 19304
rect 9916 19252 9922 19304
rect 10244 19301 10272 19332
rect 10229 19295 10287 19301
rect 10229 19261 10241 19295
rect 10275 19261 10287 19295
rect 10229 19255 10287 19261
rect 10318 19252 10324 19304
rect 10376 19252 10382 19304
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19261 10471 19295
rect 10413 19255 10471 19261
rect 7929 19227 7987 19233
rect 7929 19193 7941 19227
rect 7975 19193 7987 19227
rect 8849 19227 8907 19233
rect 8849 19224 8861 19227
rect 7929 19187 7987 19193
rect 8266 19196 8861 19224
rect 8266 19156 8294 19196
rect 8849 19193 8861 19196
rect 8895 19224 8907 19227
rect 8938 19224 8944 19236
rect 8895 19196 8944 19224
rect 8895 19193 8907 19196
rect 8849 19187 8907 19193
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 10428 19224 10456 19255
rect 10520 19236 10548 19332
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 14185 19363 14243 19369
rect 14185 19360 14197 19363
rect 14148 19332 14197 19360
rect 14148 19320 14154 19332
rect 14185 19329 14197 19332
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19360 14427 19363
rect 14918 19360 14924 19372
rect 14415 19332 14924 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 14918 19320 14924 19332
rect 14976 19360 14982 19372
rect 15930 19360 15936 19372
rect 14976 19332 15936 19360
rect 14976 19320 14982 19332
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 10594 19252 10600 19304
rect 10652 19252 10658 19304
rect 10686 19252 10692 19304
rect 10744 19252 10750 19304
rect 14734 19252 14740 19304
rect 14792 19252 14798 19304
rect 15010 19252 15016 19304
rect 15068 19252 15074 19304
rect 16224 19292 16252 19400
rect 16761 19363 16819 19369
rect 16761 19329 16773 19363
rect 16807 19360 16819 19363
rect 16942 19360 16948 19372
rect 16807 19332 16948 19360
rect 16807 19329 16819 19332
rect 16761 19323 16819 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 16298 19292 16304 19304
rect 16224 19264 16304 19292
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 10244 19196 10456 19224
rect 7668 19128 8294 19156
rect 8665 19159 8723 19165
rect 8665 19125 8677 19159
rect 8711 19156 8723 19159
rect 10244 19156 10272 19196
rect 10502 19184 10508 19236
rect 10560 19224 10566 19236
rect 10781 19227 10839 19233
rect 10781 19224 10793 19227
rect 10560 19196 10793 19224
rect 10560 19184 10566 19196
rect 10781 19193 10793 19196
rect 10827 19193 10839 19227
rect 10781 19187 10839 19193
rect 13906 19184 13912 19236
rect 13964 19224 13970 19236
rect 14093 19227 14151 19233
rect 14093 19224 14105 19227
rect 13964 19196 14105 19224
rect 13964 19184 13970 19196
rect 14093 19193 14105 19196
rect 14139 19193 14151 19227
rect 14093 19187 14151 19193
rect 16022 19184 16028 19236
rect 16080 19224 16086 19236
rect 16500 19224 16528 19255
rect 16666 19252 16672 19304
rect 16724 19252 16730 19304
rect 17052 19301 17080 19400
rect 17494 19320 17500 19372
rect 17552 19360 17558 19372
rect 18892 19360 18920 19468
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 21453 19499 21511 19505
rect 21453 19465 21465 19499
rect 21499 19496 21511 19499
rect 21634 19496 21640 19508
rect 21499 19468 21640 19496
rect 21499 19465 21511 19468
rect 21453 19459 21511 19465
rect 21634 19456 21640 19468
rect 21692 19456 21698 19508
rect 25590 19456 25596 19508
rect 25648 19496 25654 19508
rect 25869 19499 25927 19505
rect 25869 19496 25881 19499
rect 25648 19468 25881 19496
rect 25648 19456 25654 19468
rect 25869 19465 25881 19468
rect 25915 19465 25927 19499
rect 25869 19459 25927 19465
rect 25958 19456 25964 19508
rect 26016 19496 26022 19508
rect 26786 19496 26792 19508
rect 26016 19468 26792 19496
rect 26016 19456 26022 19468
rect 26786 19456 26792 19468
rect 26844 19496 26850 19508
rect 27985 19499 28043 19505
rect 27985 19496 27997 19499
rect 26844 19468 27997 19496
rect 26844 19456 26850 19468
rect 27985 19465 27997 19468
rect 28031 19496 28043 19499
rect 28166 19496 28172 19508
rect 28031 19468 28172 19496
rect 28031 19465 28043 19468
rect 27985 19459 28043 19465
rect 28166 19456 28172 19468
rect 28224 19456 28230 19508
rect 20438 19388 20444 19440
rect 20496 19428 20502 19440
rect 20496 19400 24808 19428
rect 20496 19388 20502 19400
rect 17552 19332 18920 19360
rect 17552 19320 17558 19332
rect 17880 19301 17908 19332
rect 19702 19320 19708 19372
rect 19760 19360 19766 19372
rect 20349 19363 20407 19369
rect 20349 19360 20361 19363
rect 19760 19332 20361 19360
rect 19760 19320 19766 19332
rect 20349 19329 20361 19332
rect 20395 19329 20407 19363
rect 20349 19323 20407 19329
rect 20622 19320 20628 19372
rect 20680 19360 20686 19372
rect 24780 19360 24808 19400
rect 24854 19388 24860 19440
rect 24912 19428 24918 19440
rect 27706 19428 27712 19440
rect 24912 19400 27712 19428
rect 24912 19388 24918 19400
rect 27706 19388 27712 19400
rect 27764 19388 27770 19440
rect 28077 19431 28135 19437
rect 28077 19397 28089 19431
rect 28123 19428 28135 19431
rect 29178 19428 29184 19440
rect 28123 19400 29184 19428
rect 28123 19397 28135 19400
rect 28077 19391 28135 19397
rect 20680 19332 22094 19360
rect 24780 19332 25820 19360
rect 20680 19320 20686 19332
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 17037 19295 17095 19301
rect 17037 19261 17049 19295
rect 17083 19261 17095 19295
rect 17037 19255 17095 19261
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19261 17923 19295
rect 17865 19255 17923 19261
rect 16080 19196 16528 19224
rect 16080 19184 16086 19196
rect 8711 19128 10272 19156
rect 13725 19159 13783 19165
rect 8711 19125 8723 19128
rect 8665 19119 8723 19125
rect 13725 19125 13737 19159
rect 13771 19156 13783 19159
rect 13998 19156 14004 19168
rect 13771 19128 14004 19156
rect 13771 19125 13783 19128
rect 13725 19119 13783 19125
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 15654 19116 15660 19168
rect 15712 19156 15718 19168
rect 16868 19156 16896 19255
rect 18046 19252 18052 19304
rect 18104 19252 18110 19304
rect 18138 19252 18144 19304
rect 18196 19252 18202 19304
rect 18233 19295 18291 19301
rect 18233 19261 18245 19295
rect 18279 19292 18291 19295
rect 18322 19292 18328 19304
rect 18279 19264 18328 19292
rect 18279 19261 18291 19264
rect 18233 19255 18291 19261
rect 17218 19184 17224 19236
rect 17276 19184 17282 19236
rect 17310 19184 17316 19236
rect 17368 19224 17374 19236
rect 18248 19224 18276 19255
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 18524 19264 20085 19292
rect 18524 19233 18552 19264
rect 20073 19261 20085 19264
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21361 19295 21419 19301
rect 21361 19292 21373 19295
rect 21140 19264 21373 19292
rect 21140 19252 21146 19264
rect 21361 19261 21373 19264
rect 21407 19261 21419 19295
rect 21361 19255 21419 19261
rect 21542 19252 21548 19304
rect 21600 19252 21606 19304
rect 22066 19292 22094 19332
rect 24213 19295 24271 19301
rect 24213 19292 24225 19295
rect 22066 19264 24225 19292
rect 24213 19261 24225 19264
rect 24259 19292 24271 19295
rect 25682 19292 25688 19304
rect 24259 19264 25688 19292
rect 24259 19261 24271 19264
rect 24213 19255 24271 19261
rect 25682 19252 25688 19264
rect 25740 19252 25746 19304
rect 25792 19292 25820 19332
rect 25866 19320 25872 19372
rect 25924 19360 25930 19372
rect 25924 19332 26234 19360
rect 25924 19320 25930 19332
rect 25958 19292 25964 19304
rect 25792 19264 25964 19292
rect 25958 19252 25964 19264
rect 26016 19252 26022 19304
rect 26206 19292 26234 19332
rect 26326 19320 26332 19372
rect 26384 19360 26390 19372
rect 28092 19360 28120 19391
rect 29178 19388 29184 19400
rect 29236 19388 29242 19440
rect 26384 19332 28120 19360
rect 26384 19320 26390 19332
rect 26697 19295 26755 19301
rect 26697 19292 26709 19295
rect 26206 19264 26709 19292
rect 26697 19261 26709 19264
rect 26743 19292 26755 19295
rect 27338 19292 27344 19304
rect 26743 19264 27344 19292
rect 26743 19261 26755 19264
rect 26697 19255 26755 19261
rect 27338 19252 27344 19264
rect 27396 19292 27402 19304
rect 28629 19295 28687 19301
rect 28629 19292 28641 19295
rect 27396 19264 28641 19292
rect 27396 19252 27402 19264
rect 28629 19261 28641 19264
rect 28675 19292 28687 19295
rect 28994 19292 29000 19304
rect 28675 19264 29000 19292
rect 28675 19261 28687 19264
rect 28629 19255 28687 19261
rect 28994 19252 29000 19264
rect 29052 19252 29058 19304
rect 29273 19295 29331 19301
rect 29273 19261 29285 19295
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 17368 19196 18276 19224
rect 18509 19227 18567 19233
rect 17368 19184 17374 19196
rect 18509 19193 18521 19227
rect 18555 19193 18567 19227
rect 18509 19187 18567 19193
rect 26050 19184 26056 19236
rect 26108 19184 26114 19236
rect 28442 19184 28448 19236
rect 28500 19184 28506 19236
rect 28721 19227 28779 19233
rect 28721 19193 28733 19227
rect 28767 19224 28779 19227
rect 29288 19224 29316 19255
rect 29546 19233 29552 19236
rect 28767 19196 29316 19224
rect 28767 19193 28779 19196
rect 28721 19187 28779 19193
rect 29540 19187 29552 19233
rect 29546 19184 29552 19187
rect 29604 19184 29610 19236
rect 17126 19156 17132 19168
rect 15712 19128 17132 19156
rect 15712 19116 15718 19128
rect 17126 19116 17132 19128
rect 17184 19116 17190 19168
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 24305 19159 24363 19165
rect 24305 19156 24317 19159
rect 19024 19128 24317 19156
rect 19024 19116 19030 19128
rect 24305 19125 24317 19128
rect 24351 19156 24363 19159
rect 24946 19156 24952 19168
rect 24351 19128 24952 19156
rect 24351 19125 24363 19128
rect 24305 19119 24363 19125
rect 24946 19116 24952 19128
rect 25004 19116 25010 19168
rect 25314 19116 25320 19168
rect 25372 19156 25378 19168
rect 25685 19159 25743 19165
rect 25685 19156 25697 19159
rect 25372 19128 25697 19156
rect 25372 19116 25378 19128
rect 25685 19125 25697 19128
rect 25731 19125 25743 19159
rect 25685 19119 25743 19125
rect 25853 19159 25911 19165
rect 25853 19125 25865 19159
rect 25899 19156 25911 19159
rect 26234 19156 26240 19168
rect 25899 19128 26240 19156
rect 25899 19125 25911 19128
rect 25853 19119 25911 19125
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 26418 19116 26424 19168
rect 26476 19156 26482 19168
rect 26605 19159 26663 19165
rect 26605 19156 26617 19159
rect 26476 19128 26617 19156
rect 26476 19116 26482 19128
rect 26605 19125 26617 19128
rect 26651 19125 26663 19159
rect 26605 19119 26663 19125
rect 26878 19116 26884 19168
rect 26936 19156 26942 19168
rect 28994 19156 29000 19168
rect 26936 19128 29000 19156
rect 26936 19116 26942 19128
rect 28994 19116 29000 19128
rect 29052 19116 29058 19168
rect 29089 19159 29147 19165
rect 29089 19125 29101 19159
rect 29135 19156 29147 19159
rect 29362 19156 29368 19168
rect 29135 19128 29368 19156
rect 29135 19125 29147 19128
rect 29089 19119 29147 19125
rect 29362 19116 29368 19128
rect 29420 19116 29426 19168
rect 29454 19116 29460 19168
rect 29512 19156 29518 19168
rect 30653 19159 30711 19165
rect 30653 19156 30665 19159
rect 29512 19128 30665 19156
rect 29512 19116 29518 19128
rect 30653 19125 30665 19128
rect 30699 19125 30711 19159
rect 30653 19119 30711 19125
rect 552 19066 31648 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 12096 19066
rect 12148 19014 12160 19066
rect 12212 19014 12224 19066
rect 12276 19014 12288 19066
rect 12340 19014 12352 19066
rect 12404 19014 19870 19066
rect 19922 19014 19934 19066
rect 19986 19014 19998 19066
rect 20050 19014 20062 19066
rect 20114 19014 20126 19066
rect 20178 19014 27644 19066
rect 27696 19014 27708 19066
rect 27760 19014 27772 19066
rect 27824 19014 27836 19066
rect 27888 19014 27900 19066
rect 27952 19014 31648 19066
rect 552 18992 31648 19014
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 3234 18952 3240 18964
rect 3007 18924 3240 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 5718 18912 5724 18964
rect 5776 18952 5782 18964
rect 5813 18955 5871 18961
rect 5813 18952 5825 18955
rect 5776 18924 5825 18952
rect 5776 18912 5782 18924
rect 5813 18921 5825 18924
rect 5859 18952 5871 18955
rect 8386 18952 8392 18964
rect 5859 18924 8392 18952
rect 5859 18921 5871 18924
rect 5813 18915 5871 18921
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 8665 18955 8723 18961
rect 8665 18921 8677 18955
rect 8711 18952 8723 18955
rect 9122 18952 9128 18964
rect 8711 18924 9128 18952
rect 8711 18921 8723 18924
rect 8665 18915 8723 18921
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 9306 18912 9312 18964
rect 9364 18952 9370 18964
rect 10502 18952 10508 18964
rect 9364 18924 10508 18952
rect 9364 18912 9370 18924
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 10652 18924 12572 18952
rect 10652 18912 10658 18924
rect 1848 18887 1906 18893
rect 1848 18853 1860 18887
rect 1894 18884 1906 18887
rect 3053 18887 3111 18893
rect 3053 18884 3065 18887
rect 1894 18856 3065 18884
rect 1894 18853 1906 18856
rect 1848 18847 1906 18853
rect 3053 18853 3065 18856
rect 3099 18853 3111 18887
rect 3053 18847 3111 18853
rect 3142 18844 3148 18896
rect 3200 18884 3206 18896
rect 8938 18884 8944 18896
rect 3200 18856 8944 18884
rect 3200 18844 3206 18856
rect 1578 18776 1584 18828
rect 1636 18776 1642 18828
rect 3326 18776 3332 18828
rect 3384 18776 3390 18828
rect 3418 18776 3424 18828
rect 3476 18776 3482 18828
rect 3712 18825 3740 18856
rect 8938 18844 8944 18856
rect 8996 18844 9002 18896
rect 9401 18887 9459 18893
rect 9401 18884 9413 18887
rect 9140 18856 9413 18884
rect 3513 18819 3571 18825
rect 3513 18785 3525 18819
rect 3559 18785 3571 18819
rect 3513 18779 3571 18785
rect 3697 18819 3755 18825
rect 3697 18785 3709 18819
rect 3743 18785 3755 18819
rect 3697 18779 3755 18785
rect 3528 18748 3556 18779
rect 4062 18776 4068 18828
rect 4120 18816 4126 18828
rect 5353 18819 5411 18825
rect 5353 18816 5365 18819
rect 4120 18788 5365 18816
rect 4120 18776 4126 18788
rect 5353 18785 5365 18788
rect 5399 18785 5411 18819
rect 5353 18779 5411 18785
rect 5537 18819 5595 18825
rect 5537 18785 5549 18819
rect 5583 18816 5595 18819
rect 5902 18816 5908 18828
rect 5583 18788 5908 18816
rect 5583 18785 5595 18788
rect 5537 18779 5595 18785
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18816 6147 18819
rect 6454 18816 6460 18828
rect 6135 18788 6460 18816
rect 6135 18785 6147 18788
rect 6089 18779 6147 18785
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 8849 18819 8907 18825
rect 8849 18816 8861 18819
rect 7800 18788 8861 18816
rect 7800 18776 7806 18788
rect 8849 18785 8861 18788
rect 8895 18816 8907 18819
rect 9030 18816 9036 18828
rect 8895 18788 9036 18816
rect 8895 18785 8907 18788
rect 8849 18779 8907 18785
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 9140 18825 9168 18856
rect 9401 18853 9413 18856
rect 9447 18853 9459 18887
rect 10226 18884 10232 18896
rect 9401 18847 9459 18853
rect 9508 18856 10232 18884
rect 9125 18819 9183 18825
rect 9125 18785 9137 18819
rect 9171 18785 9183 18819
rect 9125 18779 9183 18785
rect 9306 18776 9312 18828
rect 9364 18776 9370 18828
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 3528 18720 4537 18748
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18717 4859 18751
rect 4801 18711 4859 18717
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18717 4951 18751
rect 4893 18711 4951 18717
rect 4246 18640 4252 18692
rect 4304 18680 4310 18692
rect 4816 18680 4844 18711
rect 4304 18652 4844 18680
rect 4908 18680 4936 18711
rect 4982 18708 4988 18760
rect 5040 18708 5046 18760
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 6972 18720 8953 18748
rect 6972 18708 6978 18720
rect 8941 18717 8953 18720
rect 8987 18748 8999 18751
rect 9508 18748 9536 18856
rect 10226 18844 10232 18856
rect 10284 18844 10290 18896
rect 10318 18844 10324 18896
rect 10376 18884 10382 18896
rect 10965 18887 11023 18893
rect 10965 18884 10977 18887
rect 10376 18856 10977 18884
rect 10376 18844 10382 18856
rect 10965 18853 10977 18856
rect 11011 18853 11023 18887
rect 10965 18847 11023 18853
rect 11054 18844 11060 18896
rect 11112 18884 11118 18896
rect 11333 18887 11391 18893
rect 11333 18884 11345 18887
rect 11112 18856 11345 18884
rect 11112 18844 11118 18856
rect 11333 18853 11345 18856
rect 11379 18884 11391 18887
rect 11425 18887 11483 18893
rect 11425 18884 11437 18887
rect 11379 18856 11437 18884
rect 11379 18853 11391 18856
rect 11333 18847 11391 18853
rect 11425 18853 11437 18856
rect 11471 18853 11483 18887
rect 11425 18847 11483 18853
rect 12544 18884 12572 18924
rect 14734 18912 14740 18964
rect 14792 18952 14798 18964
rect 14921 18955 14979 18961
rect 14921 18952 14933 18955
rect 14792 18924 14933 18952
rect 14792 18912 14798 18924
rect 14921 18921 14933 18924
rect 14967 18921 14979 18955
rect 14921 18915 14979 18921
rect 15194 18912 15200 18964
rect 15252 18952 15258 18964
rect 15746 18952 15752 18964
rect 15252 18924 15752 18952
rect 15252 18912 15258 18924
rect 15746 18912 15752 18924
rect 15804 18952 15810 18964
rect 16482 18952 16488 18964
rect 15804 18924 16488 18952
rect 15804 18912 15810 18924
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 16666 18912 16672 18964
rect 16724 18952 16730 18964
rect 16761 18955 16819 18961
rect 16761 18952 16773 18955
rect 16724 18924 16773 18952
rect 16724 18912 16730 18924
rect 16761 18921 16773 18924
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 18693 18955 18751 18961
rect 18693 18952 18705 18955
rect 18196 18924 18705 18952
rect 18196 18912 18202 18924
rect 18693 18921 18705 18924
rect 18739 18921 18751 18955
rect 24854 18952 24860 18964
rect 18693 18915 18751 18921
rect 21192 18924 24860 18952
rect 12618 18884 12624 18896
rect 12544 18856 12624 18884
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10137 18819 10195 18825
rect 10060 18816 10149 18819
rect 9824 18791 10149 18816
rect 9824 18788 10088 18791
rect 9824 18776 9830 18788
rect 10137 18785 10149 18791
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 10502 18776 10508 18828
rect 10560 18776 10566 18828
rect 11146 18776 11152 18828
rect 11204 18776 11210 18828
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 11790 18816 11796 18828
rect 11655 18788 11796 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 11974 18776 11980 18828
rect 12032 18816 12038 18828
rect 12115 18819 12173 18825
rect 12115 18816 12127 18819
rect 12032 18788 12127 18816
rect 12032 18776 12038 18788
rect 12115 18785 12127 18788
rect 12161 18785 12173 18819
rect 12115 18779 12173 18785
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18785 12311 18819
rect 12253 18779 12311 18785
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18816 12403 18819
rect 12434 18816 12440 18828
rect 12391 18788 12440 18816
rect 12391 18785 12403 18788
rect 12345 18779 12403 18785
rect 8987 18720 9536 18748
rect 8987 18717 8999 18720
rect 8941 18711 8999 18717
rect 9582 18708 9588 18760
rect 9640 18708 9646 18760
rect 9674 18708 9680 18760
rect 9732 18708 9738 18760
rect 10042 18708 10048 18760
rect 10100 18708 10106 18760
rect 10686 18708 10692 18760
rect 10744 18748 10750 18760
rect 12268 18748 12296 18779
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 12544 18825 12572 18856
rect 12618 18844 12624 18856
rect 12676 18884 12682 18896
rect 13814 18884 13820 18896
rect 12676 18856 13820 18884
rect 12676 18844 12682 18856
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 17034 18884 17040 18896
rect 16316 18856 17040 18884
rect 12529 18819 12587 18825
rect 12529 18785 12541 18819
rect 12575 18785 12587 18819
rect 12529 18779 12587 18785
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 13722 18816 13728 18828
rect 12860 18788 13728 18816
rect 12860 18776 12866 18788
rect 13722 18776 13728 18788
rect 13780 18816 13786 18828
rect 14829 18819 14887 18825
rect 14829 18816 14841 18819
rect 13780 18788 14841 18816
rect 13780 18776 13786 18788
rect 14829 18785 14841 18788
rect 14875 18816 14887 18819
rect 14918 18816 14924 18828
rect 14875 18788 14924 18816
rect 14875 18785 14887 18788
rect 14829 18779 14887 18785
rect 14918 18776 14924 18788
rect 14976 18776 14982 18828
rect 15562 18776 15568 18828
rect 15620 18776 15626 18828
rect 15930 18776 15936 18828
rect 15988 18816 15994 18828
rect 16316 18825 16344 18856
rect 17034 18844 17040 18856
rect 17092 18844 17098 18896
rect 21082 18884 21088 18896
rect 19076 18856 21088 18884
rect 19076 18828 19104 18856
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 16117 18819 16175 18825
rect 16117 18816 16129 18819
rect 15988 18788 16129 18816
rect 15988 18776 15994 18788
rect 16117 18785 16129 18788
rect 16163 18785 16175 18819
rect 16117 18779 16175 18785
rect 16301 18819 16359 18825
rect 16301 18785 16313 18819
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 16393 18819 16451 18825
rect 16393 18785 16405 18819
rect 16439 18785 16451 18819
rect 16393 18779 16451 18785
rect 12986 18748 12992 18760
rect 10744 18720 12992 18748
rect 10744 18708 10750 18720
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 15654 18748 15660 18760
rect 14608 18720 15660 18748
rect 14608 18708 14614 18720
rect 15654 18708 15660 18720
rect 15712 18748 15718 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15712 18720 15853 18748
rect 15712 18708 15718 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 16408 18748 16436 18779
rect 16482 18776 16488 18828
rect 16540 18816 16546 18828
rect 17218 18816 17224 18828
rect 16540 18788 17224 18816
rect 16540 18776 16546 18788
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 18690 18776 18696 18828
rect 18748 18776 18754 18828
rect 18782 18776 18788 18828
rect 18840 18816 18846 18828
rect 18877 18819 18935 18825
rect 18877 18816 18889 18819
rect 18840 18788 18889 18816
rect 18840 18776 18846 18788
rect 18877 18785 18889 18788
rect 18923 18816 18935 18819
rect 19058 18816 19064 18828
rect 18923 18788 19064 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 19058 18776 19064 18788
rect 19116 18776 19122 18828
rect 19521 18819 19579 18825
rect 19521 18785 19533 18819
rect 19567 18816 19579 18819
rect 20622 18816 20628 18828
rect 19567 18788 20628 18816
rect 19567 18785 19579 18788
rect 19521 18779 19579 18785
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 16758 18748 16764 18760
rect 16408 18720 16764 18748
rect 15841 18711 15899 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 21192 18748 21220 18924
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 27982 18952 27988 18964
rect 25740 18924 27988 18952
rect 25740 18912 25746 18924
rect 27982 18912 27988 18924
rect 28040 18912 28046 18964
rect 28074 18912 28080 18964
rect 28132 18952 28138 18964
rect 29273 18955 29331 18961
rect 28132 18924 28856 18952
rect 28132 18912 28138 18924
rect 22370 18844 22376 18896
rect 22428 18893 22434 18896
rect 22428 18884 22440 18893
rect 28718 18884 28724 18896
rect 22428 18856 22473 18884
rect 25700 18856 28724 18884
rect 22428 18847 22440 18856
rect 22428 18844 22434 18847
rect 22002 18776 22008 18828
rect 22060 18816 22066 18828
rect 25700 18825 25728 18856
rect 28718 18844 28724 18856
rect 28776 18844 28782 18896
rect 28828 18884 28856 18924
rect 29273 18921 29285 18955
rect 29319 18952 29331 18955
rect 29546 18952 29552 18964
rect 29319 18924 29552 18952
rect 29319 18921 29331 18924
rect 29273 18915 29331 18921
rect 29546 18912 29552 18924
rect 29604 18912 29610 18964
rect 29454 18884 29460 18896
rect 28828 18856 28948 18884
rect 25685 18819 25743 18825
rect 22060 18788 24164 18816
rect 22060 18776 22066 18788
rect 19260 18720 21220 18748
rect 22649 18751 22707 18757
rect 8846 18680 8852 18692
rect 4908 18652 8852 18680
rect 4304 18640 4310 18652
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 9033 18683 9091 18689
rect 9033 18649 9045 18683
rect 9079 18680 9091 18683
rect 9490 18680 9496 18692
rect 9079 18652 9496 18680
rect 9079 18649 9091 18652
rect 9033 18643 9091 18649
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 11793 18683 11851 18689
rect 9646 18652 10732 18680
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4798 18612 4804 18624
rect 4212 18584 4804 18612
rect 4212 18572 4218 18584
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 5166 18572 5172 18624
rect 5224 18572 5230 18624
rect 5994 18572 6000 18624
rect 6052 18572 6058 18624
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 9646 18612 9674 18652
rect 8628 18584 9674 18612
rect 8628 18572 8634 18584
rect 10226 18572 10232 18624
rect 10284 18572 10290 18624
rect 10704 18621 10732 18652
rect 11793 18649 11805 18683
rect 11839 18680 11851 18683
rect 13078 18680 13084 18692
rect 11839 18652 13084 18680
rect 11839 18649 11851 18652
rect 11793 18643 11851 18649
rect 13078 18640 13084 18652
rect 13136 18640 13142 18692
rect 15749 18683 15807 18689
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 16942 18680 16948 18692
rect 15795 18652 16948 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 10689 18615 10747 18621
rect 10689 18581 10701 18615
rect 10735 18581 10747 18615
rect 10689 18575 10747 18581
rect 11885 18615 11943 18621
rect 11885 18581 11897 18615
rect 11931 18612 11943 18615
rect 11974 18612 11980 18624
rect 11931 18584 11980 18612
rect 11931 18581 11943 18584
rect 11885 18575 11943 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 15657 18615 15715 18621
rect 15657 18581 15669 18615
rect 15703 18612 15715 18615
rect 15838 18612 15844 18624
rect 15703 18584 15844 18612
rect 15703 18581 15715 18584
rect 15657 18575 15715 18581
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16114 18572 16120 18624
rect 16172 18612 16178 18624
rect 17034 18612 17040 18624
rect 16172 18584 17040 18612
rect 16172 18572 16178 18584
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 19058 18572 19064 18624
rect 19116 18612 19122 18624
rect 19260 18621 19288 18720
rect 22649 18717 22661 18751
rect 22695 18748 22707 18751
rect 23474 18748 23480 18760
rect 22695 18720 23480 18748
rect 22695 18717 22707 18720
rect 22649 18711 22707 18717
rect 19245 18615 19303 18621
rect 19245 18612 19257 18615
rect 19116 18584 19257 18612
rect 19116 18572 19122 18584
rect 19245 18581 19257 18584
rect 19291 18581 19303 18615
rect 19245 18575 19303 18581
rect 21266 18572 21272 18624
rect 21324 18572 21330 18624
rect 21358 18572 21364 18624
rect 21416 18612 21422 18624
rect 22664 18612 22692 18711
rect 23474 18708 23480 18720
rect 23532 18708 23538 18760
rect 24026 18708 24032 18760
rect 24084 18708 24090 18760
rect 24136 18748 24164 18788
rect 25685 18785 25697 18819
rect 25731 18785 25743 18819
rect 25685 18779 25743 18785
rect 26418 18776 26424 18828
rect 26476 18776 26482 18828
rect 26510 18776 26516 18828
rect 26568 18816 26574 18828
rect 26677 18819 26735 18825
rect 26677 18816 26689 18819
rect 26568 18788 26689 18816
rect 26568 18776 26574 18788
rect 26677 18785 26689 18788
rect 26723 18785 26735 18819
rect 26677 18779 26735 18785
rect 28629 18819 28687 18825
rect 28629 18785 28641 18819
rect 28675 18785 28687 18819
rect 28629 18779 28687 18785
rect 24854 18757 24860 18760
rect 24673 18751 24731 18757
rect 24673 18748 24685 18751
rect 24136 18720 24685 18748
rect 24673 18717 24685 18720
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 24832 18751 24860 18757
rect 24832 18717 24844 18751
rect 24832 18711 24860 18717
rect 24854 18708 24860 18711
rect 24912 18708 24918 18760
rect 24946 18708 24952 18760
rect 25004 18708 25010 18760
rect 25866 18708 25872 18760
rect 25924 18708 25930 18760
rect 28644 18748 28672 18779
rect 28810 18776 28816 18828
rect 28868 18776 28874 18828
rect 28920 18825 28948 18856
rect 29012 18856 29460 18884
rect 29012 18828 29040 18856
rect 29454 18844 29460 18856
rect 29512 18844 29518 18896
rect 29564 18856 31064 18884
rect 28905 18819 28963 18825
rect 28905 18785 28917 18819
rect 28951 18785 28963 18819
rect 28905 18779 28963 18785
rect 28994 18776 29000 18828
rect 29052 18776 29058 18828
rect 29362 18776 29368 18828
rect 29420 18776 29426 18828
rect 29564 18816 29592 18856
rect 29638 18825 29644 18828
rect 29472 18788 29592 18816
rect 29178 18748 29184 18760
rect 28644 18720 29184 18748
rect 29178 18708 29184 18720
rect 29236 18748 29242 18760
rect 29472 18748 29500 18788
rect 29632 18779 29644 18825
rect 29638 18776 29644 18779
rect 29696 18776 29702 18828
rect 30190 18776 30196 18828
rect 30248 18816 30254 18828
rect 30837 18819 30895 18825
rect 30837 18816 30849 18819
rect 30248 18788 30849 18816
rect 30248 18776 30254 18788
rect 30837 18785 30849 18788
rect 30883 18785 30895 18819
rect 30837 18779 30895 18785
rect 29236 18720 29500 18748
rect 29236 18708 29242 18720
rect 25222 18640 25228 18692
rect 25280 18640 25286 18692
rect 31036 18624 31064 18856
rect 21416 18584 22692 18612
rect 21416 18572 21422 18584
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 27801 18615 27859 18621
rect 27801 18612 27813 18615
rect 27764 18584 27813 18612
rect 27764 18572 27770 18584
rect 27801 18581 27813 18584
rect 27847 18612 27859 18615
rect 28350 18612 28356 18624
rect 27847 18584 28356 18612
rect 27847 18581 27859 18584
rect 27801 18575 27859 18581
rect 28350 18572 28356 18584
rect 28408 18572 28414 18624
rect 28718 18572 28724 18624
rect 28776 18612 28782 18624
rect 30745 18615 30803 18621
rect 30745 18612 30757 18615
rect 28776 18584 30757 18612
rect 28776 18572 28782 18584
rect 30745 18581 30757 18584
rect 30791 18581 30803 18615
rect 30745 18575 30803 18581
rect 31018 18572 31024 18624
rect 31076 18572 31082 18624
rect 552 18522 31648 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 11436 18522
rect 11488 18470 11500 18522
rect 11552 18470 11564 18522
rect 11616 18470 11628 18522
rect 11680 18470 11692 18522
rect 11744 18470 19210 18522
rect 19262 18470 19274 18522
rect 19326 18470 19338 18522
rect 19390 18470 19402 18522
rect 19454 18470 19466 18522
rect 19518 18470 26984 18522
rect 27036 18470 27048 18522
rect 27100 18470 27112 18522
rect 27164 18470 27176 18522
rect 27228 18470 27240 18522
rect 27292 18470 31648 18522
rect 552 18448 31648 18470
rect 4801 18411 4859 18417
rect 4801 18377 4813 18411
rect 4847 18408 4859 18411
rect 4982 18408 4988 18420
rect 4847 18380 4988 18408
rect 4847 18377 4859 18380
rect 4801 18371 4859 18377
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 5166 18368 5172 18420
rect 5224 18368 5230 18420
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6328 18380 6561 18408
rect 6328 18368 6334 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 6549 18371 6607 18377
rect 8018 18368 8024 18420
rect 8076 18408 8082 18420
rect 9858 18408 9864 18420
rect 8076 18380 9864 18408
rect 8076 18368 8082 18380
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 10042 18408 10048 18420
rect 9968 18380 10048 18408
rect 6288 18340 6316 18368
rect 3988 18312 5120 18340
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3234 18204 3240 18216
rect 2915 18176 3240 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 3234 18164 3240 18176
rect 3292 18164 3298 18216
rect 3510 18164 3516 18216
rect 3568 18164 3574 18216
rect 3878 18164 3884 18216
rect 3936 18204 3942 18216
rect 3988 18213 4016 18312
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4249 18275 4307 18281
rect 4249 18272 4261 18275
rect 4120 18244 4261 18272
rect 4120 18232 4126 18244
rect 4249 18241 4261 18244
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 3973 18207 4031 18213
rect 3973 18204 3985 18207
rect 3936 18176 3985 18204
rect 3936 18164 3942 18176
rect 3973 18173 3985 18176
rect 4019 18173 4031 18207
rect 4525 18207 4583 18213
rect 4525 18204 4537 18207
rect 3973 18167 4031 18173
rect 4265 18176 4537 18204
rect 4265 18148 4293 18176
rect 4525 18173 4537 18176
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 4709 18207 4767 18213
rect 4709 18173 4721 18207
rect 4755 18204 4767 18207
rect 4798 18204 4804 18216
rect 4755 18176 4804 18204
rect 4755 18173 4767 18176
rect 4709 18167 4767 18173
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 4982 18164 4988 18216
rect 5040 18164 5046 18216
rect 5092 18204 5120 18312
rect 5184 18312 6316 18340
rect 5184 18281 5212 18312
rect 9030 18300 9036 18352
rect 9088 18340 9094 18352
rect 9306 18340 9312 18352
rect 9088 18312 9312 18340
rect 9088 18300 9094 18312
rect 9306 18300 9312 18312
rect 9364 18340 9370 18352
rect 9968 18340 9996 18380
rect 10042 18368 10048 18380
rect 10100 18408 10106 18420
rect 10100 18380 20576 18408
rect 10100 18368 10106 18380
rect 10502 18340 10508 18352
rect 9364 18312 9996 18340
rect 10060 18312 10508 18340
rect 9364 18300 9370 18312
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18241 5227 18275
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5169 18235 5227 18241
rect 5460 18244 5641 18272
rect 5350 18204 5356 18216
rect 5092 18176 5356 18204
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 2774 18096 2780 18148
rect 2832 18136 2838 18148
rect 3329 18139 3387 18145
rect 3329 18136 3341 18139
rect 2832 18108 3341 18136
rect 2832 18096 2838 18108
rect 3329 18105 3341 18108
rect 3375 18136 3387 18139
rect 3418 18136 3424 18148
rect 3375 18108 3424 18136
rect 3375 18105 3387 18108
rect 3329 18099 3387 18105
rect 3418 18096 3424 18108
rect 3476 18096 3482 18148
rect 4246 18096 4252 18148
rect 4304 18096 4310 18148
rect 5460 18145 5488 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 5810 18272 5816 18284
rect 5767 18244 5816 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 6089 18275 6147 18281
rect 6089 18272 6101 18275
rect 5951 18244 6101 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 6089 18241 6101 18244
rect 6135 18272 6147 18275
rect 6135 18244 6592 18272
rect 6135 18241 6147 18244
rect 6089 18235 6147 18241
rect 5994 18164 6000 18216
rect 6052 18164 6058 18216
rect 6178 18164 6184 18216
rect 6236 18204 6242 18216
rect 6303 18207 6361 18213
rect 6303 18204 6315 18207
rect 6236 18176 6315 18204
rect 6236 18164 6242 18176
rect 6303 18173 6315 18176
rect 6349 18173 6361 18207
rect 6303 18167 6361 18173
rect 6454 18164 6460 18216
rect 6512 18164 6518 18216
rect 6564 18213 6592 18244
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 9214 18272 9220 18284
rect 8996 18244 9220 18272
rect 8996 18232 9002 18244
rect 9214 18232 9220 18244
rect 9272 18272 9278 18284
rect 9272 18244 9904 18272
rect 9272 18232 9278 18244
rect 6549 18207 6607 18213
rect 6549 18173 6561 18207
rect 6595 18173 6607 18207
rect 6549 18167 6607 18173
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18173 6791 18207
rect 6733 18167 6791 18173
rect 5445 18139 5503 18145
rect 5445 18136 5457 18139
rect 4356 18108 5457 18136
rect 2961 18071 3019 18077
rect 2961 18037 2973 18071
rect 3007 18068 3019 18071
rect 3234 18068 3240 18080
rect 3007 18040 3240 18068
rect 3007 18037 3019 18040
rect 2961 18031 3019 18037
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 3436 18068 3464 18096
rect 4356 18068 4384 18108
rect 5445 18105 5457 18108
rect 5491 18105 5503 18139
rect 5445 18099 5503 18105
rect 5626 18096 5632 18148
rect 5684 18136 5690 18148
rect 6748 18136 6776 18167
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8352 18176 8493 18204
rect 8352 18164 8358 18176
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 9401 18207 9459 18213
rect 9401 18173 9413 18207
rect 9447 18204 9459 18207
rect 9876 18204 9904 18244
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 10060 18281 10088 18312
rect 10502 18300 10508 18312
rect 10560 18300 10566 18352
rect 15470 18340 15476 18352
rect 11440 18312 15476 18340
rect 10045 18275 10103 18281
rect 10045 18272 10057 18275
rect 10008 18244 10057 18272
rect 10008 18232 10014 18244
rect 10045 18241 10057 18244
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 10192 18244 10640 18272
rect 10192 18232 10198 18244
rect 10612 18216 10640 18244
rect 9447 18176 9812 18204
rect 9876 18176 9996 18204
rect 9447 18173 9459 18176
rect 9401 18167 9459 18173
rect 5684 18108 6776 18136
rect 5684 18096 5690 18108
rect 3436 18040 4384 18068
rect 4709 18071 4767 18077
rect 4709 18037 4721 18071
rect 4755 18068 4767 18071
rect 4798 18068 4804 18080
rect 4755 18040 4804 18068
rect 4755 18037 4767 18040
rect 4709 18031 4767 18037
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 5166 18028 5172 18080
rect 5224 18068 5230 18080
rect 5537 18071 5595 18077
rect 5537 18068 5549 18071
rect 5224 18040 5549 18068
rect 5224 18028 5230 18040
rect 5537 18037 5549 18040
rect 5583 18037 5595 18071
rect 5537 18031 5595 18037
rect 6178 18028 6184 18080
rect 6236 18068 6242 18080
rect 6454 18068 6460 18080
rect 6236 18040 6460 18068
rect 6236 18028 6242 18040
rect 6454 18028 6460 18040
rect 6512 18068 6518 18080
rect 6822 18068 6828 18080
rect 6512 18040 6828 18068
rect 6512 18028 6518 18040
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 8573 18071 8631 18077
rect 8573 18037 8585 18071
rect 8619 18068 8631 18071
rect 8662 18068 8668 18080
rect 8619 18040 8668 18068
rect 8619 18037 8631 18040
rect 8573 18031 8631 18037
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 8754 18028 8760 18080
rect 8812 18028 8818 18080
rect 9490 18028 9496 18080
rect 9548 18028 9554 18080
rect 9784 18068 9812 18176
rect 9858 18096 9864 18148
rect 9916 18096 9922 18148
rect 9968 18136 9996 18176
rect 10594 18164 10600 18216
rect 10652 18164 10658 18216
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 10778 18164 10784 18216
rect 10836 18164 10842 18216
rect 10870 18164 10876 18216
rect 10928 18204 10934 18216
rect 11440 18213 11468 18312
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 15562 18300 15568 18352
rect 15620 18340 15626 18352
rect 18966 18340 18972 18352
rect 15620 18312 18972 18340
rect 15620 18300 15626 18312
rect 18966 18300 18972 18312
rect 19024 18300 19030 18352
rect 20548 18340 20576 18380
rect 20622 18368 20628 18420
rect 20680 18368 20686 18420
rect 24578 18368 24584 18420
rect 24636 18408 24642 18420
rect 25774 18408 25780 18420
rect 24636 18380 25780 18408
rect 24636 18368 24642 18380
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 26510 18408 26516 18420
rect 26283 18380 26516 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 28810 18368 28816 18420
rect 28868 18368 28874 18420
rect 28920 18380 29132 18408
rect 20898 18340 20904 18352
rect 20548 18312 20904 18340
rect 20898 18300 20904 18312
rect 20956 18340 20962 18352
rect 22002 18340 22008 18352
rect 20956 18312 22008 18340
rect 20956 18300 20962 18312
rect 22002 18300 22008 18312
rect 22060 18300 22066 18352
rect 28350 18300 28356 18352
rect 28408 18340 28414 18352
rect 28920 18340 28948 18380
rect 28408 18312 28948 18340
rect 28997 18343 29055 18349
rect 28408 18300 28414 18312
rect 28997 18309 29009 18343
rect 29043 18309 29055 18343
rect 28997 18303 29055 18309
rect 11790 18232 11796 18284
rect 11848 18232 11854 18284
rect 14182 18272 14188 18284
rect 13280 18244 14188 18272
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10928 18176 10977 18204
rect 10928 18164 10934 18176
rect 10965 18173 10977 18176
rect 11011 18204 11023 18207
rect 11057 18207 11115 18213
rect 11057 18204 11069 18207
rect 11011 18176 11069 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 11057 18173 11069 18176
rect 11103 18173 11115 18207
rect 11057 18167 11115 18173
rect 11425 18207 11483 18213
rect 11425 18173 11437 18207
rect 11471 18173 11483 18207
rect 11425 18167 11483 18173
rect 11440 18136 11468 18167
rect 11606 18164 11612 18216
rect 11664 18204 11670 18216
rect 12345 18207 12403 18213
rect 12345 18204 12357 18207
rect 11664 18176 12357 18204
rect 11664 18164 11670 18176
rect 12345 18173 12357 18176
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 12894 18164 12900 18216
rect 12952 18164 12958 18216
rect 12986 18164 12992 18216
rect 13044 18164 13050 18216
rect 13078 18164 13084 18216
rect 13136 18164 13142 18216
rect 13280 18213 13308 18244
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 13354 18164 13360 18216
rect 13412 18204 13418 18216
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 13412 18176 13553 18204
rect 13412 18164 13418 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 15580 18213 15608 18300
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 15930 18272 15936 18284
rect 15703 18244 15936 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16117 18275 16175 18281
rect 16117 18272 16129 18275
rect 16040 18244 16129 18272
rect 15565 18207 15623 18213
rect 13964 18176 15240 18204
rect 13964 18164 13970 18176
rect 9968 18108 11468 18136
rect 15010 18096 15016 18148
rect 15068 18096 15074 18148
rect 15212 18145 15240 18176
rect 15565 18173 15577 18207
rect 15611 18173 15623 18207
rect 15565 18167 15623 18173
rect 15746 18164 15752 18216
rect 15804 18164 15810 18216
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16040 18213 16068 18244
rect 16117 18241 16129 18244
rect 16163 18241 16175 18275
rect 16393 18275 16451 18281
rect 16393 18272 16405 18275
rect 16117 18235 16175 18241
rect 16224 18244 16405 18272
rect 16224 18216 16252 18244
rect 16393 18241 16405 18244
rect 16439 18241 16451 18275
rect 16393 18235 16451 18241
rect 16577 18275 16635 18281
rect 16577 18241 16589 18275
rect 16623 18272 16635 18275
rect 17034 18272 17040 18284
rect 16623 18244 17040 18272
rect 16623 18241 16635 18244
rect 16577 18235 16635 18241
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 28074 18272 28080 18284
rect 22572 18244 23971 18272
rect 16025 18207 16083 18213
rect 15896 18176 15976 18204
rect 15896 18164 15902 18176
rect 15197 18139 15255 18145
rect 15197 18105 15209 18139
rect 15243 18136 15255 18139
rect 15948 18136 15976 18176
rect 16025 18173 16037 18207
rect 16071 18173 16083 18207
rect 16025 18167 16083 18173
rect 16206 18164 16212 18216
rect 16264 18164 16270 18216
rect 16298 18164 16304 18216
rect 16356 18164 16362 18216
rect 16482 18164 16488 18216
rect 16540 18204 16546 18216
rect 16850 18204 16856 18216
rect 16540 18176 16856 18204
rect 16540 18164 16546 18176
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 18785 18207 18843 18213
rect 18785 18173 18797 18207
rect 18831 18204 18843 18207
rect 18874 18204 18880 18216
rect 18831 18176 18880 18204
rect 18831 18173 18843 18176
rect 18785 18167 18843 18173
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 18966 18164 18972 18216
rect 19024 18164 19030 18216
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19334 18204 19340 18216
rect 19291 18176 19340 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18204 21327 18207
rect 21358 18204 21364 18216
rect 21315 18176 21364 18204
rect 21315 18173 21327 18176
rect 21269 18167 21327 18173
rect 17129 18139 17187 18145
rect 15243 18108 15884 18136
rect 15948 18108 17080 18136
rect 15243 18105 15255 18108
rect 15197 18099 15255 18105
rect 15856 18080 15884 18108
rect 9950 18068 9956 18080
rect 9784 18040 9956 18068
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10321 18071 10379 18077
rect 10321 18068 10333 18071
rect 10192 18040 10333 18068
rect 10192 18028 10198 18040
rect 10321 18037 10333 18040
rect 10367 18037 10379 18071
rect 10321 18031 10379 18037
rect 12618 18028 12624 18080
rect 12676 18028 12682 18080
rect 13630 18028 13636 18080
rect 13688 18068 13694 18080
rect 14185 18071 14243 18077
rect 14185 18068 14197 18071
rect 13688 18040 14197 18068
rect 13688 18028 13694 18040
rect 14185 18037 14197 18040
rect 14231 18037 14243 18071
rect 14185 18031 14243 18037
rect 15381 18071 15439 18077
rect 15381 18037 15393 18071
rect 15427 18068 15439 18071
rect 15654 18068 15660 18080
rect 15427 18040 15660 18068
rect 15427 18037 15439 18040
rect 15381 18031 15439 18037
rect 15654 18028 15660 18040
rect 15712 18028 15718 18080
rect 15838 18028 15844 18080
rect 15896 18028 15902 18080
rect 17052 18077 17080 18108
rect 17129 18105 17141 18139
rect 17175 18136 17187 18139
rect 17310 18136 17316 18148
rect 17175 18108 17316 18136
rect 17175 18105 17187 18108
rect 17129 18099 17187 18105
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 19518 18145 19524 18148
rect 19512 18099 19524 18145
rect 19518 18096 19524 18099
rect 19576 18096 19582 18148
rect 19610 18096 19616 18148
rect 19668 18136 19674 18148
rect 19794 18136 19800 18148
rect 19668 18108 19800 18136
rect 19668 18096 19674 18108
rect 19794 18096 19800 18108
rect 19852 18136 19858 18148
rect 20622 18136 20628 18148
rect 19852 18108 20628 18136
rect 19852 18096 19858 18108
rect 20622 18096 20628 18108
rect 20680 18136 20686 18148
rect 21284 18136 21312 18167
rect 21358 18164 21364 18176
rect 21416 18164 21422 18216
rect 21818 18164 21824 18216
rect 21876 18204 21882 18216
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 21876 18176 22293 18204
rect 21876 18164 21882 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 22462 18164 22468 18216
rect 22520 18164 22526 18216
rect 22572 18213 22600 18244
rect 22557 18207 22615 18213
rect 22557 18173 22569 18207
rect 22603 18173 22615 18207
rect 22557 18167 22615 18173
rect 22649 18207 22707 18213
rect 22649 18173 22661 18207
rect 22695 18173 22707 18207
rect 22649 18167 22707 18173
rect 20680 18108 21312 18136
rect 20680 18096 20686 18108
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 18690 18068 18696 18080
rect 17083 18040 18696 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 18969 18071 19027 18077
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 19058 18068 19064 18080
rect 19015 18040 19064 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 20438 18068 20444 18080
rect 19484 18040 20444 18068
rect 19484 18028 19490 18040
rect 20438 18028 20444 18040
rect 20496 18068 20502 18080
rect 21836 18068 21864 18164
rect 22664 18136 22692 18167
rect 23474 18164 23480 18216
rect 23532 18164 23538 18216
rect 23569 18207 23627 18213
rect 23569 18173 23581 18207
rect 23615 18204 23627 18207
rect 23845 18207 23903 18213
rect 23845 18204 23857 18207
rect 23615 18176 23857 18204
rect 23615 18173 23627 18176
rect 23569 18167 23627 18173
rect 23845 18173 23857 18176
rect 23891 18173 23903 18207
rect 23943 18204 23971 18244
rect 25424 18244 28080 18272
rect 24394 18204 24400 18216
rect 23943 18176 24400 18204
rect 23845 18167 23903 18173
rect 24394 18164 24400 18176
rect 24452 18204 24458 18216
rect 25424 18204 25452 18244
rect 24452 18176 25452 18204
rect 24452 18164 24458 18176
rect 25498 18164 25504 18216
rect 25556 18164 25562 18216
rect 25590 18164 25596 18216
rect 25648 18204 25654 18216
rect 25685 18207 25743 18213
rect 25685 18204 25697 18207
rect 25648 18176 25697 18204
rect 25648 18164 25654 18176
rect 25685 18173 25697 18176
rect 25731 18173 25743 18207
rect 25685 18167 25743 18173
rect 25774 18164 25780 18216
rect 25832 18164 25838 18216
rect 25866 18164 25872 18216
rect 25924 18164 25930 18216
rect 26620 18213 26648 18244
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 28442 18272 28448 18284
rect 28276 18244 28448 18272
rect 26513 18207 26571 18213
rect 26513 18173 26525 18207
rect 26559 18173 26571 18207
rect 26513 18167 26571 18173
rect 26605 18207 26663 18213
rect 26605 18173 26617 18207
rect 26651 18173 26663 18207
rect 26605 18167 26663 18173
rect 24118 18145 24124 18148
rect 22296 18108 22692 18136
rect 22296 18080 22324 18108
rect 24112 18099 24124 18145
rect 24118 18096 24124 18099
rect 24176 18096 24182 18148
rect 24854 18096 24860 18148
rect 24912 18136 24918 18148
rect 26528 18136 26556 18167
rect 26694 18164 26700 18216
rect 26752 18164 26758 18216
rect 26878 18164 26884 18216
rect 26936 18164 26942 18216
rect 27982 18164 27988 18216
rect 28040 18164 28046 18216
rect 28166 18164 28172 18216
rect 28224 18164 28230 18216
rect 28276 18213 28304 18244
rect 28442 18232 28448 18244
rect 28500 18232 28506 18284
rect 28261 18207 28319 18213
rect 28261 18173 28273 18207
rect 28307 18173 28319 18207
rect 28261 18167 28319 18173
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18173 28411 18207
rect 28353 18167 28411 18173
rect 26786 18136 26792 18148
rect 24912 18108 26792 18136
rect 24912 18096 24918 18108
rect 26786 18096 26792 18108
rect 26844 18136 26850 18148
rect 27706 18136 27712 18148
rect 26844 18108 27712 18136
rect 26844 18096 26850 18108
rect 27706 18096 27712 18108
rect 27764 18096 27770 18148
rect 27801 18139 27859 18145
rect 27801 18105 27813 18139
rect 27847 18136 27859 18139
rect 28184 18136 28212 18164
rect 27847 18108 28212 18136
rect 28368 18136 28396 18167
rect 28534 18164 28540 18216
rect 28592 18164 28598 18216
rect 28629 18207 28687 18213
rect 28629 18173 28641 18207
rect 28675 18204 28687 18207
rect 29012 18204 29040 18303
rect 29104 18272 29132 18380
rect 29638 18368 29644 18420
rect 29696 18408 29702 18420
rect 29825 18411 29883 18417
rect 29825 18408 29837 18411
rect 29696 18380 29837 18408
rect 29696 18368 29702 18380
rect 29825 18377 29837 18380
rect 29871 18377 29883 18411
rect 29825 18371 29883 18377
rect 29362 18300 29368 18352
rect 29420 18340 29426 18352
rect 29420 18312 30236 18340
rect 29420 18300 29426 18312
rect 29457 18275 29515 18281
rect 29457 18272 29469 18275
rect 29104 18244 29469 18272
rect 29457 18241 29469 18244
rect 29503 18241 29515 18275
rect 29457 18235 29515 18241
rect 29546 18232 29552 18284
rect 29604 18232 29610 18284
rect 30208 18213 30236 18312
rect 30101 18207 30159 18213
rect 30101 18204 30113 18207
rect 28675 18176 29040 18204
rect 29380 18176 30113 18204
rect 28675 18173 28687 18176
rect 28629 18167 28687 18173
rect 28994 18136 29000 18148
rect 28368 18108 29000 18136
rect 27847 18105 27859 18108
rect 27801 18099 27859 18105
rect 28994 18096 29000 18108
rect 29052 18096 29058 18148
rect 29086 18096 29092 18148
rect 29144 18136 29150 18148
rect 29380 18145 29408 18176
rect 30101 18173 30113 18176
rect 30147 18173 30159 18207
rect 30101 18167 30159 18173
rect 30193 18207 30251 18213
rect 30193 18173 30205 18207
rect 30239 18173 30251 18207
rect 30193 18167 30251 18173
rect 30285 18207 30343 18213
rect 30285 18173 30297 18207
rect 30331 18204 30343 18207
rect 30374 18204 30380 18216
rect 30331 18176 30380 18204
rect 30331 18173 30343 18176
rect 30285 18167 30343 18173
rect 30374 18164 30380 18176
rect 30432 18164 30438 18216
rect 30469 18207 30527 18213
rect 30469 18173 30481 18207
rect 30515 18204 30527 18207
rect 31018 18204 31024 18216
rect 30515 18176 31024 18204
rect 30515 18173 30527 18176
rect 30469 18167 30527 18173
rect 31018 18164 31024 18176
rect 31076 18164 31082 18216
rect 29365 18139 29423 18145
rect 29365 18136 29377 18139
rect 29144 18108 29377 18136
rect 29144 18096 29150 18108
rect 29365 18105 29377 18108
rect 29411 18105 29423 18139
rect 29365 18099 29423 18105
rect 20496 18040 21864 18068
rect 20496 18028 20502 18040
rect 22278 18028 22284 18080
rect 22336 18028 22342 18080
rect 22925 18071 22983 18077
rect 22925 18037 22937 18071
rect 22971 18068 22983 18071
rect 23290 18068 23296 18080
rect 22971 18040 23296 18068
rect 22971 18037 22983 18040
rect 22925 18031 22983 18037
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 24946 18028 24952 18080
rect 25004 18068 25010 18080
rect 25130 18068 25136 18080
rect 25004 18040 25136 18068
rect 25004 18028 25010 18040
rect 25130 18028 25136 18040
rect 25188 18068 25194 18080
rect 25225 18071 25283 18077
rect 25225 18068 25237 18071
rect 25188 18040 25237 18068
rect 25188 18028 25194 18040
rect 25225 18037 25237 18040
rect 25271 18037 25283 18071
rect 25225 18031 25283 18037
rect 26145 18071 26203 18077
rect 26145 18037 26157 18071
rect 26191 18068 26203 18071
rect 28074 18068 28080 18080
rect 26191 18040 28080 18068
rect 26191 18037 26203 18040
rect 26145 18031 26203 18037
rect 28074 18028 28080 18040
rect 28132 18028 28138 18080
rect 28169 18071 28227 18077
rect 28169 18037 28181 18071
rect 28215 18068 28227 18071
rect 29270 18068 29276 18080
rect 28215 18040 29276 18068
rect 28215 18037 28227 18040
rect 28169 18031 28227 18037
rect 29270 18028 29276 18040
rect 29328 18028 29334 18080
rect 552 17978 31648 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 12096 17978
rect 12148 17926 12160 17978
rect 12212 17926 12224 17978
rect 12276 17926 12288 17978
rect 12340 17926 12352 17978
rect 12404 17926 19870 17978
rect 19922 17926 19934 17978
rect 19986 17926 19998 17978
rect 20050 17926 20062 17978
rect 20114 17926 20126 17978
rect 20178 17926 27644 17978
rect 27696 17926 27708 17978
rect 27760 17926 27772 17978
rect 27824 17926 27836 17978
rect 27888 17926 27900 17978
rect 27952 17926 31648 17978
rect 552 17904 31648 17926
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 3878 17864 3884 17876
rect 3476 17836 3884 17864
rect 3476 17824 3482 17836
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 3973 17867 4031 17873
rect 3973 17833 3985 17867
rect 4019 17833 4031 17867
rect 3973 17827 4031 17833
rect 5629 17867 5687 17873
rect 5629 17833 5641 17867
rect 5675 17864 5687 17867
rect 5718 17864 5724 17876
rect 5675 17836 5724 17864
rect 5675 17833 5687 17836
rect 5629 17827 5687 17833
rect 3988 17796 4016 17827
rect 5718 17824 5724 17836
rect 5776 17824 5782 17876
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 6052 17836 6592 17864
rect 6052 17824 6058 17836
rect 2884 17768 4016 17796
rect 2682 17688 2688 17740
rect 2740 17688 2746 17740
rect 2774 17688 2780 17740
rect 2832 17688 2838 17740
rect 2884 17737 2912 17768
rect 4154 17756 4160 17808
rect 4212 17756 4218 17808
rect 4982 17756 4988 17808
rect 5040 17796 5046 17808
rect 5534 17796 5540 17808
rect 5040 17768 5540 17796
rect 5040 17756 5046 17768
rect 2869 17731 2927 17737
rect 2869 17697 2881 17731
rect 2915 17697 2927 17731
rect 2869 17691 2927 17697
rect 3050 17688 3056 17740
rect 3108 17688 3114 17740
rect 3697 17731 3755 17737
rect 3697 17697 3709 17731
rect 3743 17728 3755 17731
rect 3743 17700 3777 17728
rect 3743 17697 3755 17700
rect 3697 17691 3755 17697
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17629 3203 17663
rect 3145 17623 3203 17629
rect 3605 17663 3663 17669
rect 3605 17629 3617 17663
rect 3651 17660 3663 17663
rect 3712 17660 3740 17691
rect 3878 17688 3884 17740
rect 3936 17688 3942 17740
rect 4062 17688 4068 17740
rect 4120 17688 4126 17740
rect 4172 17728 4200 17756
rect 4341 17731 4399 17737
rect 4341 17728 4353 17731
rect 4172 17700 4353 17728
rect 4341 17697 4353 17700
rect 4387 17697 4399 17731
rect 4341 17691 4399 17697
rect 4522 17688 4528 17740
rect 4580 17728 4586 17740
rect 5092 17737 5120 17768
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 6454 17796 6460 17808
rect 6104 17768 6460 17796
rect 6104 17740 6132 17768
rect 6454 17756 6460 17768
rect 6512 17756 6518 17808
rect 6564 17805 6592 17836
rect 6914 17824 6920 17876
rect 6972 17824 6978 17876
rect 8205 17867 8263 17873
rect 8205 17833 8217 17867
rect 8251 17864 8263 17867
rect 8251 17836 9812 17864
rect 8251 17833 8263 17836
rect 8205 17827 8263 17833
rect 6549 17799 6607 17805
rect 6549 17765 6561 17799
rect 6595 17765 6607 17799
rect 6549 17759 6607 17765
rect 6638 17756 6644 17808
rect 6696 17796 6702 17808
rect 8389 17799 8447 17805
rect 6696 17768 7052 17796
rect 6696 17756 6702 17768
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4580 17700 4813 17728
rect 4580 17688 4586 17700
rect 4801 17697 4813 17700
rect 4847 17697 4859 17731
rect 4801 17691 4859 17697
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17697 4951 17731
rect 4893 17691 4951 17697
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17697 5135 17731
rect 5077 17691 5135 17697
rect 4080 17660 4108 17688
rect 3651 17632 4108 17660
rect 3651 17629 3663 17632
rect 3605 17623 3663 17629
rect 2406 17484 2412 17536
rect 2464 17484 2470 17536
rect 3160 17524 3188 17623
rect 4154 17620 4160 17672
rect 4212 17620 4218 17672
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17629 4307 17663
rect 4249 17623 4307 17629
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 4479 17632 4629 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 4908 17660 4936 17691
rect 5166 17688 5172 17740
rect 5224 17688 5230 17740
rect 5258 17688 5264 17740
rect 5316 17688 5322 17740
rect 5442 17688 5448 17740
rect 5500 17688 5506 17740
rect 5997 17731 6055 17737
rect 5997 17728 6009 17731
rect 5552 17700 6009 17728
rect 5350 17660 5356 17672
rect 4908 17632 5356 17660
rect 4617 17623 4675 17629
rect 3234 17552 3240 17604
rect 3292 17592 3298 17604
rect 3421 17595 3479 17601
rect 3421 17592 3433 17595
rect 3292 17564 3433 17592
rect 3292 17552 3298 17564
rect 3421 17561 3433 17564
rect 3467 17561 3479 17595
rect 3421 17555 3479 17561
rect 3881 17595 3939 17601
rect 3881 17561 3893 17595
rect 3927 17592 3939 17595
rect 4062 17592 4068 17604
rect 3927 17564 4068 17592
rect 3927 17561 3939 17564
rect 3881 17555 3939 17561
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 4154 17524 4160 17536
rect 3160 17496 4160 17524
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 4265 17524 4293 17623
rect 5350 17620 5356 17632
rect 5408 17660 5414 17672
rect 5552 17660 5580 17700
rect 5997 17697 6009 17700
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 6086 17688 6092 17740
rect 6144 17688 6150 17740
rect 6178 17688 6184 17740
rect 6236 17688 6242 17740
rect 6362 17737 6368 17740
rect 6319 17731 6368 17737
rect 6319 17697 6331 17731
rect 6365 17697 6368 17731
rect 6319 17691 6368 17697
rect 6362 17688 6368 17691
rect 6420 17728 6426 17740
rect 6420 17700 6684 17728
rect 6420 17688 6426 17700
rect 5408 17632 5580 17660
rect 5408 17620 5414 17632
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 6104 17660 6132 17688
rect 5868 17632 6132 17660
rect 5868 17620 5874 17632
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 6656 17660 6684 17700
rect 6730 17688 6736 17740
rect 6788 17688 6794 17740
rect 7024 17737 7052 17768
rect 8389 17765 8401 17799
rect 8435 17796 8447 17799
rect 8754 17796 8760 17808
rect 8435 17768 8760 17796
rect 8435 17765 8447 17768
rect 8389 17759 8447 17765
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 9674 17796 9680 17808
rect 8864 17768 9680 17796
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17697 7067 17731
rect 7009 17691 7067 17697
rect 7098 17688 7104 17740
rect 7156 17728 7162 17740
rect 7193 17731 7251 17737
rect 7193 17728 7205 17731
rect 7156 17700 7205 17728
rect 7156 17688 7162 17700
rect 7193 17697 7205 17700
rect 7239 17697 7251 17731
rect 7193 17691 7251 17697
rect 8570 17688 8576 17740
rect 8628 17688 8634 17740
rect 8662 17688 8668 17740
rect 8720 17688 8726 17740
rect 8864 17728 8892 17768
rect 9674 17756 9680 17768
rect 9732 17756 9738 17808
rect 9784 17796 9812 17836
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10045 17867 10103 17873
rect 10045 17864 10057 17867
rect 9916 17836 10057 17864
rect 9916 17824 9922 17836
rect 10045 17833 10057 17836
rect 10091 17833 10103 17867
rect 10045 17827 10103 17833
rect 9784 17768 9996 17796
rect 8772 17700 8892 17728
rect 8932 17731 8990 17737
rect 8772 17660 8800 17700
rect 8932 17697 8944 17731
rect 8978 17728 8990 17731
rect 9858 17728 9864 17740
rect 8978 17700 9864 17728
rect 8978 17697 8990 17700
rect 8932 17691 8990 17697
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 6656 17632 8800 17660
rect 9968 17660 9996 17768
rect 10060 17728 10088 17827
rect 10226 17824 10232 17876
rect 10284 17864 10290 17876
rect 10686 17864 10692 17876
rect 10284 17836 10692 17864
rect 10284 17824 10290 17836
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 11146 17864 11152 17876
rect 10827 17836 11152 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11425 17867 11483 17873
rect 11425 17833 11437 17867
rect 11471 17864 11483 17867
rect 11606 17864 11612 17876
rect 11471 17836 11612 17864
rect 11471 17833 11483 17836
rect 11425 17827 11483 17833
rect 11606 17824 11612 17836
rect 11664 17824 11670 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13817 17867 13875 17873
rect 13817 17864 13829 17867
rect 12492 17836 13829 17864
rect 12492 17824 12498 17836
rect 13817 17833 13829 17836
rect 13863 17833 13875 17867
rect 13817 17827 13875 17833
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 15010 17864 15016 17876
rect 14231 17836 15016 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 15930 17824 15936 17876
rect 15988 17864 15994 17876
rect 16117 17867 16175 17873
rect 16117 17864 16129 17867
rect 15988 17836 16129 17864
rect 15988 17824 15994 17836
rect 16117 17833 16129 17836
rect 16163 17833 16175 17867
rect 16117 17827 16175 17833
rect 17037 17867 17095 17873
rect 17037 17833 17049 17867
rect 17083 17864 17095 17867
rect 17126 17864 17132 17876
rect 17083 17836 17132 17864
rect 17083 17833 17095 17836
rect 17037 17827 17095 17833
rect 17126 17824 17132 17836
rect 17184 17824 17190 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19392 17836 19717 17864
rect 19392 17824 19398 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 21085 17867 21143 17873
rect 21085 17833 21097 17867
rect 21131 17864 21143 17867
rect 23934 17864 23940 17876
rect 21131 17836 23152 17864
rect 21131 17833 21143 17836
rect 21085 17827 21143 17833
rect 12710 17796 12716 17808
rect 11992 17768 12716 17796
rect 10060 17700 10272 17728
rect 10042 17660 10048 17672
rect 9968 17632 10048 17660
rect 10042 17620 10048 17632
rect 10100 17620 10106 17672
rect 10244 17669 10272 17700
rect 11330 17688 11336 17740
rect 11388 17688 11394 17740
rect 11992 17737 12020 17768
rect 12710 17756 12716 17768
rect 12768 17756 12774 17808
rect 13630 17756 13636 17808
rect 13688 17756 13694 17808
rect 16206 17796 16212 17808
rect 15396 17768 16212 17796
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 12233 17731 12291 17737
rect 12233 17728 12245 17731
rect 12124 17700 12245 17728
rect 12124 17688 12130 17700
rect 12233 17697 12245 17700
rect 12279 17697 12291 17731
rect 12233 17691 12291 17697
rect 12526 17688 12532 17740
rect 12584 17728 12590 17740
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 12584 17700 13461 17728
rect 12584 17688 12590 17700
rect 13449 17697 13461 17700
rect 13495 17697 13507 17731
rect 13449 17691 13507 17697
rect 14369 17731 14427 17737
rect 14369 17697 14381 17731
rect 14415 17697 14427 17731
rect 14369 17691 14427 17697
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17660 10287 17663
rect 10594 17660 10600 17672
rect 10275 17632 10600 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 11606 17620 11612 17672
rect 11664 17620 11670 17672
rect 14384 17660 14412 17691
rect 14458 17688 14464 17740
rect 14516 17688 14522 17740
rect 14645 17731 14703 17737
rect 14645 17697 14657 17731
rect 14691 17697 14703 17731
rect 14645 17691 14703 17697
rect 14550 17660 14556 17672
rect 14384 17632 14556 17660
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 5258 17552 5264 17604
rect 5316 17592 5322 17604
rect 7101 17595 7159 17601
rect 7101 17592 7113 17595
rect 5316 17564 7113 17592
rect 5316 17552 5322 17564
rect 7101 17561 7113 17564
rect 7147 17561 7159 17595
rect 7101 17555 7159 17561
rect 10502 17552 10508 17604
rect 10560 17592 10566 17604
rect 11624 17592 11652 17620
rect 10560 17564 11652 17592
rect 10560 17552 10566 17564
rect 13354 17552 13360 17604
rect 13412 17552 13418 17604
rect 14660 17592 14688 17691
rect 14918 17688 14924 17740
rect 14976 17688 14982 17740
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15396 17737 15424 17768
rect 16206 17756 16212 17768
rect 16264 17756 16270 17808
rect 19426 17796 19432 17808
rect 18892 17768 19432 17796
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 15252 17700 15393 17728
rect 15252 17688 15258 17700
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 15381 17691 15439 17697
rect 15562 17688 15568 17740
rect 15620 17688 15626 17740
rect 15654 17688 15660 17740
rect 15712 17688 15718 17740
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 16022 17728 16028 17740
rect 15979 17700 16028 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 15764 17660 15792 17691
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 16114 17688 16120 17740
rect 16172 17688 16178 17740
rect 16298 17688 16304 17740
rect 16356 17688 16362 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 18414 17728 18420 17740
rect 16623 17700 18420 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 18414 17688 18420 17700
rect 18472 17688 18478 17740
rect 18892 17737 18920 17768
rect 19426 17756 19432 17768
rect 19484 17756 19490 17808
rect 19518 17756 19524 17808
rect 19576 17756 19582 17808
rect 20622 17756 20628 17808
rect 20680 17796 20686 17808
rect 21361 17799 21419 17805
rect 21361 17796 21373 17799
rect 20680 17768 21373 17796
rect 20680 17756 20686 17768
rect 21361 17765 21373 17768
rect 21407 17765 21419 17799
rect 22554 17796 22560 17808
rect 21361 17759 21419 17765
rect 21468 17768 22560 17796
rect 18877 17731 18935 17737
rect 18877 17697 18889 17731
rect 18923 17697 18935 17731
rect 18877 17691 18935 17697
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 15764 17632 16405 17660
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16758 17660 16764 17672
rect 16715 17632 16764 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 18892 17660 18920 17691
rect 19058 17688 19064 17740
rect 19116 17688 19122 17740
rect 19153 17731 19211 17737
rect 19153 17697 19165 17731
rect 19199 17697 19211 17731
rect 19153 17691 19211 17697
rect 18196 17632 18920 17660
rect 18196 17620 18202 17632
rect 18966 17620 18972 17672
rect 19024 17660 19030 17672
rect 19168 17660 19196 17691
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19610 17728 19616 17740
rect 19300 17700 19616 17728
rect 19300 17688 19306 17700
rect 19610 17688 19616 17700
rect 19668 17688 19674 17740
rect 19702 17688 19708 17740
rect 19760 17728 19766 17740
rect 19797 17731 19855 17737
rect 19797 17728 19809 17731
rect 19760 17700 19809 17728
rect 19760 17688 19766 17700
rect 19797 17697 19809 17700
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 20714 17688 20720 17740
rect 20772 17688 20778 17740
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21082 17728 21088 17740
rect 20947 17700 21088 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21082 17688 21088 17700
rect 21140 17728 21146 17740
rect 21468 17728 21496 17768
rect 22554 17756 22560 17768
rect 22612 17756 22618 17808
rect 21140 17700 21496 17728
rect 21140 17688 21146 17700
rect 22186 17688 22192 17740
rect 22244 17688 22250 17740
rect 23124 17737 23152 17836
rect 23308 17836 23940 17864
rect 23308 17737 23336 17836
rect 23934 17824 23940 17836
rect 23992 17824 23998 17876
rect 24029 17867 24087 17873
rect 24029 17833 24041 17867
rect 24075 17864 24087 17867
rect 24118 17864 24124 17876
rect 24075 17836 24124 17864
rect 24075 17833 24087 17836
rect 24029 17827 24087 17833
rect 24118 17824 24124 17836
rect 24176 17824 24182 17876
rect 24854 17824 24860 17876
rect 24912 17864 24918 17876
rect 25225 17867 25283 17873
rect 25225 17864 25237 17867
rect 24912 17836 25237 17864
rect 24912 17824 24918 17836
rect 25225 17833 25237 17836
rect 25271 17833 25283 17867
rect 25593 17867 25651 17873
rect 25593 17864 25605 17867
rect 25225 17827 25283 17833
rect 25332 17836 25605 17864
rect 23400 17768 24164 17796
rect 23400 17737 23428 17768
rect 24136 17740 24164 17768
rect 24228 17768 24808 17796
rect 22649 17731 22707 17737
rect 22649 17697 22661 17731
rect 22695 17697 22707 17731
rect 22649 17691 22707 17697
rect 23109 17731 23167 17737
rect 23109 17697 23121 17731
rect 23155 17697 23167 17731
rect 23109 17691 23167 17697
rect 23293 17731 23351 17737
rect 23293 17697 23305 17731
rect 23339 17697 23351 17731
rect 23293 17691 23351 17697
rect 23385 17731 23443 17737
rect 23385 17697 23397 17731
rect 23431 17697 23443 17731
rect 23385 17691 23443 17697
rect 23477 17731 23535 17737
rect 23477 17697 23489 17731
rect 23523 17703 23612 17731
rect 23523 17697 23535 17703
rect 23477 17691 23535 17697
rect 20806 17660 20812 17672
rect 19024 17632 20812 17660
rect 19024 17620 19030 17632
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 22465 17663 22523 17669
rect 22465 17629 22477 17663
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 21266 17592 21272 17604
rect 14660 17564 21272 17592
rect 21266 17552 21272 17564
rect 21324 17552 21330 17604
rect 22480 17592 22508 17623
rect 22554 17620 22560 17672
rect 22612 17660 22618 17672
rect 22664 17660 22692 17691
rect 23584 17660 23612 17703
rect 24118 17688 24124 17740
rect 24176 17688 24182 17740
rect 24228 17660 24256 17768
rect 24780 17740 24808 17768
rect 24305 17731 24363 17737
rect 24305 17697 24317 17731
rect 24351 17697 24363 17731
rect 24305 17691 24363 17697
rect 22612 17632 24256 17660
rect 24320 17660 24348 17691
rect 24394 17688 24400 17740
rect 24452 17688 24458 17740
rect 24489 17731 24547 17737
rect 24489 17697 24501 17731
rect 24535 17697 24547 17731
rect 24489 17691 24547 17697
rect 24320 17632 24440 17660
rect 22612 17620 22618 17632
rect 24302 17592 24308 17604
rect 22480 17564 24308 17592
rect 24302 17552 24308 17564
rect 24360 17552 24366 17604
rect 4338 17524 4344 17536
rect 4265 17496 4344 17524
rect 4338 17484 4344 17496
rect 4396 17484 4402 17536
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5592 17496 5825 17524
rect 5592 17484 5598 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 5813 17487 5871 17493
rect 6270 17484 6276 17536
rect 6328 17524 6334 17536
rect 6914 17524 6920 17536
rect 6328 17496 6920 17524
rect 6328 17484 6334 17496
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 10965 17527 11023 17533
rect 10965 17524 10977 17527
rect 9640 17496 10977 17524
rect 9640 17484 9646 17496
rect 10965 17493 10977 17496
rect 11011 17493 11023 17527
rect 10965 17487 11023 17493
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 13372 17524 13400 17552
rect 11388 17496 13400 17524
rect 11388 17484 11394 17496
rect 14366 17484 14372 17536
rect 14424 17524 14430 17536
rect 14829 17527 14887 17533
rect 14829 17524 14841 17527
rect 14424 17496 14841 17524
rect 14424 17484 14430 17496
rect 14829 17493 14841 17496
rect 14875 17493 14887 17527
rect 14829 17487 14887 17493
rect 14918 17484 14924 17536
rect 14976 17524 14982 17536
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 14976 17496 15025 17524
rect 14976 17484 14982 17496
rect 15013 17493 15025 17496
rect 15059 17493 15071 17527
rect 15013 17487 15071 17493
rect 15194 17484 15200 17536
rect 15252 17484 15258 17536
rect 18690 17484 18696 17536
rect 18748 17524 18754 17536
rect 22002 17524 22008 17536
rect 18748 17496 22008 17524
rect 18748 17484 18754 17496
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 22922 17484 22928 17536
rect 22980 17524 22986 17536
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 22980 17496 23029 17524
rect 22980 17484 22986 17496
rect 23017 17493 23029 17496
rect 23063 17493 23075 17527
rect 23017 17487 23075 17493
rect 23198 17484 23204 17536
rect 23256 17524 23262 17536
rect 23753 17527 23811 17533
rect 23753 17524 23765 17527
rect 23256 17496 23765 17524
rect 23256 17484 23262 17496
rect 23753 17493 23765 17496
rect 23799 17493 23811 17527
rect 24412 17524 24440 17632
rect 24504 17592 24532 17691
rect 24670 17688 24676 17740
rect 24728 17688 24734 17740
rect 24762 17688 24768 17740
rect 24820 17728 24826 17740
rect 25133 17731 25191 17737
rect 25133 17728 25145 17731
rect 24820 17700 25145 17728
rect 24820 17688 24826 17700
rect 25133 17697 25145 17700
rect 25179 17697 25191 17731
rect 25332 17728 25360 17836
rect 25593 17833 25605 17836
rect 25639 17833 25651 17867
rect 25593 17827 25651 17833
rect 25976 17836 26556 17864
rect 25406 17756 25412 17808
rect 25464 17796 25470 17808
rect 25976 17796 26004 17836
rect 25464 17768 26004 17796
rect 25464 17756 25470 17768
rect 25976 17737 26004 17768
rect 26050 17756 26056 17808
rect 26108 17796 26114 17808
rect 26421 17799 26479 17805
rect 26421 17796 26433 17799
rect 26108 17768 26433 17796
rect 26108 17756 26114 17768
rect 26421 17765 26433 17768
rect 26467 17765 26479 17799
rect 26421 17759 26479 17765
rect 25869 17731 25927 17737
rect 25869 17728 25881 17731
rect 25332 17700 25881 17728
rect 25133 17691 25191 17697
rect 25869 17697 25881 17700
rect 25915 17697 25927 17731
rect 25869 17691 25927 17697
rect 25961 17731 26019 17737
rect 25961 17697 25973 17731
rect 26007 17697 26019 17731
rect 25961 17691 26019 17697
rect 26142 17688 26148 17740
rect 26200 17688 26206 17740
rect 26234 17688 26240 17740
rect 26292 17688 26298 17740
rect 26528 17728 26556 17836
rect 26694 17824 26700 17876
rect 26752 17864 26758 17876
rect 27433 17867 27491 17873
rect 27433 17864 27445 17867
rect 26752 17836 27445 17864
rect 26752 17824 26758 17836
rect 27433 17833 27445 17836
rect 27479 17833 27491 17867
rect 28534 17864 28540 17876
rect 27433 17827 27491 17833
rect 27724 17836 28540 17864
rect 27249 17799 27307 17805
rect 27249 17765 27261 17799
rect 27295 17796 27307 17799
rect 27338 17796 27344 17808
rect 27295 17768 27344 17796
rect 27295 17765 27307 17768
rect 27249 17759 27307 17765
rect 27338 17756 27344 17768
rect 27396 17756 27402 17808
rect 27724 17796 27752 17836
rect 28534 17824 28540 17836
rect 28592 17864 28598 17876
rect 28592 17836 28672 17864
rect 28592 17824 28598 17836
rect 28074 17796 28080 17808
rect 27448 17768 27752 17796
rect 27448 17728 27476 17768
rect 27724 17737 27752 17768
rect 27908 17768 28080 17796
rect 27908 17737 27936 17768
rect 28074 17756 28080 17768
rect 28132 17756 28138 17808
rect 28644 17796 28672 17836
rect 28994 17824 29000 17876
rect 29052 17824 29058 17876
rect 29454 17824 29460 17876
rect 29512 17864 29518 17876
rect 29549 17867 29607 17873
rect 29549 17864 29561 17867
rect 29512 17836 29561 17864
rect 29512 17824 29518 17836
rect 29549 17833 29561 17836
rect 29595 17833 29607 17867
rect 29549 17827 29607 17833
rect 29641 17867 29699 17873
rect 29641 17833 29653 17867
rect 29687 17864 29699 17867
rect 30282 17864 30288 17876
rect 29687 17836 30288 17864
rect 29687 17833 29699 17836
rect 29641 17827 29699 17833
rect 30282 17824 30288 17836
rect 30340 17824 30346 17876
rect 28644 17768 28994 17796
rect 26528 17700 27476 17728
rect 27617 17731 27675 17737
rect 27617 17697 27629 17731
rect 27663 17697 27675 17731
rect 27617 17691 27675 17697
rect 27709 17731 27767 17737
rect 27709 17697 27721 17731
rect 27755 17697 27767 17731
rect 27709 17691 27767 17697
rect 27893 17731 27951 17737
rect 27893 17697 27905 17731
rect 27939 17697 27951 17731
rect 27893 17691 27951 17697
rect 27985 17731 28043 17737
rect 27985 17697 27997 17731
rect 28031 17726 28043 17731
rect 28031 17698 28120 17726
rect 28031 17697 28043 17698
rect 27985 17691 28043 17697
rect 24946 17620 24952 17672
rect 25004 17620 25010 17672
rect 25774 17620 25780 17672
rect 25832 17660 25838 17672
rect 27632 17660 27660 17691
rect 25832 17632 27660 17660
rect 25832 17620 25838 17632
rect 28092 17604 28120 17698
rect 28350 17688 28356 17740
rect 28408 17688 28414 17740
rect 28534 17688 28540 17740
rect 28592 17688 28598 17740
rect 28626 17688 28632 17740
rect 28684 17688 28690 17740
rect 28718 17688 28724 17740
rect 28776 17688 28782 17740
rect 28966 17728 28994 17768
rect 29270 17756 29276 17808
rect 29328 17796 29334 17808
rect 30300 17796 30328 17824
rect 29328 17768 30144 17796
rect 30300 17768 30512 17796
rect 29328 17756 29334 17768
rect 30006 17728 30012 17740
rect 28966 17700 30012 17728
rect 30006 17688 30012 17700
rect 30064 17688 30070 17740
rect 30116 17737 30144 17768
rect 30101 17731 30159 17737
rect 30101 17697 30113 17731
rect 30147 17697 30159 17731
rect 30101 17691 30159 17697
rect 30190 17688 30196 17740
rect 30248 17728 30254 17740
rect 30484 17737 30512 17768
rect 30285 17731 30343 17737
rect 30285 17728 30297 17731
rect 30248 17700 30297 17728
rect 30248 17688 30254 17700
rect 30285 17697 30297 17700
rect 30331 17697 30343 17731
rect 30285 17691 30343 17697
rect 30377 17731 30435 17737
rect 30377 17697 30389 17731
rect 30423 17697 30435 17731
rect 30377 17691 30435 17697
rect 30469 17731 30527 17737
rect 30469 17697 30481 17731
rect 30515 17697 30527 17731
rect 30469 17691 30527 17697
rect 28166 17620 28172 17672
rect 28224 17660 28230 17672
rect 28736 17660 28764 17688
rect 28224 17632 28764 17660
rect 29457 17663 29515 17669
rect 28224 17620 28230 17632
rect 29457 17629 29469 17663
rect 29503 17660 29515 17663
rect 29546 17660 29552 17672
rect 29503 17632 29552 17660
rect 29503 17629 29515 17632
rect 29457 17623 29515 17629
rect 29546 17620 29552 17632
rect 29604 17620 29610 17672
rect 25685 17595 25743 17601
rect 25685 17592 25697 17595
rect 24504 17564 25697 17592
rect 25685 17561 25697 17564
rect 25731 17561 25743 17595
rect 25685 17555 25743 17561
rect 28074 17552 28080 17604
rect 28132 17592 28138 17604
rect 28442 17592 28448 17604
rect 28132 17564 28448 17592
rect 28132 17552 28138 17564
rect 28442 17552 28448 17564
rect 28500 17552 28506 17604
rect 28718 17552 28724 17604
rect 28776 17592 28782 17604
rect 30392 17592 30420 17691
rect 28776 17564 30420 17592
rect 28776 17552 28782 17564
rect 25222 17524 25228 17536
rect 24412 17496 25228 17524
rect 23753 17487 23811 17493
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 27614 17484 27620 17536
rect 27672 17524 27678 17536
rect 28736 17524 28764 17552
rect 27672 17496 28764 17524
rect 30009 17527 30067 17533
rect 27672 17484 27678 17496
rect 30009 17493 30021 17527
rect 30055 17524 30067 17527
rect 30466 17524 30472 17536
rect 30055 17496 30472 17524
rect 30055 17493 30067 17496
rect 30009 17487 30067 17493
rect 30466 17484 30472 17496
rect 30524 17484 30530 17536
rect 30558 17484 30564 17536
rect 30616 17524 30622 17536
rect 30745 17527 30803 17533
rect 30745 17524 30757 17527
rect 30616 17496 30757 17524
rect 30616 17484 30622 17496
rect 30745 17493 30757 17496
rect 30791 17493 30803 17527
rect 30745 17487 30803 17493
rect 552 17434 31648 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 11436 17434
rect 11488 17382 11500 17434
rect 11552 17382 11564 17434
rect 11616 17382 11628 17434
rect 11680 17382 11692 17434
rect 11744 17382 19210 17434
rect 19262 17382 19274 17434
rect 19326 17382 19338 17434
rect 19390 17382 19402 17434
rect 19454 17382 19466 17434
rect 19518 17382 26984 17434
rect 27036 17382 27048 17434
rect 27100 17382 27112 17434
rect 27164 17382 27176 17434
rect 27228 17382 27240 17434
rect 27292 17382 31648 17434
rect 552 17360 31648 17382
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 3697 17323 3755 17329
rect 3697 17320 3709 17323
rect 3568 17292 3709 17320
rect 3568 17280 3574 17292
rect 3697 17289 3709 17292
rect 3743 17289 3755 17323
rect 3697 17283 3755 17289
rect 3789 17323 3847 17329
rect 3789 17289 3801 17323
rect 3835 17320 3847 17323
rect 4062 17320 4068 17332
rect 3835 17292 4068 17320
rect 3835 17289 3847 17292
rect 3789 17283 3847 17289
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4709 17323 4767 17329
rect 4709 17289 4721 17323
rect 4755 17320 4767 17323
rect 5166 17320 5172 17332
rect 4755 17292 5172 17320
rect 4755 17289 4767 17292
rect 4709 17283 4767 17289
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 5994 17320 6000 17332
rect 5951 17292 6000 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 5994 17280 6000 17292
rect 6052 17320 6058 17332
rect 6052 17292 6592 17320
rect 6052 17280 6058 17292
rect 2777 17255 2835 17261
rect 2777 17221 2789 17255
rect 2823 17252 2835 17255
rect 3878 17252 3884 17264
rect 2823 17224 3884 17252
rect 2823 17221 2835 17224
rect 2777 17215 2835 17221
rect 1213 17187 1271 17193
rect 1213 17153 1225 17187
rect 1259 17184 1271 17187
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 1259 17156 1409 17184
rect 1259 17153 1271 17156
rect 1213 17147 1271 17153
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 2682 17144 2688 17196
rect 2740 17184 2746 17196
rect 2792 17184 2820 17215
rect 3878 17212 3884 17224
rect 3936 17212 3942 17264
rect 4525 17255 4583 17261
rect 4525 17221 4537 17255
rect 4571 17252 4583 17255
rect 6089 17255 6147 17261
rect 6089 17252 6101 17255
rect 4571 17224 6101 17252
rect 4571 17221 4583 17224
rect 4525 17215 4583 17221
rect 6089 17221 6101 17224
rect 6135 17221 6147 17255
rect 6089 17215 6147 17221
rect 6362 17212 6368 17264
rect 6420 17252 6426 17264
rect 6420 17224 6500 17252
rect 6420 17212 6426 17224
rect 2740 17156 2820 17184
rect 3605 17187 3663 17193
rect 2740 17144 2746 17156
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 3651 17156 4629 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 4617 17153 4629 17156
rect 4663 17184 4675 17187
rect 5077 17187 5135 17193
rect 5077 17184 5089 17187
rect 4663 17156 5089 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 5077 17153 5089 17156
rect 5123 17153 5135 17187
rect 5721 17187 5779 17193
rect 5077 17147 5135 17153
rect 5184 17156 5580 17184
rect 1305 17119 1363 17125
rect 1305 17085 1317 17119
rect 1351 17116 1363 17119
rect 1664 17119 1722 17125
rect 1351 17088 1440 17116
rect 1351 17085 1363 17088
rect 1305 17079 1363 17085
rect 1412 17060 1440 17088
rect 1664 17085 1676 17119
rect 1710 17116 1722 17119
rect 2406 17116 2412 17128
rect 1710 17088 2412 17116
rect 1710 17085 1722 17088
rect 1664 17079 1722 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 4154 17116 4160 17128
rect 4111 17088 4160 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4154 17076 4160 17088
rect 4212 17116 4218 17128
rect 4522 17116 4528 17128
rect 4212 17088 4528 17116
rect 4212 17076 4218 17088
rect 4522 17076 4528 17088
rect 4580 17076 4586 17128
rect 4798 17076 4804 17128
rect 4856 17076 4862 17128
rect 4982 17076 4988 17128
rect 5040 17076 5046 17128
rect 1394 17008 1400 17060
rect 1452 17008 1458 17060
rect 2682 17008 2688 17060
rect 2740 17048 2746 17060
rect 4249 17051 4307 17057
rect 4249 17048 4261 17051
rect 2740 17020 4261 17048
rect 2740 17008 2746 17020
rect 4249 17017 4261 17020
rect 4295 17017 4307 17051
rect 4249 17011 4307 17017
rect 4706 17008 4712 17060
rect 4764 17048 4770 17060
rect 5184 17048 5212 17156
rect 5258 17076 5264 17128
rect 5316 17076 5322 17128
rect 5442 17076 5448 17128
rect 5500 17076 5506 17128
rect 5552 17116 5580 17156
rect 5721 17153 5733 17187
rect 5767 17184 5779 17187
rect 6178 17184 6184 17196
rect 5767 17156 6184 17184
rect 5767 17153 5779 17156
rect 5721 17147 5779 17153
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 6472 17193 6500 17224
rect 6457 17187 6515 17193
rect 6457 17153 6469 17187
rect 6503 17153 6515 17187
rect 6457 17147 6515 17153
rect 5813 17119 5871 17125
rect 5813 17116 5825 17119
rect 5552 17088 5825 17116
rect 5813 17085 5825 17088
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 5994 17076 6000 17128
rect 6052 17076 6058 17128
rect 6086 17076 6092 17128
rect 6144 17076 6150 17128
rect 6270 17076 6276 17128
rect 6328 17076 6334 17128
rect 6564 17125 6592 17292
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 10873 17323 10931 17329
rect 8352 17292 10425 17320
rect 8352 17280 8358 17292
rect 9769 17255 9827 17261
rect 9769 17221 9781 17255
rect 9815 17221 9827 17255
rect 9769 17215 9827 17221
rect 8294 17184 8300 17196
rect 8036 17156 8300 17184
rect 8036 17128 8064 17156
rect 8294 17144 8300 17156
rect 8352 17144 8358 17196
rect 9784 17184 9812 17215
rect 9858 17212 9864 17264
rect 9916 17212 9922 17264
rect 10397 17252 10425 17292
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 11330 17320 11336 17332
rect 10919 17292 11336 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 11790 17280 11796 17332
rect 11848 17280 11854 17332
rect 14001 17323 14059 17329
rect 14001 17320 14013 17323
rect 12176 17292 14013 17320
rect 11146 17252 11152 17264
rect 10397 17224 11152 17252
rect 11146 17212 11152 17224
rect 11204 17212 11210 17264
rect 9950 17184 9956 17196
rect 9784 17156 9956 17184
rect 9950 17144 9956 17156
rect 10008 17184 10014 17196
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10008 17156 10701 17184
rect 10008 17144 10014 17156
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 12176 17184 12204 17292
rect 14001 17289 14013 17292
rect 14047 17289 14059 17323
rect 15930 17320 15936 17332
rect 14001 17283 14059 17289
rect 14292 17292 15936 17320
rect 10689 17147 10747 17153
rect 10796 17156 12204 17184
rect 6365 17119 6423 17125
rect 6365 17085 6377 17119
rect 6411 17085 6423 17119
rect 6365 17079 6423 17085
rect 6549 17119 6607 17125
rect 6549 17085 6561 17119
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 5626 17057 5632 17060
rect 4764 17020 5212 17048
rect 5353 17051 5411 17057
rect 4764 17008 4770 17020
rect 5353 17017 5365 17051
rect 5399 17048 5411 17051
rect 5583 17051 5632 17057
rect 5399 17020 5488 17048
rect 5399 17017 5411 17020
rect 5353 17011 5411 17017
rect 3326 16940 3332 16992
rect 3384 16940 3390 16992
rect 3878 16940 3884 16992
rect 3936 16980 3942 16992
rect 3973 16983 4031 16989
rect 3973 16980 3985 16983
rect 3936 16952 3985 16980
rect 3936 16940 3942 16952
rect 3973 16949 3985 16952
rect 4019 16949 4031 16983
rect 3973 16943 4031 16949
rect 4338 16940 4344 16992
rect 4396 16980 4402 16992
rect 5166 16980 5172 16992
rect 4396 16952 5172 16980
rect 4396 16940 4402 16952
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 5460 16980 5488 17020
rect 5583 17017 5595 17051
rect 5629 17017 5632 17051
rect 5583 17011 5632 17017
rect 5626 17008 5632 17011
rect 5684 17048 5690 17060
rect 5902 17048 5908 17060
rect 5684 17020 5908 17048
rect 5684 17008 5690 17020
rect 5902 17008 5908 17020
rect 5960 17008 5966 17060
rect 6380 17048 6408 17079
rect 8018 17076 8024 17128
rect 8076 17076 8082 17128
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17116 8171 17119
rect 8389 17119 8447 17125
rect 8389 17116 8401 17119
rect 8159 17088 8401 17116
rect 8159 17085 8171 17088
rect 8113 17079 8171 17085
rect 8389 17085 8401 17088
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 8656 17119 8714 17125
rect 8656 17085 8668 17119
rect 8702 17116 8714 17119
rect 10042 17116 10048 17128
rect 8702 17088 10048 17116
rect 8702 17085 8714 17088
rect 8656 17079 8714 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17085 10195 17119
rect 10137 17079 10195 17085
rect 6730 17048 6736 17060
rect 6380 17020 6736 17048
rect 6380 16980 6408 17020
rect 6730 17008 6736 17020
rect 6788 17008 6794 17060
rect 9398 17008 9404 17060
rect 9456 17048 9462 17060
rect 10152 17048 10180 17079
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 10318 17076 10324 17128
rect 10376 17076 10382 17128
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 10468 17088 10517 17116
rect 10468 17076 10474 17088
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 10594 17076 10600 17128
rect 10652 17076 10658 17128
rect 10796 17048 10824 17156
rect 10873 17119 10931 17125
rect 10873 17085 10885 17119
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 9456 17020 10824 17048
rect 10888 17048 10916 17079
rect 11146 17076 11152 17128
rect 11204 17076 11210 17128
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 12906 17119 12964 17125
rect 12906 17116 12918 17119
rect 12676 17088 12918 17116
rect 12676 17076 12682 17088
rect 12906 17085 12918 17088
rect 12952 17085 12964 17119
rect 12906 17079 12964 17085
rect 13173 17119 13231 17125
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13633 17119 13691 17125
rect 13633 17116 13645 17119
rect 13219 17088 13645 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 13633 17085 13645 17088
rect 13679 17085 13691 17119
rect 13633 17079 13691 17085
rect 13722 17076 13728 17128
rect 13780 17076 13786 17128
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 13906 17116 13912 17128
rect 13863 17088 13912 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 11698 17048 11704 17060
rect 10888 17020 11704 17048
rect 9456 17008 9462 17020
rect 11698 17008 11704 17020
rect 11756 17008 11762 17060
rect 14016 17048 14044 17283
rect 14292 17252 14320 17292
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16301 17323 16359 17329
rect 16301 17320 16313 17323
rect 16264 17292 16313 17320
rect 16264 17280 16270 17292
rect 16301 17289 16313 17292
rect 16347 17289 16359 17323
rect 16301 17283 16359 17289
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 23658 17320 23664 17332
rect 20772 17292 23664 17320
rect 20772 17280 20778 17292
rect 23658 17280 23664 17292
rect 23716 17280 23722 17332
rect 24026 17280 24032 17332
rect 24084 17320 24090 17332
rect 25590 17320 25596 17332
rect 24084 17292 25596 17320
rect 24084 17280 24090 17292
rect 25590 17280 25596 17292
rect 25648 17280 25654 17332
rect 25685 17323 25743 17329
rect 25685 17289 25697 17323
rect 25731 17320 25743 17323
rect 25774 17320 25780 17332
rect 25731 17292 25780 17320
rect 25731 17289 25743 17292
rect 25685 17283 25743 17289
rect 25774 17280 25780 17292
rect 25832 17280 25838 17332
rect 26142 17280 26148 17332
rect 26200 17320 26206 17332
rect 27249 17323 27307 17329
rect 27249 17320 27261 17323
rect 26200 17292 27261 17320
rect 26200 17280 26206 17292
rect 27249 17289 27261 17292
rect 27295 17289 27307 17323
rect 27249 17283 27307 17289
rect 28350 17280 28356 17332
rect 28408 17320 28414 17332
rect 28813 17323 28871 17329
rect 28813 17320 28825 17323
rect 28408 17292 28825 17320
rect 28408 17280 28414 17292
rect 28813 17289 28825 17292
rect 28859 17289 28871 17323
rect 28813 17283 28871 17289
rect 30374 17280 30380 17332
rect 30432 17320 30438 17332
rect 31021 17323 31079 17329
rect 31021 17320 31033 17323
rect 30432 17292 31033 17320
rect 30432 17280 30438 17292
rect 31021 17289 31033 17292
rect 31067 17289 31079 17323
rect 31021 17283 31079 17289
rect 14200 17224 14320 17252
rect 14200 17128 14228 17224
rect 14826 17212 14832 17264
rect 14884 17212 14890 17264
rect 19426 17252 19432 17264
rect 18248 17224 19432 17252
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 14332 17156 14504 17184
rect 14332 17144 14338 17156
rect 14182 17076 14188 17128
rect 14240 17076 14246 17128
rect 14366 17076 14372 17128
rect 14424 17076 14430 17128
rect 14476 17125 14504 17156
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 14461 17119 14519 17125
rect 14461 17085 14473 17119
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 14568 17048 14596 17079
rect 14918 17076 14924 17128
rect 14976 17076 14982 17128
rect 16298 17116 16304 17128
rect 15028 17088 16304 17116
rect 15028 17048 15056 17088
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17116 16727 17119
rect 16942 17116 16948 17128
rect 16715 17088 16948 17116
rect 16715 17085 16727 17088
rect 16669 17079 16727 17085
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18248 17125 18276 17224
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 20254 17212 20260 17264
rect 20312 17212 20318 17264
rect 29546 17252 29552 17264
rect 26160 17224 29552 17252
rect 26160 17196 26188 17224
rect 29546 17212 29552 17224
rect 29604 17212 29610 17264
rect 30282 17212 30288 17264
rect 30340 17252 30346 17264
rect 30340 17224 30420 17252
rect 30340 17212 30346 17224
rect 18598 17144 18604 17196
rect 18656 17184 18662 17196
rect 18656 17156 19748 17184
rect 18656 17144 18662 17156
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17828 17088 18061 17116
rect 17828 17076 17834 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17085 18291 17119
rect 18233 17079 18291 17085
rect 14016 17020 15056 17048
rect 15930 17008 15936 17060
rect 15988 17048 15994 17060
rect 15988 17020 16436 17048
rect 15988 17008 15994 17020
rect 5460 16952 6408 16980
rect 11057 16983 11115 16989
rect 11057 16949 11069 16983
rect 11103 16980 11115 16983
rect 11606 16980 11612 16992
rect 11103 16952 11612 16980
rect 11103 16949 11115 16952
rect 11057 16943 11115 16949
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 16408 16980 16436 17020
rect 16758 17008 16764 17060
rect 16816 17048 16822 17060
rect 18248 17048 18276 17079
rect 18690 17076 18696 17128
rect 18748 17076 18754 17128
rect 18785 17119 18843 17125
rect 18785 17085 18797 17119
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 16816 17020 18276 17048
rect 18800 17048 18828 17079
rect 18966 17076 18972 17128
rect 19024 17076 19030 17128
rect 19058 17076 19064 17128
rect 19116 17076 19122 17128
rect 19610 17076 19616 17128
rect 19668 17076 19674 17128
rect 19150 17048 19156 17060
rect 18800 17020 19156 17048
rect 16816 17008 16822 17020
rect 19150 17008 19156 17020
rect 19208 17008 19214 17060
rect 19245 17051 19303 17057
rect 19245 17017 19257 17051
rect 19291 17048 19303 17051
rect 19291 17020 19656 17048
rect 19291 17017 19303 17020
rect 19245 17011 19303 17017
rect 19628 16992 19656 17020
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16408 16952 16865 16980
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 16853 16943 16911 16949
rect 18233 16983 18291 16989
rect 18233 16949 18245 16983
rect 18279 16980 18291 16983
rect 18874 16980 18880 16992
rect 18279 16952 18880 16980
rect 18279 16949 18291 16952
rect 18233 16943 18291 16949
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 19426 16940 19432 16992
rect 19484 16940 19490 16992
rect 19610 16940 19616 16992
rect 19668 16940 19674 16992
rect 19720 16980 19748 17156
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 21082 17193 21088 17196
rect 21060 17187 21088 17193
rect 21060 17153 21072 17187
rect 21060 17147 21088 17153
rect 21082 17144 21088 17147
rect 21140 17144 21146 17196
rect 21450 17144 21456 17196
rect 21508 17144 21514 17196
rect 21913 17187 21971 17193
rect 21913 17153 21925 17187
rect 21959 17184 21971 17187
rect 22554 17184 22560 17196
rect 21959 17156 22560 17184
rect 21959 17153 21971 17156
rect 21913 17147 21971 17153
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17184 23627 17187
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 23615 17156 23949 17184
rect 23615 17153 23627 17156
rect 23569 17147 23627 17153
rect 23937 17153 23949 17156
rect 23983 17153 23995 17187
rect 23937 17147 23995 17153
rect 24946 17144 24952 17196
rect 25004 17184 25010 17196
rect 25133 17187 25191 17193
rect 25133 17184 25145 17187
rect 25004 17156 25145 17184
rect 25004 17144 25010 17156
rect 25133 17153 25145 17156
rect 25179 17184 25191 17187
rect 25958 17184 25964 17196
rect 25179 17156 25964 17184
rect 25179 17153 25191 17156
rect 25133 17147 25191 17153
rect 25958 17144 25964 17156
rect 26016 17184 26022 17196
rect 26142 17184 26148 17196
rect 26016 17156 26148 17184
rect 26016 17144 26022 17156
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 26786 17144 26792 17196
rect 26844 17184 26850 17196
rect 27982 17184 27988 17196
rect 26844 17156 27988 17184
rect 26844 17144 26850 17156
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 19852 17088 19993 17116
rect 19852 17076 19858 17088
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 21174 17076 21180 17128
rect 21232 17076 21238 17128
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17116 22155 17119
rect 22143 17088 22232 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 20073 17051 20131 17057
rect 20073 17017 20085 17051
rect 20119 17048 20131 17051
rect 20346 17048 20352 17060
rect 20119 17020 20352 17048
rect 20119 17017 20131 17020
rect 20073 17011 20131 17017
rect 20346 17008 20352 17020
rect 20404 17008 20410 17060
rect 21450 16980 21456 16992
rect 19720 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 22204 16989 22232 17088
rect 23290 17076 23296 17128
rect 23348 17125 23354 17128
rect 23348 17116 23360 17125
rect 23348 17088 23393 17116
rect 23348 17079 23360 17088
rect 23348 17076 23354 17079
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 23845 17119 23903 17125
rect 23845 17116 23857 17119
rect 23532 17088 23857 17116
rect 23532 17076 23538 17088
rect 23845 17085 23857 17088
rect 23891 17085 23903 17119
rect 23845 17079 23903 17085
rect 24213 17119 24271 17125
rect 24213 17085 24225 17119
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 24397 17119 24455 17125
rect 24397 17085 24409 17119
rect 24443 17085 24455 17119
rect 24397 17079 24455 17085
rect 22189 16983 22247 16989
rect 22189 16949 22201 16983
rect 22235 16980 22247 16983
rect 22278 16980 22284 16992
rect 22235 16952 22284 16980
rect 22235 16949 22247 16952
rect 22189 16943 22247 16949
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 24228 16980 24256 17079
rect 24412 17048 24440 17079
rect 24486 17076 24492 17128
rect 24544 17076 24550 17128
rect 24581 17119 24639 17125
rect 24581 17085 24593 17119
rect 24627 17116 24639 17119
rect 24762 17116 24768 17128
rect 24627 17088 24768 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 24762 17076 24768 17088
rect 24820 17076 24826 17128
rect 25317 17119 25375 17125
rect 25317 17085 25329 17119
rect 25363 17116 25375 17119
rect 25866 17116 25872 17128
rect 25363 17088 25872 17116
rect 25363 17085 25375 17088
rect 25317 17079 25375 17085
rect 25866 17076 25872 17088
rect 25924 17076 25930 17128
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27338 17116 27344 17128
rect 27203 17088 27344 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 27338 17076 27344 17088
rect 27396 17076 27402 17128
rect 27540 17125 27568 17156
rect 27982 17144 27988 17156
rect 28040 17144 28046 17196
rect 28810 17184 28816 17196
rect 28276 17156 28816 17184
rect 27525 17119 27583 17125
rect 27525 17085 27537 17119
rect 27571 17085 27583 17119
rect 27525 17079 27583 17085
rect 27614 17076 27620 17128
rect 27672 17076 27678 17128
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17085 27767 17119
rect 27709 17079 27767 17085
rect 25130 17048 25136 17060
rect 24412 17020 25136 17048
rect 25130 17008 25136 17020
rect 25188 17008 25194 17060
rect 25590 17008 25596 17060
rect 25648 17048 25654 17060
rect 27724 17048 27752 17079
rect 27890 17076 27896 17128
rect 27948 17076 27954 17128
rect 25648 17020 27752 17048
rect 25648 17008 25654 17020
rect 24670 16980 24676 16992
rect 24228 16952 24676 16980
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 24854 16940 24860 16992
rect 24912 16940 24918 16992
rect 25222 16940 25228 16992
rect 25280 16940 25286 16992
rect 27724 16980 27752 17020
rect 27982 17008 27988 17060
rect 28040 17008 28046 17060
rect 28166 17008 28172 17060
rect 28224 17008 28230 17060
rect 28276 16980 28304 17156
rect 28810 17144 28816 17156
rect 28868 17184 28874 17196
rect 30190 17184 30196 17196
rect 28868 17156 30196 17184
rect 28868 17144 28874 17156
rect 30190 17144 30196 17156
rect 30248 17144 30254 17196
rect 30392 17193 30420 17224
rect 30466 17212 30472 17264
rect 30524 17212 30530 17264
rect 30377 17187 30435 17193
rect 30377 17153 30389 17187
rect 30423 17153 30435 17187
rect 30484 17184 30512 17212
rect 30484 17156 30880 17184
rect 30377 17147 30435 17153
rect 28353 17119 28411 17125
rect 28353 17085 28365 17119
rect 28399 17116 28411 17119
rect 28902 17116 28908 17128
rect 28399 17088 28908 17116
rect 28399 17085 28411 17088
rect 28353 17079 28411 17085
rect 28902 17076 28908 17088
rect 28960 17076 28966 17128
rect 28997 17119 29055 17125
rect 28997 17085 29009 17119
rect 29043 17116 29055 17119
rect 29086 17116 29092 17128
rect 29043 17088 29092 17116
rect 29043 17085 29055 17088
rect 28997 17079 29055 17085
rect 29086 17076 29092 17088
rect 29144 17076 29150 17128
rect 29178 17076 29184 17128
rect 29236 17076 29242 17128
rect 29270 17076 29276 17128
rect 29328 17076 29334 17128
rect 29365 17119 29423 17125
rect 29365 17085 29377 17119
rect 29411 17116 29423 17119
rect 29733 17119 29791 17125
rect 29733 17116 29745 17119
rect 29411 17088 29745 17116
rect 29411 17085 29423 17088
rect 29365 17079 29423 17085
rect 29733 17085 29745 17088
rect 29779 17085 29791 17119
rect 30469 17119 30527 17125
rect 30469 17116 30481 17119
rect 29733 17079 29791 17085
rect 29840 17088 30481 17116
rect 28442 17008 28448 17060
rect 28500 17008 28506 17060
rect 28626 17008 28632 17060
rect 28684 17008 28690 17060
rect 29840 17048 29868 17088
rect 30469 17085 30481 17088
rect 30515 17085 30527 17119
rect 30469 17079 30527 17085
rect 30558 17076 30564 17128
rect 30616 17076 30622 17128
rect 30742 17076 30748 17128
rect 30800 17076 30806 17128
rect 30852 17125 30880 17156
rect 30837 17119 30895 17125
rect 30837 17085 30849 17119
rect 30883 17085 30895 17119
rect 30837 17079 30895 17085
rect 31113 17119 31171 17125
rect 31113 17085 31125 17119
rect 31159 17085 31171 17119
rect 31113 17079 31171 17085
rect 28966 17020 29868 17048
rect 27724 16952 28304 16980
rect 28534 16940 28540 16992
rect 28592 16980 28598 16992
rect 28966 16980 28994 17020
rect 30006 17008 30012 17060
rect 30064 17048 30070 17060
rect 31128 17048 31156 17079
rect 30064 17020 31156 17048
rect 30064 17008 30070 17020
rect 28592 16952 28994 16980
rect 29641 16983 29699 16989
rect 28592 16940 28598 16952
rect 29641 16949 29653 16983
rect 29687 16980 29699 16983
rect 30190 16980 30196 16992
rect 29687 16952 30196 16980
rect 29687 16949 29699 16952
rect 29641 16943 29699 16949
rect 30190 16940 30196 16952
rect 30248 16940 30254 16992
rect 31202 16940 31208 16992
rect 31260 16940 31266 16992
rect 552 16890 31648 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 12096 16890
rect 12148 16838 12160 16890
rect 12212 16838 12224 16890
rect 12276 16838 12288 16890
rect 12340 16838 12352 16890
rect 12404 16838 19870 16890
rect 19922 16838 19934 16890
rect 19986 16838 19998 16890
rect 20050 16838 20062 16890
rect 20114 16838 20126 16890
rect 20178 16838 27644 16890
rect 27696 16838 27708 16890
rect 27760 16838 27772 16890
rect 27824 16838 27836 16890
rect 27888 16838 27900 16890
rect 27952 16838 31648 16890
rect 552 16816 31648 16838
rect 3234 16736 3240 16788
rect 3292 16776 3298 16788
rect 4062 16776 4068 16788
rect 3292 16748 4068 16776
rect 3292 16736 3298 16748
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4154 16736 4160 16788
rect 4212 16736 4218 16788
rect 4985 16779 5043 16785
rect 4985 16745 4997 16779
rect 5031 16776 5043 16779
rect 5350 16776 5356 16788
rect 5031 16748 5356 16776
rect 5031 16745 5043 16748
rect 4985 16739 5043 16745
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 6181 16779 6239 16785
rect 6181 16745 6193 16779
rect 6227 16776 6239 16779
rect 6270 16776 6276 16788
rect 6227 16748 6276 16776
rect 6227 16745 6239 16748
rect 6181 16739 6239 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 6457 16779 6515 16785
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 6730 16776 6736 16788
rect 6503 16748 6736 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 2869 16711 2927 16717
rect 2869 16708 2881 16711
rect 2424 16680 2881 16708
rect 2424 16649 2452 16680
rect 2869 16677 2881 16680
rect 2915 16677 2927 16711
rect 3605 16711 3663 16717
rect 3605 16708 3617 16711
rect 2869 16671 2927 16677
rect 3528 16680 3617 16708
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16609 2467 16643
rect 2409 16603 2467 16609
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16609 2559 16643
rect 2501 16603 2559 16609
rect 2593 16643 2651 16649
rect 2593 16609 2605 16643
rect 2639 16640 2651 16643
rect 2682 16640 2688 16652
rect 2639 16612 2688 16640
rect 2639 16609 2651 16612
rect 2593 16603 2651 16609
rect 2516 16504 2544 16603
rect 2682 16600 2688 16612
rect 2740 16600 2746 16652
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 2958 16640 2964 16652
rect 2823 16612 2964 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3418 16600 3424 16652
rect 3476 16600 3482 16652
rect 3528 16649 3556 16680
rect 3605 16677 3617 16680
rect 3651 16708 3663 16711
rect 4525 16711 4583 16717
rect 4525 16708 4537 16711
rect 3651 16680 4537 16708
rect 3651 16677 3663 16680
rect 3605 16671 3663 16677
rect 4525 16677 4537 16680
rect 4571 16708 4583 16711
rect 4706 16708 4712 16720
rect 4571 16680 4712 16708
rect 4571 16677 4583 16680
rect 4525 16671 4583 16677
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 5368 16708 5396 16736
rect 5368 16680 5856 16708
rect 3513 16643 3571 16649
rect 3513 16609 3525 16643
rect 3559 16609 3571 16643
rect 3513 16603 3571 16609
rect 3789 16643 3847 16649
rect 3789 16609 3801 16643
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4154 16640 4160 16652
rect 4111 16612 4160 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 2774 16504 2780 16516
rect 2516 16476 2780 16504
rect 2774 16464 2780 16476
rect 2832 16464 2838 16516
rect 3436 16504 3464 16600
rect 3804 16572 3832 16603
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4798 16640 4804 16652
rect 4304 16612 4804 16640
rect 4304 16600 4310 16612
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 5169 16643 5227 16649
rect 5169 16640 5181 16643
rect 4948 16612 5181 16640
rect 4948 16600 4954 16612
rect 5169 16609 5181 16612
rect 5215 16640 5227 16643
rect 5258 16640 5264 16652
rect 5215 16612 5264 16640
rect 5215 16609 5227 16612
rect 5169 16603 5227 16609
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 5368 16649 5396 16680
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16609 5595 16643
rect 5537 16603 5595 16609
rect 3878 16572 3884 16584
rect 3804 16544 3884 16572
rect 3878 16532 3884 16544
rect 3936 16572 3942 16584
rect 5552 16572 5580 16603
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 5828 16649 5856 16680
rect 5902 16668 5908 16720
rect 5960 16708 5966 16720
rect 6362 16708 6368 16720
rect 5960 16680 6368 16708
rect 5960 16668 5966 16680
rect 6362 16668 6368 16680
rect 6420 16668 6426 16720
rect 5813 16643 5871 16649
rect 5813 16609 5825 16643
rect 5859 16609 5871 16643
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 5813 16603 5871 16609
rect 5920 16612 6193 16640
rect 5920 16572 5948 16612
rect 6181 16609 6193 16612
rect 6227 16640 6239 16643
rect 6472 16640 6500 16739
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 8941 16779 8999 16785
rect 8941 16745 8953 16779
rect 8987 16776 8999 16779
rect 9766 16776 9772 16788
rect 8987 16748 9772 16776
rect 8987 16745 8999 16748
rect 8941 16739 8999 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 10410 16736 10416 16788
rect 10468 16776 10474 16788
rect 10870 16776 10876 16788
rect 10468 16748 10876 16776
rect 10468 16736 10474 16748
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 14550 16736 14556 16788
rect 14608 16736 14614 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 18509 16779 18567 16785
rect 18509 16776 18521 16779
rect 16356 16748 18521 16776
rect 16356 16736 16362 16748
rect 18509 16745 18521 16748
rect 18555 16745 18567 16779
rect 18509 16739 18567 16745
rect 18969 16779 19027 16785
rect 18969 16745 18981 16779
rect 19015 16776 19027 16779
rect 19058 16776 19064 16788
rect 19015 16748 19064 16776
rect 19015 16745 19027 16748
rect 18969 16739 19027 16745
rect 19058 16736 19064 16748
rect 19116 16736 19122 16788
rect 19150 16736 19156 16788
rect 19208 16736 19214 16788
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 20990 16776 20996 16788
rect 19576 16748 20996 16776
rect 19576 16736 19582 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 22646 16736 22652 16788
rect 22704 16736 22710 16788
rect 24489 16779 24547 16785
rect 24489 16745 24501 16779
rect 24535 16776 24547 16779
rect 25774 16776 25780 16788
rect 24535 16748 25780 16776
rect 24535 16745 24547 16748
rect 24489 16739 24547 16745
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 28169 16779 28227 16785
rect 28169 16745 28181 16779
rect 28215 16776 28227 16779
rect 29730 16776 29736 16788
rect 28215 16748 29736 16776
rect 28215 16745 28227 16748
rect 28169 16739 28227 16745
rect 29730 16736 29736 16748
rect 29788 16736 29794 16788
rect 30098 16736 30104 16788
rect 30156 16776 30162 16788
rect 30742 16776 30748 16788
rect 30156 16748 30748 16776
rect 30156 16736 30162 16748
rect 30742 16736 30748 16748
rect 30800 16736 30806 16788
rect 6546 16668 6552 16720
rect 6604 16708 6610 16720
rect 6825 16711 6883 16717
rect 6825 16708 6837 16711
rect 6604 16680 6837 16708
rect 6604 16668 6610 16680
rect 6825 16677 6837 16680
rect 6871 16677 6883 16711
rect 6825 16671 6883 16677
rect 11333 16711 11391 16717
rect 11333 16677 11345 16711
rect 11379 16708 11391 16711
rect 11790 16708 11796 16720
rect 11379 16680 11796 16708
rect 11379 16677 11391 16680
rect 11333 16671 11391 16677
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 13633 16711 13691 16717
rect 13633 16677 13645 16711
rect 13679 16708 13691 16711
rect 13722 16708 13728 16720
rect 13679 16680 13728 16708
rect 13679 16677 13691 16680
rect 13633 16671 13691 16677
rect 13722 16668 13728 16680
rect 13780 16668 13786 16720
rect 14826 16668 14832 16720
rect 14884 16708 14890 16720
rect 15666 16711 15724 16717
rect 15666 16708 15678 16711
rect 14884 16680 15678 16708
rect 14884 16668 14890 16680
rect 15666 16677 15678 16680
rect 15712 16677 15724 16711
rect 19702 16708 19708 16720
rect 15666 16671 15724 16677
rect 17144 16680 19708 16708
rect 17144 16652 17172 16680
rect 19702 16668 19708 16680
rect 19760 16708 19766 16720
rect 19760 16680 19840 16708
rect 19760 16668 19766 16680
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 6227 16612 6500 16640
rect 6564 16612 6653 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 3936 16544 4292 16572
rect 5552 16544 5948 16572
rect 3936 16532 3942 16544
rect 3973 16507 4031 16513
rect 3973 16504 3985 16507
rect 3436 16476 3985 16504
rect 3973 16473 3985 16476
rect 4019 16473 4031 16507
rect 3973 16467 4031 16473
rect 4264 16448 4292 16544
rect 6362 16532 6368 16584
rect 6420 16532 6426 16584
rect 4893 16507 4951 16513
rect 4893 16473 4905 16507
rect 4939 16473 4951 16507
rect 4893 16467 4951 16473
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 2133 16439 2191 16445
rect 2133 16436 2145 16439
rect 2004 16408 2145 16436
rect 2004 16396 2010 16408
rect 2133 16405 2145 16408
rect 2179 16405 2191 16439
rect 2133 16399 2191 16405
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 4908 16436 4936 16467
rect 5350 16464 5356 16516
rect 5408 16504 5414 16516
rect 6564 16504 6592 16612
rect 6641 16609 6653 16612
rect 6687 16640 6699 16643
rect 6730 16640 6736 16652
rect 6687 16612 6736 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 10520 16612 10793 16640
rect 10520 16584 10548 16612
rect 10781 16609 10793 16612
rect 10827 16609 10839 16643
rect 10781 16603 10839 16609
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16640 11023 16643
rect 11054 16640 11060 16652
rect 11011 16612 11060 16640
rect 11011 16609 11023 16612
rect 10965 16603 11023 16609
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11146 16600 11152 16652
rect 11204 16600 11210 16652
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 11296 16612 11437 16640
rect 11296 16600 11302 16612
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 11606 16600 11612 16652
rect 11664 16600 11670 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 12492 16612 12725 16640
rect 12492 16600 12498 16612
rect 12713 16609 12725 16612
rect 12759 16640 12771 16643
rect 12805 16643 12863 16649
rect 12805 16640 12817 16643
rect 12759 16612 12817 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 12805 16609 12817 16612
rect 12851 16609 12863 16643
rect 12805 16603 12863 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 15979 16612 16221 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16209 16609 16221 16612
rect 16255 16609 16267 16643
rect 16209 16603 16267 16609
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16640 16359 16643
rect 17126 16640 17132 16652
rect 16347 16612 17132 16640
rect 16347 16609 16359 16612
rect 16301 16603 16359 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 17678 16600 17684 16652
rect 17736 16640 17742 16652
rect 17773 16643 17831 16649
rect 17773 16640 17785 16643
rect 17736 16612 17785 16640
rect 17736 16600 17742 16612
rect 17773 16609 17785 16612
rect 17819 16609 17831 16643
rect 17773 16603 17831 16609
rect 17862 16600 17868 16652
rect 17920 16600 17926 16652
rect 17957 16643 18015 16649
rect 17957 16609 17969 16643
rect 18003 16640 18015 16643
rect 18003 16612 18092 16640
rect 18003 16609 18015 16612
rect 17957 16603 18015 16609
rect 9766 16581 9772 16584
rect 9744 16575 9772 16581
rect 9744 16541 9756 16575
rect 9744 16535 9772 16541
rect 9766 16532 9772 16535
rect 9824 16532 9830 16584
rect 9858 16532 9864 16584
rect 9916 16532 9922 16584
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16572 10195 16575
rect 10410 16572 10416 16584
rect 10183 16544 10416 16572
rect 10183 16541 10195 16544
rect 10137 16535 10195 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10502 16532 10508 16584
rect 10560 16532 10566 16584
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 5408 16476 6592 16504
rect 10612 16504 10640 16535
rect 11974 16532 11980 16584
rect 12032 16532 12038 16584
rect 10962 16504 10968 16516
rect 10612 16476 10968 16504
rect 5408 16464 5414 16476
rect 10962 16464 10968 16476
rect 11020 16464 11026 16516
rect 11422 16464 11428 16516
rect 11480 16464 11486 16516
rect 18064 16504 18092 16612
rect 18138 16600 18144 16652
rect 18196 16600 18202 16652
rect 18248 16612 18460 16640
rect 18248 16504 18276 16612
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18432 16572 18460 16612
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 18601 16643 18659 16649
rect 18601 16640 18613 16643
rect 18564 16612 18613 16640
rect 18564 16600 18570 16612
rect 18601 16609 18613 16612
rect 18647 16609 18659 16643
rect 18601 16603 18659 16609
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19518 16640 19524 16652
rect 19024 16612 19524 16640
rect 19024 16600 19030 16612
rect 19518 16600 19524 16612
rect 19576 16640 19582 16652
rect 19613 16643 19671 16649
rect 19613 16640 19625 16643
rect 19576 16612 19625 16640
rect 19576 16600 19582 16612
rect 19613 16609 19625 16612
rect 19659 16609 19671 16643
rect 19812 16640 19840 16680
rect 19886 16668 19892 16720
rect 19944 16708 19950 16720
rect 22186 16708 22192 16720
rect 19944 16680 22192 16708
rect 19944 16668 19950 16680
rect 22186 16668 22192 16680
rect 22244 16668 22250 16720
rect 23385 16711 23443 16717
rect 23385 16677 23397 16711
rect 23431 16708 23443 16711
rect 23658 16708 23664 16720
rect 23431 16680 23664 16708
rect 23431 16677 23443 16680
rect 23385 16671 23443 16677
rect 23658 16668 23664 16680
rect 23716 16668 23722 16720
rect 24854 16668 24860 16720
rect 24912 16708 24918 16720
rect 25694 16711 25752 16717
rect 25694 16708 25706 16711
rect 24912 16680 25706 16708
rect 24912 16668 24918 16680
rect 25694 16677 25706 16680
rect 25740 16677 25752 16711
rect 30006 16708 30012 16720
rect 25694 16671 25752 16677
rect 26712 16680 30012 16708
rect 26712 16652 26740 16680
rect 30006 16668 30012 16680
rect 30064 16668 30070 16720
rect 30190 16668 30196 16720
rect 30248 16717 30254 16720
rect 30248 16708 30260 16717
rect 30248 16680 30293 16708
rect 30248 16671 30260 16680
rect 30248 16668 30254 16671
rect 20070 16640 20076 16652
rect 19812 16612 20076 16640
rect 19613 16603 19671 16609
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 20346 16600 20352 16652
rect 20404 16640 20410 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 20404 16612 21281 16640
rect 20404 16600 20410 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 21525 16643 21583 16649
rect 21525 16640 21537 16643
rect 21416 16612 21537 16640
rect 21416 16600 21422 16612
rect 21525 16609 21537 16612
rect 21571 16609 21583 16643
rect 21525 16603 21583 16609
rect 22922 16600 22928 16652
rect 22980 16600 22986 16652
rect 23014 16600 23020 16652
rect 23072 16600 23078 16652
rect 23198 16600 23204 16652
rect 23256 16600 23262 16652
rect 23293 16643 23351 16649
rect 23293 16609 23305 16643
rect 23339 16640 23351 16643
rect 23474 16640 23480 16652
rect 23339 16612 23480 16640
rect 23339 16609 23351 16612
rect 23293 16603 23351 16609
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16640 23811 16643
rect 23845 16643 23903 16649
rect 23845 16640 23857 16643
rect 23799 16612 23857 16640
rect 23799 16609 23811 16612
rect 23753 16603 23811 16609
rect 23845 16609 23857 16612
rect 23891 16609 23903 16643
rect 23845 16603 23903 16609
rect 18432 16544 20300 16572
rect 18325 16535 18383 16541
rect 18064 16476 18276 16504
rect 5994 16436 6000 16448
rect 4304 16408 6000 16436
rect 4304 16396 4310 16408
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 17494 16396 17500 16448
rect 17552 16396 17558 16448
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 18340 16436 18368 16535
rect 19058 16464 19064 16516
rect 19116 16504 19122 16516
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 19116 16476 19257 16504
rect 19116 16464 19122 16476
rect 19245 16473 19257 16476
rect 19291 16473 19303 16507
rect 19245 16467 19303 16473
rect 19426 16464 19432 16516
rect 19484 16504 19490 16516
rect 19702 16504 19708 16516
rect 19484 16476 19708 16504
rect 19484 16464 19490 16476
rect 19702 16464 19708 16476
rect 19760 16464 19766 16516
rect 20272 16448 20300 16544
rect 22462 16532 22468 16584
rect 22520 16572 22526 16584
rect 22741 16575 22799 16581
rect 22741 16572 22753 16575
rect 22520 16544 22753 16572
rect 22520 16532 22526 16544
rect 22741 16541 22753 16544
rect 22787 16541 22799 16575
rect 23584 16572 23612 16603
rect 24026 16600 24032 16652
rect 24084 16600 24090 16652
rect 24118 16600 24124 16652
rect 24176 16600 24182 16652
rect 24213 16643 24271 16649
rect 24213 16609 24225 16643
rect 24259 16640 24271 16643
rect 25222 16640 25228 16652
rect 24259 16638 24900 16640
rect 25056 16638 25228 16640
rect 24259 16612 25228 16638
rect 24259 16609 24271 16612
rect 24872 16610 25084 16612
rect 24213 16603 24271 16609
rect 25222 16600 25228 16612
rect 25280 16600 25286 16652
rect 25961 16643 26019 16649
rect 25961 16609 25973 16643
rect 26007 16640 26019 16643
rect 26145 16643 26203 16649
rect 26145 16640 26157 16643
rect 26007 16612 26157 16640
rect 26007 16609 26019 16612
rect 25961 16603 26019 16609
rect 26145 16609 26157 16612
rect 26191 16609 26203 16643
rect 26145 16603 26203 16609
rect 26237 16643 26295 16649
rect 26237 16609 26249 16643
rect 26283 16640 26295 16643
rect 26694 16640 26700 16652
rect 26283 16612 26700 16640
rect 26283 16609 26295 16612
rect 26237 16603 26295 16609
rect 26694 16600 26700 16612
rect 26752 16600 26758 16652
rect 27801 16643 27859 16649
rect 27801 16609 27813 16643
rect 27847 16640 27859 16643
rect 27890 16640 27896 16652
rect 27847 16612 27896 16640
rect 27847 16609 27859 16612
rect 27801 16603 27859 16609
rect 22741 16535 22799 16541
rect 23400 16544 23612 16572
rect 24136 16572 24164 16600
rect 27816 16572 27844 16603
rect 27890 16600 27896 16612
rect 27948 16600 27954 16652
rect 27985 16643 28043 16649
rect 27985 16609 27997 16643
rect 28031 16640 28043 16643
rect 28031 16612 28580 16640
rect 28031 16609 28043 16612
rect 27985 16603 28043 16609
rect 28442 16572 28448 16584
rect 24136 16544 24900 16572
rect 23400 16516 23428 16544
rect 22554 16464 22560 16516
rect 22612 16504 22618 16516
rect 22612 16476 23336 16504
rect 22612 16464 22618 16476
rect 17736 16408 18368 16436
rect 17736 16396 17742 16408
rect 20254 16396 20260 16448
rect 20312 16396 20318 16448
rect 23308 16436 23336 16476
rect 23382 16464 23388 16516
rect 23440 16464 23446 16516
rect 24486 16504 24492 16516
rect 23860 16476 24492 16504
rect 23860 16436 23888 16476
rect 24486 16464 24492 16476
rect 24544 16464 24550 16516
rect 24581 16507 24639 16513
rect 24581 16473 24593 16507
rect 24627 16504 24639 16507
rect 24762 16504 24768 16516
rect 24627 16476 24768 16504
rect 24627 16473 24639 16476
rect 24581 16467 24639 16473
rect 24762 16464 24768 16476
rect 24820 16464 24826 16516
rect 23308 16408 23888 16436
rect 24872 16436 24900 16544
rect 27356 16544 28448 16572
rect 27356 16516 27384 16544
rect 28442 16532 28448 16544
rect 28500 16532 28506 16584
rect 28552 16572 28580 16612
rect 28626 16600 28632 16652
rect 28684 16600 28690 16652
rect 28718 16600 28724 16652
rect 28776 16600 28782 16652
rect 28810 16600 28816 16652
rect 28868 16600 28874 16652
rect 28902 16600 28908 16652
rect 28960 16640 28966 16652
rect 28997 16643 29055 16649
rect 28997 16640 29009 16643
rect 28960 16612 29009 16640
rect 28960 16600 28966 16612
rect 28997 16609 29009 16612
rect 29043 16609 29055 16643
rect 28997 16603 29055 16609
rect 30469 16643 30527 16649
rect 30469 16609 30481 16643
rect 30515 16640 30527 16643
rect 31202 16640 31208 16652
rect 30515 16612 31208 16640
rect 30515 16609 30527 16612
rect 30469 16603 30527 16609
rect 31202 16600 31208 16612
rect 31260 16600 31266 16652
rect 28552 16544 29132 16572
rect 27338 16464 27344 16516
rect 27396 16464 27402 16516
rect 27614 16464 27620 16516
rect 27672 16504 27678 16516
rect 28353 16507 28411 16513
rect 28353 16504 28365 16507
rect 27672 16476 28365 16504
rect 27672 16464 27678 16476
rect 28353 16473 28365 16476
rect 28399 16473 28411 16507
rect 28353 16467 28411 16473
rect 25958 16436 25964 16448
rect 24872 16408 25964 16436
rect 25958 16396 25964 16408
rect 26016 16396 26022 16448
rect 27522 16396 27528 16448
rect 27580 16436 27586 16448
rect 28994 16436 29000 16448
rect 27580 16408 29000 16436
rect 27580 16396 27586 16408
rect 28994 16396 29000 16408
rect 29052 16396 29058 16448
rect 29104 16445 29132 16544
rect 29089 16439 29147 16445
rect 29089 16405 29101 16439
rect 29135 16436 29147 16439
rect 30282 16436 30288 16448
rect 29135 16408 30288 16436
rect 29135 16405 29147 16408
rect 29089 16399 29147 16405
rect 30282 16396 30288 16408
rect 30340 16396 30346 16448
rect 552 16346 31648 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 11436 16346
rect 11488 16294 11500 16346
rect 11552 16294 11564 16346
rect 11616 16294 11628 16346
rect 11680 16294 11692 16346
rect 11744 16294 19210 16346
rect 19262 16294 19274 16346
rect 19326 16294 19338 16346
rect 19390 16294 19402 16346
rect 19454 16294 19466 16346
rect 19518 16294 26984 16346
rect 27036 16294 27048 16346
rect 27100 16294 27112 16346
rect 27164 16294 27176 16346
rect 27228 16294 27240 16346
rect 27292 16294 31648 16346
rect 552 16272 31648 16294
rect 4890 16192 4896 16244
rect 4948 16232 4954 16244
rect 4985 16235 5043 16241
rect 4985 16232 4997 16235
rect 4948 16204 4997 16232
rect 4948 16192 4954 16204
rect 4985 16201 4997 16204
rect 5031 16201 5043 16235
rect 4985 16195 5043 16201
rect 2682 16124 2688 16176
rect 2740 16164 2746 16176
rect 3053 16167 3111 16173
rect 3053 16164 3065 16167
rect 2740 16136 3065 16164
rect 2740 16124 2746 16136
rect 3053 16133 3065 16136
rect 3099 16164 3111 16167
rect 4617 16167 4675 16173
rect 4617 16164 4629 16167
rect 3099 16136 4629 16164
rect 3099 16133 3111 16136
rect 3053 16127 3111 16133
rect 4617 16133 4629 16136
rect 4663 16164 4675 16167
rect 4706 16164 4712 16176
rect 4663 16136 4712 16164
rect 4663 16133 4675 16136
rect 4617 16127 4675 16133
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 5000 16164 5028 16195
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 5537 16235 5595 16241
rect 5537 16232 5549 16235
rect 5224 16204 5549 16232
rect 5224 16192 5230 16204
rect 5537 16201 5549 16204
rect 5583 16201 5595 16235
rect 5537 16195 5595 16201
rect 8941 16235 8999 16241
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 9490 16232 9496 16244
rect 8987 16204 9496 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17276 16204 17509 16232
rect 17276 16192 17282 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 18414 16192 18420 16244
rect 18472 16192 18478 16244
rect 19058 16192 19064 16244
rect 19116 16192 19122 16244
rect 19518 16192 19524 16244
rect 19576 16232 19582 16244
rect 20162 16232 20168 16244
rect 19576 16204 20168 16232
rect 19576 16192 19582 16204
rect 20162 16192 20168 16204
rect 20220 16232 20226 16244
rect 20622 16232 20628 16244
rect 20220 16204 20628 16232
rect 20220 16192 20226 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 22278 16232 22284 16244
rect 21192 16204 22284 16232
rect 5810 16164 5816 16176
rect 5000 16136 5816 16164
rect 5810 16124 5816 16136
rect 5868 16124 5874 16176
rect 8570 16124 8576 16176
rect 8628 16164 8634 16176
rect 11054 16164 11060 16176
rect 8628 16136 11060 16164
rect 8628 16124 8634 16136
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 17678 16124 17684 16176
rect 17736 16164 17742 16176
rect 20346 16164 20352 16176
rect 17736 16136 20352 16164
rect 17736 16124 17742 16136
rect 4246 16056 4252 16108
rect 4304 16056 4310 16108
rect 1394 15988 1400 16040
rect 1452 15988 1458 16040
rect 1946 16037 1952 16040
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1673 16031 1731 16037
rect 1673 16028 1685 16031
rect 1535 16000 1685 16028
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 1673 15997 1685 16000
rect 1719 15997 1731 16031
rect 1940 16028 1952 16037
rect 1907 16000 1952 16028
rect 1673 15991 1731 15997
rect 1940 15991 1952 16000
rect 1946 15988 1952 15991
rect 2004 15988 2010 16040
rect 4154 15988 4160 16040
rect 4212 16028 4218 16040
rect 5350 16028 5356 16040
rect 4212 16000 5356 16028
rect 4212 15988 4218 16000
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5626 15988 5632 16040
rect 5684 15988 5690 16040
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 6604 16000 6745 16028
rect 6604 15988 6610 16000
rect 6733 15997 6745 16000
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 8018 15988 8024 16040
rect 8076 15988 8082 16040
rect 8588 16037 8616 16124
rect 9950 16096 9956 16108
rect 9416 16068 9956 16096
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 9306 15988 9312 16040
rect 9364 15988 9370 16040
rect 9416 16037 9444 16068
rect 9950 16056 9956 16068
rect 10008 16096 10014 16108
rect 10226 16096 10232 16108
rect 10008 16068 10232 16096
rect 10008 16056 10014 16068
rect 10226 16056 10232 16068
rect 10284 16096 10290 16108
rect 10284 16068 13952 16096
rect 10284 16056 10290 16068
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9490 15988 9496 16040
rect 9548 15988 9554 16040
rect 9674 15988 9680 16040
rect 9732 15988 9738 16040
rect 9766 15988 9772 16040
rect 9824 16028 9830 16040
rect 10597 16031 10655 16037
rect 10597 16028 10609 16031
rect 9824 16000 10609 16028
rect 9824 15988 9830 16000
rect 10597 15997 10609 16000
rect 10643 15997 10655 16031
rect 10597 15991 10655 15997
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 11020 16000 11069 16028
rect 11020 15988 11026 16000
rect 11057 15997 11069 16000
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 11974 15988 11980 16040
rect 12032 16028 12038 16040
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 12032 16000 13001 16028
rect 12032 15988 12038 16000
rect 12989 15997 13001 16000
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 4985 15963 5043 15969
rect 4985 15960 4997 15963
rect 4724 15932 4997 15960
rect 4724 15901 4752 15932
rect 4985 15929 4997 15932
rect 5031 15960 5043 15963
rect 5534 15960 5540 15972
rect 5031 15932 5540 15960
rect 5031 15929 5043 15932
rect 4985 15923 5043 15929
rect 5534 15920 5540 15932
rect 5592 15920 5598 15972
rect 5718 15920 5724 15972
rect 5776 15960 5782 15972
rect 5813 15963 5871 15969
rect 5813 15960 5825 15963
rect 5776 15932 5825 15960
rect 5776 15920 5782 15932
rect 5813 15929 5825 15932
rect 5859 15929 5871 15963
rect 5813 15923 5871 15929
rect 6638 15920 6644 15972
rect 6696 15920 6702 15972
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15960 8815 15963
rect 10045 15963 10103 15969
rect 10045 15960 10057 15963
rect 8803 15932 10057 15960
rect 8803 15929 8815 15932
rect 8757 15923 8815 15929
rect 10045 15929 10057 15932
rect 10091 15929 10103 15963
rect 13004 15960 13032 15991
rect 13262 15988 13268 16040
rect 13320 16028 13326 16040
rect 13924 16037 13952 16068
rect 19518 16056 19524 16108
rect 19576 16056 19582 16108
rect 19628 16105 19656 16136
rect 20346 16124 20352 16136
rect 20404 16164 20410 16176
rect 21082 16164 21088 16176
rect 20404 16136 21088 16164
rect 20404 16124 20410 16136
rect 21082 16124 21088 16136
rect 21140 16124 21146 16176
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19702 16056 19708 16108
rect 19760 16056 19766 16108
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 20993 16099 21051 16105
rect 20993 16096 21005 16099
rect 20772 16068 21005 16096
rect 20772 16056 20778 16068
rect 20993 16065 21005 16068
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13320 16000 13829 16028
rect 13320 15988 13326 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 13998 15988 14004 16040
rect 14056 15988 14062 16040
rect 14182 15988 14188 16040
rect 14240 15988 14246 16040
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 17586 15988 17592 16040
rect 17644 16037 17650 16040
rect 17644 16031 17693 16037
rect 17644 15997 17647 16031
rect 17681 15997 17693 16031
rect 17644 15991 17693 15997
rect 17644 15988 17650 15991
rect 17770 15988 17776 16040
rect 17828 15988 17834 16040
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 17920 16000 18337 16028
rect 17920 15988 17926 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 19429 16031 19487 16037
rect 19429 15997 19441 16031
rect 19475 16028 19487 16031
rect 19720 16028 19748 16056
rect 19475 16000 19748 16028
rect 19475 15997 19487 16000
rect 19429 15991 19487 15997
rect 19886 15988 19892 16040
rect 19944 15988 19950 16040
rect 21100 16028 21128 16124
rect 21192 16105 21220 16204
rect 22278 16192 22284 16204
rect 22336 16232 22342 16244
rect 23382 16232 23388 16244
rect 22336 16204 23388 16232
rect 22336 16192 22342 16204
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 25317 16235 25375 16241
rect 25317 16232 25329 16235
rect 25188 16204 25329 16232
rect 25188 16192 25194 16204
rect 25317 16201 25329 16204
rect 25363 16201 25375 16235
rect 25317 16195 25375 16201
rect 25498 16192 25504 16244
rect 25556 16232 25562 16244
rect 27065 16235 27123 16241
rect 27065 16232 27077 16235
rect 25556 16204 27077 16232
rect 25556 16192 25562 16204
rect 27065 16201 27077 16204
rect 27111 16201 27123 16235
rect 27065 16195 27123 16201
rect 28077 16235 28135 16241
rect 28077 16201 28089 16235
rect 28123 16232 28135 16235
rect 29178 16232 29184 16244
rect 28123 16204 29184 16232
rect 28123 16201 28135 16204
rect 28077 16195 28135 16201
rect 29178 16192 29184 16204
rect 29236 16192 29242 16244
rect 21637 16167 21695 16173
rect 21637 16133 21649 16167
rect 21683 16133 21695 16167
rect 21637 16127 21695 16133
rect 21177 16099 21235 16105
rect 21177 16065 21189 16099
rect 21223 16065 21235 16099
rect 21177 16059 21235 16065
rect 21269 16031 21327 16037
rect 21269 16028 21281 16031
rect 21100 16000 21281 16028
rect 21269 15997 21281 16000
rect 21315 15997 21327 16031
rect 21652 16028 21680 16127
rect 21818 16124 21824 16176
rect 21876 16164 21882 16176
rect 22557 16167 22615 16173
rect 22557 16164 22569 16167
rect 21876 16136 22569 16164
rect 21876 16124 21882 16136
rect 22557 16133 22569 16136
rect 22603 16164 22615 16167
rect 24118 16164 24124 16176
rect 22603 16136 24124 16164
rect 22603 16133 22615 16136
rect 22557 16127 22615 16133
rect 24118 16124 24124 16136
rect 24176 16124 24182 16176
rect 26142 16164 26148 16176
rect 24688 16136 26148 16164
rect 24688 16105 24716 16136
rect 26142 16124 26148 16136
rect 26200 16124 26206 16176
rect 28997 16167 29055 16173
rect 28997 16164 29009 16167
rect 28092 16136 29009 16164
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16065 24731 16099
rect 25222 16096 25228 16108
rect 24673 16059 24731 16065
rect 24872 16068 25228 16096
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21652 16000 21925 16028
rect 21269 15991 21327 15997
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 22002 15988 22008 16040
rect 22060 15988 22066 16040
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 22189 16031 22247 16037
rect 22189 16028 22201 16031
rect 22152 16000 22201 16028
rect 22152 15988 22158 16000
rect 22189 15997 22201 16000
rect 22235 15997 22247 16031
rect 22189 15991 22247 15997
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 22373 16031 22431 16037
rect 22373 15997 22385 16031
rect 22419 16028 22431 16031
rect 22554 16028 22560 16040
rect 22419 16000 22560 16028
rect 22419 15997 22431 16000
rect 22373 15991 22431 15997
rect 14918 15960 14924 15972
rect 13004 15932 14924 15960
rect 10045 15923 10103 15929
rect 14918 15920 14924 15932
rect 14976 15920 14982 15972
rect 18049 15963 18107 15969
rect 18049 15929 18061 15963
rect 18095 15929 18107 15963
rect 18049 15923 18107 15929
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15861 4767 15895
rect 4709 15855 4767 15861
rect 4798 15852 4804 15904
rect 4856 15852 4862 15904
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 7340 15864 7389 15892
rect 7340 15852 7346 15864
rect 7377 15861 7389 15864
rect 7423 15861 7435 15895
rect 7377 15855 7435 15861
rect 8110 15852 8116 15904
rect 8168 15852 8174 15904
rect 9030 15852 9036 15904
rect 9088 15852 9094 15904
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 10318 15892 10324 15904
rect 9364 15864 10324 15892
rect 9364 15852 9370 15864
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 11701 15895 11759 15901
rect 11701 15861 11713 15895
rect 11747 15892 11759 15895
rect 11882 15892 11888 15904
rect 11747 15864 11888 15892
rect 11747 15861 11759 15864
rect 11701 15855 11759 15861
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 13078 15852 13084 15904
rect 13136 15852 13142 15904
rect 13538 15852 13544 15904
rect 13596 15852 13602 15904
rect 17218 15852 17224 15904
rect 17276 15852 17282 15904
rect 17770 15852 17776 15904
rect 17828 15892 17834 15904
rect 18064 15892 18092 15923
rect 18138 15920 18144 15972
rect 18196 15920 18202 15972
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 20128 15932 20729 15960
rect 20128 15920 20134 15932
rect 20717 15929 20729 15932
rect 20763 15960 20775 15963
rect 22296 15960 22324 15991
rect 22554 15988 22560 16000
rect 22612 15988 22618 16040
rect 22646 15988 22652 16040
rect 22704 16028 22710 16040
rect 22741 16031 22799 16037
rect 22741 16028 22753 16031
rect 22704 16000 22753 16028
rect 22704 15988 22710 16000
rect 22741 15997 22753 16000
rect 22787 15997 22799 16031
rect 22741 15991 22799 15997
rect 23658 15988 23664 16040
rect 23716 16028 23722 16040
rect 24029 16031 24087 16037
rect 24029 16028 24041 16031
rect 23716 16000 24041 16028
rect 23716 15988 23722 16000
rect 24029 15997 24041 16000
rect 24075 15997 24087 16031
rect 24029 15991 24087 15997
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 16028 24271 16031
rect 24762 16028 24768 16040
rect 24259 16000 24768 16028
rect 24259 15997 24271 16000
rect 24213 15991 24271 15997
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 24872 16037 24900 16068
rect 25222 16056 25228 16068
rect 25280 16096 25286 16108
rect 25280 16068 26188 16096
rect 25280 16056 25286 16068
rect 24857 16031 24915 16037
rect 24857 15997 24869 16031
rect 24903 15997 24915 16031
rect 25501 16031 25559 16037
rect 25501 16028 25513 16031
rect 24857 15991 24915 15997
rect 25240 16000 25513 16028
rect 22462 15960 22468 15972
rect 20763 15932 21864 15960
rect 22296 15932 22468 15960
rect 20763 15929 20775 15932
rect 20717 15923 20775 15929
rect 17828 15864 18092 15892
rect 17828 15852 17834 15864
rect 18414 15852 18420 15904
rect 18472 15892 18478 15904
rect 18690 15892 18696 15904
rect 18472 15864 18696 15892
rect 18472 15852 18478 15864
rect 18690 15852 18696 15864
rect 18748 15892 18754 15904
rect 21266 15892 21272 15904
rect 18748 15864 21272 15892
rect 18748 15852 18754 15864
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 21726 15852 21732 15904
rect 21784 15852 21790 15904
rect 21836 15892 21864 15932
rect 22462 15920 22468 15932
rect 22520 15960 22526 15972
rect 23474 15960 23480 15972
rect 22520 15932 23480 15960
rect 22520 15920 22526 15932
rect 23474 15920 23480 15932
rect 23532 15920 23538 15972
rect 24397 15963 24455 15969
rect 24397 15929 24409 15963
rect 24443 15960 24455 15963
rect 24946 15960 24952 15972
rect 24443 15932 24952 15960
rect 24443 15929 24455 15932
rect 24397 15923 24455 15929
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 22370 15892 22376 15904
rect 21836 15864 22376 15892
rect 22370 15852 22376 15864
rect 22428 15852 22434 15904
rect 22922 15852 22928 15904
rect 22980 15852 22986 15904
rect 23382 15852 23388 15904
rect 23440 15892 23446 15904
rect 25240 15901 25268 16000
rect 25501 15997 25513 16000
rect 25547 15997 25559 16031
rect 25501 15991 25559 15997
rect 25593 16031 25651 16037
rect 25593 15997 25605 16031
rect 25639 15997 25651 16031
rect 25593 15991 25651 15997
rect 25406 15920 25412 15972
rect 25464 15960 25470 15972
rect 25608 15960 25636 15991
rect 25774 15988 25780 16040
rect 25832 15988 25838 16040
rect 25869 16031 25927 16037
rect 25869 15997 25881 16031
rect 25915 15997 25927 16031
rect 25869 15991 25927 15997
rect 25464 15932 25636 15960
rect 25884 15960 25912 15991
rect 26050 15988 26056 16040
rect 26108 15988 26114 16040
rect 26160 16028 26188 16068
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 26160 16000 27261 16028
rect 27249 15997 27261 16000
rect 27295 15997 27307 16031
rect 27249 15991 27307 15997
rect 27525 16031 27583 16037
rect 27525 15997 27537 16031
rect 27571 15997 27583 16031
rect 27525 15991 27583 15997
rect 25884 15932 26280 15960
rect 25464 15920 25470 15932
rect 26252 15904 26280 15932
rect 26694 15920 26700 15972
rect 26752 15960 26758 15972
rect 26789 15963 26847 15969
rect 26789 15960 26801 15963
rect 26752 15932 26801 15960
rect 26752 15920 26758 15932
rect 26789 15929 26801 15932
rect 26835 15929 26847 15963
rect 26789 15923 26847 15929
rect 27338 15920 27344 15972
rect 27396 15960 27402 15972
rect 27433 15963 27491 15969
rect 27433 15960 27445 15963
rect 27396 15932 27445 15960
rect 27396 15920 27402 15932
rect 27433 15929 27445 15932
rect 27479 15929 27491 15963
rect 27433 15923 27491 15929
rect 24765 15895 24823 15901
rect 24765 15892 24777 15895
rect 23440 15864 24777 15892
rect 23440 15852 23446 15864
rect 24765 15861 24777 15864
rect 24811 15861 24823 15895
rect 24765 15855 24823 15861
rect 25225 15895 25283 15901
rect 25225 15861 25237 15895
rect 25271 15861 25283 15895
rect 25225 15855 25283 15861
rect 26234 15852 26240 15904
rect 26292 15892 26298 15904
rect 27540 15892 27568 15991
rect 27614 15988 27620 16040
rect 27672 15988 27678 16040
rect 27798 15988 27804 16040
rect 27856 15988 27862 16040
rect 27893 16031 27951 16037
rect 27893 15997 27905 16031
rect 27939 16028 27951 16031
rect 28092 16028 28120 16136
rect 28997 16133 29009 16136
rect 29043 16133 29055 16167
rect 28997 16127 29055 16133
rect 28166 16056 28172 16108
rect 28224 16096 28230 16108
rect 29457 16099 29515 16105
rect 29457 16096 29469 16099
rect 28224 16068 29469 16096
rect 28224 16056 28230 16068
rect 29457 16065 29469 16068
rect 29503 16065 29515 16099
rect 29457 16059 29515 16065
rect 29546 16056 29552 16108
rect 29604 16056 29610 16108
rect 27939 16000 28120 16028
rect 27939 15997 27951 16000
rect 27893 15991 27951 15997
rect 28626 15988 28632 16040
rect 28684 16028 28690 16040
rect 28813 16031 28871 16037
rect 28813 16028 28825 16031
rect 28684 16000 28825 16028
rect 28684 15988 28690 16000
rect 28813 15997 28825 16000
rect 28859 16028 28871 16031
rect 28859 16000 28948 16028
rect 28859 15997 28871 16000
rect 28813 15991 28871 15997
rect 27816 15960 27844 15988
rect 28534 15960 28540 15972
rect 27816 15932 28540 15960
rect 28534 15920 28540 15932
rect 28592 15920 28598 15972
rect 28920 15904 28948 16000
rect 30006 15988 30012 16040
rect 30064 15988 30070 16040
rect 28074 15892 28080 15904
rect 26292 15864 28080 15892
rect 26292 15852 26298 15864
rect 28074 15852 28080 15864
rect 28132 15852 28138 15904
rect 28166 15852 28172 15904
rect 28224 15852 28230 15904
rect 28902 15852 28908 15904
rect 28960 15892 28966 15904
rect 29365 15895 29423 15901
rect 29365 15892 29377 15895
rect 28960 15864 29377 15892
rect 28960 15852 28966 15864
rect 29365 15861 29377 15864
rect 29411 15861 29423 15895
rect 29365 15855 29423 15861
rect 29822 15852 29828 15904
rect 29880 15892 29886 15904
rect 29917 15895 29975 15901
rect 29917 15892 29929 15895
rect 29880 15864 29929 15892
rect 29880 15852 29886 15864
rect 29917 15861 29929 15864
rect 29963 15861 29975 15895
rect 29917 15855 29975 15861
rect 552 15802 31648 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 12096 15802
rect 12148 15750 12160 15802
rect 12212 15750 12224 15802
rect 12276 15750 12288 15802
rect 12340 15750 12352 15802
rect 12404 15750 19870 15802
rect 19922 15750 19934 15802
rect 19986 15750 19998 15802
rect 20050 15750 20062 15802
rect 20114 15750 20126 15802
rect 20178 15750 27644 15802
rect 27696 15750 27708 15802
rect 27760 15750 27772 15802
rect 27824 15750 27836 15802
rect 27888 15750 27900 15802
rect 27952 15750 31648 15802
rect 552 15728 31648 15750
rect 2682 15648 2688 15700
rect 2740 15648 2746 15700
rect 5994 15648 6000 15700
rect 6052 15688 6058 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 6052 15660 7205 15688
rect 6052 15648 6058 15660
rect 7193 15657 7205 15660
rect 7239 15657 7251 15691
rect 7193 15651 7251 15657
rect 7282 15648 7288 15700
rect 7340 15648 7346 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 9824 15660 10149 15688
rect 9824 15648 9830 15660
rect 10137 15657 10149 15660
rect 10183 15688 10195 15691
rect 10410 15688 10416 15700
rect 10183 15660 10416 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 10888 15660 11100 15688
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 5534 15620 5540 15632
rect 1452 15592 5540 15620
rect 1452 15580 1458 15592
rect 1302 15512 1308 15564
rect 1360 15512 1366 15564
rect 4448 15561 4476 15592
rect 5534 15580 5540 15592
rect 5592 15620 5598 15632
rect 5718 15620 5724 15632
rect 5592 15592 5724 15620
rect 5592 15580 5598 15592
rect 5718 15580 5724 15592
rect 5776 15580 5782 15632
rect 5813 15623 5871 15629
rect 5813 15589 5825 15623
rect 5859 15620 5871 15623
rect 6638 15620 6644 15632
rect 5859 15592 6644 15620
rect 5859 15589 5871 15592
rect 5813 15583 5871 15589
rect 6638 15580 6644 15592
rect 6696 15620 6702 15632
rect 10888 15620 10916 15660
rect 6696 15592 10916 15620
rect 11072 15620 11100 15660
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11204 15660 11621 15688
rect 11204 15648 11210 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 12161 15691 12219 15697
rect 12161 15657 12173 15691
rect 12207 15688 12219 15691
rect 13998 15688 14004 15700
rect 12207 15660 14004 15688
rect 12207 15657 12219 15660
rect 12161 15651 12219 15657
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 14182 15648 14188 15700
rect 14240 15648 14246 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 18601 15691 18659 15697
rect 18601 15688 18613 15691
rect 17828 15660 18613 15688
rect 17828 15648 17834 15660
rect 18601 15657 18613 15660
rect 18647 15657 18659 15691
rect 18969 15691 19027 15697
rect 18969 15688 18981 15691
rect 18601 15651 18659 15657
rect 18708 15660 18981 15688
rect 12434 15620 12440 15632
rect 11072 15592 12440 15620
rect 6696 15580 6702 15592
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 13078 15580 13084 15632
rect 13136 15620 13142 15632
rect 14200 15620 14228 15648
rect 13136 15592 13676 15620
rect 13136 15580 13142 15592
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 3145 15555 3203 15561
rect 3145 15552 3157 15555
rect 2823 15524 3157 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3145 15521 3157 15524
rect 3191 15521 3203 15555
rect 3145 15515 3203 15521
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 5500 15524 6561 15552
rect 5500 15512 5506 15524
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 9030 15561 9036 15564
rect 8757 15555 8815 15561
rect 8757 15552 8769 15555
rect 8168 15524 8769 15552
rect 8168 15512 8174 15524
rect 8757 15521 8769 15524
rect 8803 15521 8815 15555
rect 9024 15552 9036 15561
rect 8991 15524 9036 15552
rect 8757 15515 8815 15521
rect 9024 15515 9036 15524
rect 9030 15512 9036 15515
rect 9088 15512 9094 15564
rect 9858 15512 9864 15564
rect 9916 15552 9922 15564
rect 10413 15555 10471 15561
rect 10413 15552 10425 15555
rect 9916 15524 10425 15552
rect 9916 15512 9922 15524
rect 10413 15521 10425 15524
rect 10459 15552 10471 15555
rect 10689 15555 10747 15561
rect 10459 15524 10640 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15453 2283 15487
rect 2225 15447 2283 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3050 15484 3056 15496
rect 3007 15456 3056 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 2240 15416 2268 15447
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 3789 15487 3847 15493
rect 3789 15453 3801 15487
rect 3835 15484 3847 15487
rect 4062 15484 4068 15496
rect 3835 15456 4068 15484
rect 3835 15453 3847 15456
rect 3789 15447 3847 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 7156 15456 7389 15484
rect 7156 15444 7162 15456
rect 7377 15453 7389 15456
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 10612 15484 10640 15524
rect 10689 15521 10701 15555
rect 10735 15552 10747 15555
rect 10870 15552 10876 15564
rect 10735 15524 10876 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11793 15555 11851 15561
rect 11793 15552 11805 15555
rect 11112 15524 11805 15552
rect 11112 15512 11118 15524
rect 11793 15521 11805 15524
rect 11839 15521 11851 15555
rect 11793 15515 11851 15521
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10612 15456 10977 15484
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 11808 15484 11836 15515
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 11977 15555 12035 15561
rect 11977 15552 11989 15555
rect 11940 15524 11989 15552
rect 11940 15512 11946 15524
rect 11977 15521 11989 15524
rect 12023 15521 12035 15555
rect 11977 15515 12035 15521
rect 13377 15555 13435 15561
rect 13377 15521 13389 15555
rect 13423 15552 13435 15555
rect 13538 15552 13544 15564
rect 13423 15524 13544 15552
rect 13423 15521 13435 15524
rect 13377 15515 13435 15521
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 13648 15561 13676 15592
rect 13832 15592 14228 15620
rect 13832 15564 13860 15592
rect 15562 15580 15568 15632
rect 15620 15620 15626 15632
rect 17494 15629 17500 15632
rect 16485 15623 16543 15629
rect 16485 15620 16497 15623
rect 15620 15592 16497 15620
rect 15620 15580 15626 15592
rect 16485 15589 16497 15592
rect 16531 15589 16543 15623
rect 17488 15620 17500 15629
rect 16485 15583 16543 15589
rect 16868 15592 17356 15620
rect 17455 15592 17500 15620
rect 13633 15555 13691 15561
rect 13633 15521 13645 15555
rect 13679 15521 13691 15555
rect 13633 15515 13691 15521
rect 13814 15512 13820 15564
rect 13872 15512 13878 15564
rect 13998 15512 14004 15564
rect 14056 15512 14062 15564
rect 14090 15512 14096 15564
rect 14148 15512 14154 15564
rect 14185 15555 14243 15561
rect 14185 15521 14197 15555
rect 14231 15521 14243 15555
rect 14185 15515 14243 15521
rect 12526 15484 12532 15496
rect 11808 15456 12532 15484
rect 10965 15447 11023 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13722 15444 13728 15496
rect 13780 15484 13786 15496
rect 14200 15484 14228 15515
rect 14826 15512 14832 15564
rect 14884 15512 14890 15564
rect 14918 15512 14924 15564
rect 14976 15512 14982 15564
rect 16758 15552 16764 15564
rect 16719 15524 16764 15552
rect 16758 15512 16764 15524
rect 16816 15512 16822 15564
rect 16868 15561 16896 15592
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15521 16911 15555
rect 16853 15515 16911 15521
rect 16945 15555 17003 15561
rect 16945 15521 16957 15555
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 15746 15484 15752 15496
rect 13780 15456 15752 15484
rect 13780 15444 13786 15456
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 2317 15419 2375 15425
rect 2317 15416 2329 15419
rect 2240 15388 2329 15416
rect 2317 15385 2329 15388
rect 2363 15385 2375 15419
rect 2317 15379 2375 15385
rect 10229 15419 10287 15425
rect 10229 15385 10241 15419
rect 10275 15416 10287 15419
rect 11238 15416 11244 15428
rect 10275 15388 11244 15416
rect 10275 15385 10287 15388
rect 10229 15379 10287 15385
rect 11238 15376 11244 15388
rect 11296 15376 11302 15428
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 15013 15419 15071 15425
rect 15013 15416 15025 15419
rect 14148 15388 15025 15416
rect 14148 15376 14154 15388
rect 15013 15385 15025 15388
rect 15059 15385 15071 15419
rect 15013 15379 15071 15385
rect 1394 15308 1400 15360
rect 1452 15308 1458 15360
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 6822 15308 6828 15360
rect 6880 15308 6886 15360
rect 10410 15308 10416 15360
rect 10468 15308 10474 15360
rect 10962 15308 10968 15360
rect 11020 15348 11026 15360
rect 12253 15351 12311 15357
rect 12253 15348 12265 15351
rect 11020 15320 12265 15348
rect 11020 15308 11026 15320
rect 12253 15317 12265 15320
rect 12299 15317 12311 15351
rect 12253 15311 12311 15317
rect 14366 15308 14372 15360
rect 14424 15348 14430 15360
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 14424 15320 14473 15348
rect 14424 15308 14430 15320
rect 14461 15317 14473 15320
rect 14507 15317 14519 15351
rect 14461 15311 14519 15317
rect 14642 15308 14648 15360
rect 14700 15308 14706 15360
rect 16960 15348 16988 15515
rect 17034 15512 17040 15564
rect 17092 15552 17098 15564
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 17092 15524 17141 15552
rect 17092 15512 17098 15524
rect 17129 15521 17141 15524
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 17328 15552 17356 15592
rect 17488 15583 17500 15592
rect 17494 15580 17500 15583
rect 17552 15580 17558 15632
rect 18322 15580 18328 15632
rect 18380 15620 18386 15632
rect 18506 15620 18512 15632
rect 18380 15592 18512 15620
rect 18380 15580 18386 15592
rect 18506 15580 18512 15592
rect 18564 15620 18570 15632
rect 18708 15620 18736 15660
rect 18969 15657 18981 15660
rect 19015 15657 19027 15691
rect 18969 15651 19027 15657
rect 19061 15691 19119 15697
rect 19061 15657 19073 15691
rect 19107 15688 19119 15691
rect 20714 15688 20720 15700
rect 19107 15660 20720 15688
rect 19107 15657 19119 15660
rect 19061 15651 19119 15657
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 21358 15688 21364 15700
rect 21131 15660 21364 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 21726 15688 21732 15700
rect 21468 15660 21732 15688
rect 18564 15592 18736 15620
rect 18564 15580 18570 15592
rect 18782 15580 18788 15632
rect 18840 15620 18846 15632
rect 19429 15623 19487 15629
rect 19429 15620 19441 15623
rect 18840 15592 19441 15620
rect 18840 15580 18846 15592
rect 19429 15589 19441 15592
rect 19475 15589 19487 15623
rect 19429 15583 19487 15589
rect 19610 15580 19616 15632
rect 19668 15620 19674 15632
rect 19797 15623 19855 15629
rect 19797 15620 19809 15623
rect 19668 15592 19809 15620
rect 19668 15580 19674 15592
rect 19797 15589 19809 15592
rect 19843 15589 19855 15623
rect 19797 15583 19855 15589
rect 20165 15623 20223 15629
rect 20165 15589 20177 15623
rect 20211 15620 20223 15623
rect 20254 15620 20260 15632
rect 20211 15592 20260 15620
rect 20211 15589 20223 15592
rect 20165 15583 20223 15589
rect 20254 15580 20260 15592
rect 20312 15580 20318 15632
rect 21468 15620 21496 15660
rect 21726 15648 21732 15660
rect 21784 15648 21790 15700
rect 21913 15691 21971 15697
rect 21913 15657 21925 15691
rect 21959 15688 21971 15691
rect 22094 15688 22100 15700
rect 21959 15660 22100 15688
rect 21959 15657 21971 15660
rect 21913 15651 21971 15657
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22189 15691 22247 15697
rect 22189 15657 22201 15691
rect 22235 15688 22247 15691
rect 22462 15688 22468 15700
rect 22235 15660 22468 15688
rect 22235 15657 22247 15660
rect 22189 15651 22247 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 24302 15648 24308 15700
rect 24360 15688 24366 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 24360 15660 24501 15688
rect 24360 15648 24366 15660
rect 24489 15657 24501 15660
rect 24535 15688 24547 15691
rect 28445 15691 28503 15697
rect 24535 15660 28304 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 22278 15620 22284 15632
rect 20640 15592 21496 15620
rect 21652 15592 22284 15620
rect 18046 15552 18052 15564
rect 17328 15524 18052 15552
rect 18046 15512 18052 15524
rect 18104 15512 18110 15564
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 18877 15555 18935 15561
rect 18877 15552 18889 15555
rect 18288 15524 18889 15552
rect 18288 15512 18294 15524
rect 18877 15521 18889 15524
rect 18923 15521 18935 15555
rect 18877 15515 18935 15521
rect 19702 15512 19708 15564
rect 19760 15512 19766 15564
rect 19981 15555 20039 15561
rect 19981 15521 19993 15555
rect 20027 15521 20039 15555
rect 19981 15515 20039 15521
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15453 19671 15487
rect 19996 15484 20024 15515
rect 20438 15512 20444 15564
rect 20496 15512 20502 15564
rect 20640 15561 20668 15592
rect 20625 15555 20683 15561
rect 20625 15521 20637 15555
rect 20671 15521 20683 15555
rect 20625 15515 20683 15521
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15521 20775 15555
rect 20717 15515 20775 15521
rect 20855 15555 20913 15561
rect 20855 15521 20867 15555
rect 20901 15552 20913 15555
rect 20990 15552 20996 15564
rect 20901 15524 20996 15552
rect 20901 15521 20913 15524
rect 20855 15515 20913 15521
rect 20732 15484 20760 15515
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 21652 15561 21680 15592
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 27430 15620 27436 15632
rect 24044 15592 27436 15620
rect 21453 15555 21511 15561
rect 21453 15521 21465 15555
rect 21499 15521 21511 15555
rect 21453 15515 21511 15521
rect 21545 15555 21603 15561
rect 21545 15521 21557 15555
rect 21591 15521 21603 15555
rect 21545 15515 21603 15521
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15521 21695 15555
rect 21637 15515 21695 15521
rect 22005 15555 22063 15561
rect 22005 15521 22017 15555
rect 22051 15521 22063 15555
rect 22005 15515 22063 15521
rect 21082 15484 21088 15496
rect 19996 15456 20116 15484
rect 20732 15456 21088 15484
rect 19613 15447 19671 15453
rect 18322 15376 18328 15428
rect 18380 15416 18386 15428
rect 19628 15416 19656 15447
rect 19978 15416 19984 15428
rect 18380 15388 19984 15416
rect 18380 15376 18386 15388
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 17954 15348 17960 15360
rect 16960 15320 17960 15348
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 19702 15308 19708 15360
rect 19760 15348 19766 15360
rect 20088 15348 20116 15456
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 20898 15376 20904 15428
rect 20956 15416 20962 15428
rect 21468 15416 21496 15515
rect 21560 15484 21588 15515
rect 21818 15484 21824 15496
rect 21560 15456 21824 15484
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 22020 15484 22048 15515
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 24044 15552 24072 15592
rect 27430 15580 27436 15592
rect 27488 15580 27494 15632
rect 27798 15580 27804 15632
rect 27856 15620 27862 15632
rect 27856 15592 28028 15620
rect 27856 15580 27862 15592
rect 23992 15524 24072 15552
rect 24305 15555 24363 15561
rect 23992 15512 23998 15524
rect 24305 15521 24317 15555
rect 24351 15521 24363 15555
rect 24305 15515 24363 15521
rect 22278 15484 22284 15496
rect 22020 15456 22284 15484
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 23198 15444 23204 15496
rect 23256 15484 23262 15496
rect 24320 15484 24348 15515
rect 24394 15512 24400 15564
rect 24452 15552 24458 15564
rect 24946 15552 24952 15564
rect 24452 15524 24952 15552
rect 24452 15512 24458 15524
rect 24946 15512 24952 15524
rect 25004 15512 25010 15564
rect 25133 15555 25191 15561
rect 25133 15521 25145 15555
rect 25179 15552 25191 15555
rect 26694 15552 26700 15564
rect 25179 15524 26700 15552
rect 25179 15521 25191 15524
rect 25133 15515 25191 15521
rect 23256 15456 24348 15484
rect 23256 15444 23262 15456
rect 24578 15444 24584 15496
rect 24636 15484 24642 15496
rect 25148 15484 25176 15515
rect 26694 15512 26700 15524
rect 26752 15512 26758 15564
rect 26786 15512 26792 15564
rect 26844 15552 26850 15564
rect 27522 15552 27528 15564
rect 26844 15524 27528 15552
rect 26844 15512 26850 15524
rect 27522 15512 27528 15524
rect 27580 15552 27586 15564
rect 27709 15555 27767 15561
rect 27709 15552 27721 15555
rect 27580 15524 27721 15552
rect 27580 15512 27586 15524
rect 27709 15521 27721 15524
rect 27755 15521 27767 15555
rect 27709 15515 27767 15521
rect 27890 15512 27896 15564
rect 27948 15512 27954 15564
rect 28000 15561 28028 15592
rect 27985 15555 28043 15561
rect 27985 15521 27997 15555
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 28077 15555 28135 15561
rect 28077 15521 28089 15555
rect 28123 15552 28135 15555
rect 28166 15552 28172 15564
rect 28123 15524 28172 15552
rect 28123 15521 28135 15524
rect 28077 15515 28135 15521
rect 28166 15512 28172 15524
rect 28224 15512 28230 15564
rect 28276 15552 28304 15660
rect 28445 15657 28457 15691
rect 28491 15688 28503 15691
rect 28902 15688 28908 15700
rect 28491 15660 28908 15688
rect 28491 15657 28503 15660
rect 28445 15651 28503 15657
rect 28902 15648 28908 15660
rect 28960 15648 28966 15700
rect 28994 15648 29000 15700
rect 29052 15688 29058 15700
rect 29917 15691 29975 15697
rect 29917 15688 29929 15691
rect 29052 15660 29929 15688
rect 29052 15648 29058 15660
rect 29917 15657 29929 15660
rect 29963 15657 29975 15691
rect 29917 15651 29975 15657
rect 30282 15648 30288 15700
rect 30340 15688 30346 15700
rect 30377 15691 30435 15697
rect 30377 15688 30389 15691
rect 30340 15660 30389 15688
rect 30340 15648 30346 15660
rect 30377 15657 30389 15660
rect 30423 15657 30435 15691
rect 30377 15651 30435 15657
rect 28353 15623 28411 15629
rect 28353 15589 28365 15623
rect 28399 15620 28411 15623
rect 29558 15623 29616 15629
rect 29558 15620 29570 15623
rect 28399 15592 29570 15620
rect 28399 15589 28411 15592
rect 28353 15583 28411 15589
rect 29558 15589 29570 15592
rect 29604 15589 29616 15623
rect 29558 15583 29616 15589
rect 29270 15552 29276 15564
rect 28276 15524 29276 15552
rect 29270 15512 29276 15524
rect 29328 15552 29334 15564
rect 29328 15524 29776 15552
rect 29328 15512 29334 15524
rect 24636 15456 25176 15484
rect 26712 15484 26740 15512
rect 29748 15484 29776 15524
rect 29822 15512 29828 15564
rect 29880 15512 29886 15564
rect 30285 15555 30343 15561
rect 30285 15521 30297 15555
rect 30331 15552 30343 15555
rect 30742 15552 30748 15564
rect 30331 15524 30748 15552
rect 30331 15521 30343 15524
rect 30285 15515 30343 15521
rect 30742 15512 30748 15524
rect 30800 15512 30806 15564
rect 30469 15487 30527 15493
rect 30469 15484 30481 15487
rect 26712 15456 28028 15484
rect 29748 15456 30481 15484
rect 24636 15444 24642 15456
rect 28000 15428 28028 15456
rect 30469 15453 30481 15456
rect 30515 15453 30527 15487
rect 30469 15447 30527 15453
rect 20956 15388 21496 15416
rect 20956 15376 20962 15388
rect 22646 15376 22652 15428
rect 22704 15416 22710 15428
rect 27798 15416 27804 15428
rect 22704 15388 27804 15416
rect 22704 15376 22710 15388
rect 27798 15376 27804 15388
rect 27856 15376 27862 15428
rect 27982 15376 27988 15428
rect 28040 15376 28046 15428
rect 19760 15320 20116 15348
rect 19760 15308 19766 15320
rect 23290 15308 23296 15360
rect 23348 15348 23354 15360
rect 24026 15348 24032 15360
rect 23348 15320 24032 15348
rect 23348 15308 23354 15320
rect 24026 15308 24032 15320
rect 24084 15348 24090 15360
rect 24121 15351 24179 15357
rect 24121 15348 24133 15351
rect 24084 15320 24133 15348
rect 24084 15308 24090 15320
rect 24121 15317 24133 15320
rect 24167 15317 24179 15351
rect 24121 15311 24179 15317
rect 24854 15308 24860 15360
rect 24912 15348 24918 15360
rect 25041 15351 25099 15357
rect 25041 15348 25053 15351
rect 24912 15320 25053 15348
rect 24912 15308 24918 15320
rect 25041 15317 25053 15320
rect 25087 15317 25099 15351
rect 27816 15348 27844 15376
rect 28442 15348 28448 15360
rect 27816 15320 28448 15348
rect 25041 15311 25099 15317
rect 28442 15308 28448 15320
rect 28500 15348 28506 15360
rect 29178 15348 29184 15360
rect 28500 15320 29184 15348
rect 28500 15308 28506 15320
rect 29178 15308 29184 15320
rect 29236 15308 29242 15360
rect 552 15258 31648 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 11436 15258
rect 11488 15206 11500 15258
rect 11552 15206 11564 15258
rect 11616 15206 11628 15258
rect 11680 15206 11692 15258
rect 11744 15206 19210 15258
rect 19262 15206 19274 15258
rect 19326 15206 19338 15258
rect 19390 15206 19402 15258
rect 19454 15206 19466 15258
rect 19518 15206 26984 15258
rect 27036 15206 27048 15258
rect 27100 15206 27112 15258
rect 27164 15206 27176 15258
rect 27228 15206 27240 15258
rect 27292 15206 31648 15258
rect 552 15184 31648 15206
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 9858 15144 9864 15156
rect 9815 15116 9864 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 11606 15144 11612 15156
rect 10008 15116 11612 15144
rect 10008 15104 10014 15116
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12069 15147 12127 15153
rect 12069 15113 12081 15147
rect 12115 15113 12127 15147
rect 13722 15144 13728 15156
rect 12069 15107 12127 15113
rect 12176 15116 13728 15144
rect 4341 15079 4399 15085
rect 4341 15045 4353 15079
rect 4387 15076 4399 15079
rect 5626 15076 5632 15088
rect 4387 15048 5632 15076
rect 4387 15045 4399 15048
rect 4341 15039 4399 15045
rect 5626 15036 5632 15048
rect 5684 15036 5690 15088
rect 12084 15076 12112 15107
rect 11164 15048 12112 15076
rect 1394 14968 1400 15020
rect 1452 15008 1458 15020
rect 1581 15011 1639 15017
rect 1581 15008 1593 15011
rect 1452 14980 1593 15008
rect 1452 14968 1458 14980
rect 1581 14977 1593 14980
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 3326 14968 3332 15020
rect 3384 15008 3390 15020
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3384 14980 3709 15008
rect 3384 14968 3390 14980
rect 3697 14977 3709 14980
rect 3743 14977 3755 15011
rect 4065 15011 4123 15017
rect 4065 15008 4077 15011
rect 3697 14971 3755 14977
rect 3804 14980 4077 15008
rect 1302 14900 1308 14952
rect 1360 14900 1366 14952
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 1848 14875 1906 14881
rect 1848 14841 1860 14875
rect 1894 14872 1906 14875
rect 3237 14875 3295 14881
rect 3237 14872 3249 14875
rect 1894 14844 3249 14872
rect 1894 14841 1906 14844
rect 1848 14835 1906 14841
rect 3237 14841 3249 14844
rect 3283 14841 3295 14875
rect 3237 14835 3295 14841
rect 3436 14872 3464 14903
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 3804 14949 3832 14980
rect 4065 14977 4077 14980
rect 4111 14977 4123 15011
rect 4798 15008 4804 15020
rect 4065 14971 4123 14977
rect 4540 14980 4804 15008
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3568 14912 3617 14940
rect 3568 14900 3574 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 3970 14900 3976 14952
rect 4028 14900 4034 14952
rect 4540 14949 4568 14980
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 7101 15011 7159 15017
rect 7101 14977 7113 15011
rect 7147 15008 7159 15011
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 7147 14980 7297 15008
rect 7147 14977 7159 14980
rect 7101 14971 7159 14977
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 9950 15008 9956 15020
rect 7285 14971 7343 14977
rect 9416 14980 9956 15008
rect 4249 14943 4307 14949
rect 4249 14909 4261 14943
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 4154 14872 4160 14884
rect 3436 14844 4160 14872
rect 1397 14807 1455 14813
rect 1397 14773 1409 14807
rect 1443 14804 1455 14807
rect 1486 14804 1492 14816
rect 1443 14776 1492 14804
rect 1443 14773 1455 14776
rect 1397 14767 1455 14773
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 2961 14807 3019 14813
rect 2961 14773 2973 14807
rect 3007 14804 3019 14807
rect 3436 14804 3464 14844
rect 4154 14832 4160 14844
rect 4212 14832 4218 14884
rect 3007 14776 3464 14804
rect 4264 14804 4292 14903
rect 4448 14872 4476 14903
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 4709 14943 4767 14949
rect 4709 14940 4721 14943
rect 4672 14912 4721 14940
rect 4672 14900 4678 14912
rect 4709 14909 4721 14912
rect 4755 14940 4767 14943
rect 4890 14940 4896 14952
rect 4755 14912 4896 14940
rect 4755 14909 4767 14912
rect 4709 14903 4767 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 5592 14912 7205 14940
rect 5592 14900 5598 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 5166 14872 5172 14884
rect 4448 14844 5172 14872
rect 5166 14832 5172 14844
rect 5224 14832 5230 14884
rect 6822 14832 6828 14884
rect 6880 14881 6886 14884
rect 6880 14872 6892 14881
rect 8956 14872 8984 14903
rect 9306 14900 9312 14952
rect 9364 14900 9370 14952
rect 9416 14949 9444 14980
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 11164 15017 11192 15048
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 14977 11207 15011
rect 12176 15008 12204 15116
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 13998 15104 14004 15156
rect 14056 15104 14062 15156
rect 16666 15104 16672 15156
rect 16724 15144 16730 15156
rect 16942 15144 16948 15156
rect 16724 15116 16948 15144
rect 16724 15104 16730 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17034 15104 17040 15156
rect 17092 15104 17098 15156
rect 17773 15147 17831 15153
rect 17773 15113 17785 15147
rect 17819 15113 17831 15147
rect 17773 15107 17831 15113
rect 17957 15147 18015 15153
rect 17957 15113 17969 15147
rect 18003 15144 18015 15147
rect 18138 15144 18144 15156
rect 18003 15116 18144 15144
rect 18003 15113 18015 15116
rect 17957 15107 18015 15113
rect 11149 14971 11207 14977
rect 11532 14980 12204 15008
rect 12406 15048 12756 15076
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 9490 14900 9496 14952
rect 9548 14900 9554 14952
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 11054 14940 11060 14952
rect 9784 14912 11060 14940
rect 9784 14872 9812 14912
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11532 14949 11560 14980
rect 11517 14943 11575 14949
rect 11517 14909 11529 14943
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 11606 14900 11612 14952
rect 11664 14900 11670 14952
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14940 11759 14943
rect 11790 14940 11796 14952
rect 11747 14912 11796 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 11885 14943 11943 14949
rect 11885 14909 11897 14943
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 6880 14844 6925 14872
rect 8956 14844 9812 14872
rect 10904 14875 10962 14881
rect 6880 14835 6892 14844
rect 10904 14841 10916 14875
rect 10950 14872 10962 14875
rect 11241 14875 11299 14881
rect 11241 14872 11253 14875
rect 10950 14844 11253 14872
rect 10950 14841 10962 14844
rect 10904 14835 10962 14841
rect 11241 14841 11253 14844
rect 11287 14841 11299 14875
rect 11241 14835 11299 14841
rect 6880 14832 6886 14835
rect 4706 14804 4712 14816
rect 4264 14776 4712 14804
rect 3007 14773 3019 14776
rect 2961 14767 3019 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5350 14764 5356 14816
rect 5408 14764 5414 14816
rect 5721 14807 5779 14813
rect 5721 14773 5733 14807
rect 5767 14804 5779 14807
rect 6546 14804 6552 14816
rect 5767 14776 6552 14804
rect 5767 14773 5779 14776
rect 5721 14767 5779 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 8846 14764 8852 14816
rect 8904 14764 8910 14816
rect 9030 14764 9036 14816
rect 9088 14764 9094 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 11900 14804 11928 14903
rect 11974 14900 11980 14952
rect 12032 14940 12038 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 12032 14912 12173 14940
rect 12032 14900 12038 14912
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 12161 14903 12219 14909
rect 12406 14804 12434 15048
rect 12728 15008 12756 15048
rect 13446 15008 13452 15020
rect 12728 14980 13452 15008
rect 12728 14949 12756 14980
rect 13446 14968 13452 14980
rect 13504 15008 13510 15020
rect 13722 15008 13728 15020
rect 13504 14980 13728 15008
rect 13504 14968 13510 14980
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 17788 15008 17816 15107
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 19242 15144 19248 15156
rect 18248 15116 19248 15144
rect 18248 15076 18276 15116
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 19337 15147 19395 15153
rect 19337 15113 19349 15147
rect 19383 15144 19395 15147
rect 19610 15144 19616 15156
rect 19383 15116 19616 15144
rect 19383 15113 19395 15116
rect 19337 15107 19395 15113
rect 19610 15104 19616 15116
rect 19668 15104 19674 15156
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20714 15144 20720 15156
rect 19935 15116 20720 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 17972 15048 18276 15076
rect 17972 15008 18000 15048
rect 18138 15008 18144 15020
rect 16684 14980 17448 15008
rect 17788 14980 18000 15008
rect 18055 14980 18144 15008
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 12894 14900 12900 14952
rect 12952 14900 12958 14952
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14940 13139 14943
rect 13262 14940 13268 14952
rect 13127 14912 13268 14940
rect 13127 14909 13139 14912
rect 13081 14903 13139 14909
rect 13004 14872 13032 14903
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 14366 14949 14372 14952
rect 14360 14940 14372 14949
rect 13688 14912 13952 14940
rect 14327 14912 14372 14940
rect 13688 14900 13694 14912
rect 13170 14872 13176 14884
rect 13004 14844 13176 14872
rect 13170 14832 13176 14844
rect 13228 14872 13234 14884
rect 13228 14844 13768 14872
rect 13228 14832 13234 14844
rect 9732 14776 12434 14804
rect 9732 14764 9738 14776
rect 13354 14764 13360 14816
rect 13412 14764 13418 14816
rect 13740 14804 13768 14844
rect 13814 14832 13820 14884
rect 13872 14832 13878 14884
rect 13924 14872 13952 14912
rect 14360 14903 14372 14912
rect 14366 14900 14372 14903
rect 14424 14900 14430 14952
rect 16684 14949 16712 14980
rect 17420 14952 17448 14980
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 15488 14912 15577 14940
rect 14458 14872 14464 14884
rect 13924 14844 14464 14872
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 14182 14804 14188 14816
rect 13740 14776 14188 14804
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 15488 14813 15516 14912
rect 15565 14909 15577 14912
rect 15611 14909 15623 14943
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 15565 14903 15623 14909
rect 15764 14912 16313 14940
rect 15764 14816 15792 14912
rect 16301 14909 16313 14912
rect 16347 14909 16359 14943
rect 16301 14903 16359 14909
rect 16669 14943 16727 14949
rect 16669 14909 16681 14943
rect 16715 14909 16727 14943
rect 16669 14903 16727 14909
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 16868 14872 16896 14903
rect 16942 14900 16948 14952
rect 17000 14940 17006 14952
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 17000 14912 17325 14940
rect 17000 14900 17006 14912
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 17402 14900 17408 14952
rect 17460 14900 17466 14952
rect 18055 14949 18083 14980
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18248 14949 18276 15048
rect 18966 15036 18972 15088
rect 19024 15076 19030 15088
rect 19904 15076 19932 15107
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 21358 15104 21364 15156
rect 21416 15104 21422 15156
rect 21729 15147 21787 15153
rect 21729 15113 21741 15147
rect 21775 15144 21787 15147
rect 23198 15144 23204 15156
rect 21775 15116 23204 15144
rect 21775 15113 21787 15116
rect 21729 15107 21787 15113
rect 23198 15104 23204 15116
rect 23256 15104 23262 15156
rect 23658 15104 23664 15156
rect 23716 15144 23722 15156
rect 25406 15144 25412 15156
rect 23716 15116 25412 15144
rect 23716 15104 23722 15116
rect 25406 15104 25412 15116
rect 25464 15104 25470 15156
rect 25498 15104 25504 15156
rect 25556 15144 25562 15156
rect 26145 15147 26203 15153
rect 26145 15144 26157 15147
rect 25556 15116 26157 15144
rect 25556 15104 25562 15116
rect 26145 15113 26157 15116
rect 26191 15113 26203 15147
rect 26145 15107 26203 15113
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 28261 15147 28319 15153
rect 28261 15144 28273 15147
rect 27948 15116 28273 15144
rect 27948 15104 27954 15116
rect 28261 15113 28273 15116
rect 28307 15113 28319 15147
rect 28718 15144 28724 15156
rect 28261 15107 28319 15113
rect 28368 15116 28724 15144
rect 19024 15048 19104 15076
rect 19024 15036 19030 15048
rect 17773 14943 17831 14949
rect 17773 14909 17785 14943
rect 17819 14909 17831 14943
rect 17773 14903 17831 14909
rect 18037 14943 18095 14949
rect 18037 14909 18049 14943
rect 18083 14909 18095 14943
rect 18037 14903 18095 14909
rect 18233 14943 18291 14949
rect 18233 14909 18245 14943
rect 18279 14940 18291 14943
rect 18598 14940 18604 14952
rect 18279 14912 18604 14940
rect 18279 14909 18291 14912
rect 18233 14903 18291 14909
rect 17494 14872 17500 14884
rect 16500 14844 17500 14872
rect 15473 14807 15531 14813
rect 15473 14773 15485 14807
rect 15519 14773 15531 14807
rect 15473 14767 15531 14773
rect 15746 14764 15752 14816
rect 15804 14764 15810 14816
rect 16500 14813 16528 14844
rect 17494 14832 17500 14844
rect 17552 14872 17558 14884
rect 17788 14872 17816 14903
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 18782 14900 18788 14952
rect 18840 14900 18846 14952
rect 18966 14949 18972 14952
rect 18923 14943 18972 14949
rect 18923 14909 18935 14943
rect 18969 14909 18972 14943
rect 18923 14903 18972 14909
rect 18966 14900 18972 14903
rect 19024 14900 19030 14952
rect 19076 14949 19104 15048
rect 19148 15048 19932 15076
rect 19148 14950 19176 15048
rect 19978 15036 19984 15088
rect 20036 15076 20042 15088
rect 20073 15079 20131 15085
rect 20073 15076 20085 15079
rect 20036 15048 20085 15076
rect 20036 15036 20042 15048
rect 20073 15045 20085 15048
rect 20119 15045 20131 15079
rect 20073 15039 20131 15045
rect 23474 15036 23480 15088
rect 23532 15076 23538 15088
rect 25590 15076 25596 15088
rect 23532 15048 25596 15076
rect 23532 15036 23538 15048
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 19797 15011 19855 15017
rect 19797 15008 19809 15011
rect 19300 14980 19809 15008
rect 19300 14968 19306 14980
rect 19797 14977 19809 14980
rect 19843 14977 19855 15011
rect 19797 14971 19855 14977
rect 19996 14980 21404 15008
rect 19148 14949 19196 14950
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14909 19119 14943
rect 19148 14943 19216 14949
rect 19148 14922 19170 14943
rect 19061 14903 19119 14909
rect 19158 14909 19170 14922
rect 19204 14909 19216 14943
rect 19158 14903 19216 14909
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19900 14943 19958 14949
rect 19392 14912 19748 14940
rect 19392 14900 19398 14912
rect 19613 14875 19671 14881
rect 19613 14872 19625 14875
rect 17552 14844 19625 14872
rect 17552 14832 17558 14844
rect 19613 14841 19625 14844
rect 19659 14841 19671 14875
rect 19720 14872 19748 14912
rect 19900 14909 19912 14943
rect 19946 14940 19958 14943
rect 19996 14940 20024 14980
rect 20916 14949 20944 14980
rect 21376 14952 21404 14980
rect 22738 14968 22744 15020
rect 22796 15008 22802 15020
rect 22796 14980 24348 15008
rect 22796 14968 22802 14980
rect 20809 14943 20867 14949
rect 20809 14940 20821 14943
rect 19946 14912 20024 14940
rect 20088 14912 20821 14940
rect 19946 14909 19958 14912
rect 19900 14903 19958 14909
rect 20088 14872 20116 14912
rect 20809 14909 20821 14912
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 20901 14943 20959 14949
rect 20901 14909 20913 14943
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 21082 14900 21088 14952
rect 21140 14900 21146 14952
rect 21358 14900 21364 14952
rect 21416 14900 21422 14952
rect 21545 14943 21603 14949
rect 21545 14909 21557 14943
rect 21591 14940 21603 14943
rect 22094 14940 22100 14952
rect 21591 14912 22100 14940
rect 21591 14909 21603 14912
rect 21545 14903 21603 14909
rect 19720 14844 20116 14872
rect 20349 14875 20407 14881
rect 19613 14835 19671 14841
rect 20349 14841 20361 14875
rect 20395 14872 20407 14875
rect 20622 14872 20628 14884
rect 20395 14844 20628 14872
rect 20395 14841 20407 14844
rect 20349 14835 20407 14841
rect 16485 14807 16543 14813
rect 16485 14773 16497 14807
rect 16531 14773 16543 14807
rect 16485 14767 16543 14773
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 17678 14804 17684 14816
rect 17000 14776 17684 14804
rect 17000 14764 17006 14776
rect 17678 14764 17684 14776
rect 17736 14764 17742 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18141 14807 18199 14813
rect 18141 14804 18153 14807
rect 18012 14776 18153 14804
rect 18012 14764 18018 14776
rect 18141 14773 18153 14776
rect 18187 14804 18199 14807
rect 19150 14804 19156 14816
rect 18187 14776 19156 14804
rect 18187 14773 18199 14776
rect 18141 14767 18199 14773
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 19628 14804 19656 14835
rect 20622 14832 20628 14844
rect 20680 14832 20686 14884
rect 20990 14832 20996 14884
rect 21048 14872 21054 14884
rect 21269 14875 21327 14881
rect 21269 14872 21281 14875
rect 21048 14844 21281 14872
rect 21048 14832 21054 14844
rect 21269 14841 21281 14844
rect 21315 14841 21327 14875
rect 21560 14872 21588 14903
rect 22094 14900 22100 14912
rect 22152 14900 22158 14952
rect 23658 14900 23664 14952
rect 23716 14900 23722 14952
rect 24026 14900 24032 14952
rect 24084 14900 24090 14952
rect 24121 14943 24179 14949
rect 24121 14909 24133 14943
rect 24167 14940 24179 14943
rect 24210 14940 24216 14952
rect 24167 14912 24216 14940
rect 24167 14909 24179 14912
rect 24121 14903 24179 14909
rect 24210 14900 24216 14912
rect 24268 14900 24274 14952
rect 24320 14949 24348 14980
rect 24412 14949 24440 15048
rect 25590 15036 25596 15048
rect 25648 15076 25654 15088
rect 26234 15076 26240 15088
rect 25648 15048 26240 15076
rect 25648 15036 25654 15048
rect 26234 15036 26240 15048
rect 26292 15036 26298 15088
rect 28368 15076 28396 15116
rect 28718 15104 28724 15116
rect 28776 15104 28782 15156
rect 30377 15147 30435 15153
rect 30377 15144 30389 15147
rect 29104 15116 30389 15144
rect 28994 15076 29000 15088
rect 28184 15048 28396 15076
rect 28460 15048 29000 15076
rect 28184 15020 28212 15048
rect 25498 15008 25504 15020
rect 25056 14980 25504 15008
rect 24305 14943 24363 14949
rect 24305 14909 24317 14943
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24397 14943 24455 14949
rect 24397 14909 24409 14943
rect 24443 14909 24455 14943
rect 24397 14903 24455 14909
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 24857 14943 24915 14949
rect 24857 14909 24869 14943
rect 24903 14909 24915 14943
rect 24857 14903 24915 14909
rect 21269 14835 21327 14841
rect 21376 14844 21588 14872
rect 20714 14804 20720 14816
rect 19628 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14804 20778 14816
rect 21376 14804 21404 14844
rect 23474 14832 23480 14884
rect 23532 14832 23538 14884
rect 23750 14832 23756 14884
rect 23808 14872 23814 14884
rect 24688 14872 24716 14900
rect 23808 14844 24716 14872
rect 23808 14832 23814 14844
rect 20772 14776 21404 14804
rect 20772 14764 20778 14776
rect 21542 14764 21548 14816
rect 21600 14804 21606 14816
rect 22646 14804 22652 14816
rect 21600 14776 22652 14804
rect 21600 14764 21606 14776
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 23293 14807 23351 14813
rect 23293 14773 23305 14807
rect 23339 14804 23351 14807
rect 23382 14804 23388 14816
rect 23339 14776 23388 14804
rect 23339 14773 23351 14776
rect 23293 14767 23351 14773
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 23566 14764 23572 14816
rect 23624 14804 23630 14816
rect 23845 14807 23903 14813
rect 23845 14804 23857 14807
rect 23624 14776 23857 14804
rect 23624 14764 23630 14776
rect 23845 14773 23857 14776
rect 23891 14773 23903 14807
rect 24872 14804 24900 14903
rect 24946 14900 24952 14952
rect 25004 14900 25010 14952
rect 25056 14949 25084 14980
rect 25498 14968 25504 14980
rect 25556 14968 25562 15020
rect 28166 15008 28172 15020
rect 27264 14980 28172 15008
rect 25041 14943 25099 14949
rect 25041 14909 25053 14943
rect 25087 14909 25099 14943
rect 25041 14903 25099 14909
rect 25222 14900 25228 14952
rect 25280 14940 25286 14952
rect 25639 14943 25697 14949
rect 25639 14940 25651 14943
rect 25280 14912 25651 14940
rect 25280 14900 25286 14912
rect 25639 14909 25651 14912
rect 25685 14909 25697 14943
rect 25639 14903 25697 14909
rect 25777 14943 25835 14949
rect 25777 14909 25789 14943
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 25038 14804 25044 14816
rect 24872 14776 25044 14804
rect 23845 14767 23903 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 25314 14764 25320 14816
rect 25372 14764 25378 14816
rect 25409 14807 25467 14813
rect 25409 14773 25421 14807
rect 25455 14804 25467 14807
rect 25498 14804 25504 14816
rect 25455 14776 25504 14804
rect 25455 14773 25467 14776
rect 25409 14767 25467 14773
rect 25498 14764 25504 14776
rect 25556 14764 25562 14816
rect 25792 14804 25820 14903
rect 25866 14900 25872 14952
rect 25924 14900 25930 14952
rect 26050 14900 26056 14952
rect 26108 14900 26114 14952
rect 26694 14900 26700 14952
rect 26752 14940 26758 14952
rect 27264 14949 27292 14980
rect 28166 14968 28172 14980
rect 28224 14968 28230 15020
rect 27157 14943 27215 14949
rect 27157 14940 27169 14943
rect 26752 14912 27169 14940
rect 26752 14900 26758 14912
rect 27157 14909 27169 14912
rect 27203 14909 27215 14943
rect 27157 14903 27215 14909
rect 27249 14943 27307 14949
rect 27249 14909 27261 14943
rect 27295 14909 27307 14943
rect 27249 14903 27307 14909
rect 27341 14943 27399 14949
rect 27341 14909 27353 14943
rect 27387 14940 27399 14943
rect 27430 14940 27436 14952
rect 27387 14912 27436 14940
rect 27387 14909 27399 14912
rect 27341 14903 27399 14909
rect 27264 14872 27292 14903
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 27522 14900 27528 14952
rect 27580 14900 27586 14952
rect 28258 14940 28264 14952
rect 27816 14912 28264 14940
rect 27816 14881 27844 14912
rect 28258 14900 28264 14912
rect 28316 14900 28322 14952
rect 28460 14949 28488 15048
rect 28994 15036 29000 15048
rect 29052 15036 29058 15088
rect 29104 15008 29132 15116
rect 30377 15113 30389 15116
rect 30423 15113 30435 15147
rect 30377 15107 30435 15113
rect 29454 15008 29460 15020
rect 28736 14980 29132 15008
rect 29288 14980 29460 15008
rect 28445 14943 28503 14949
rect 28445 14909 28457 14943
rect 28491 14909 28503 14943
rect 28445 14903 28503 14909
rect 28534 14900 28540 14952
rect 28592 14900 28598 14952
rect 28736 14949 28764 14980
rect 28721 14943 28779 14949
rect 28721 14909 28733 14943
rect 28767 14909 28779 14943
rect 28721 14903 28779 14909
rect 28810 14900 28816 14952
rect 28868 14900 28874 14952
rect 28997 14943 29055 14949
rect 28997 14909 29009 14943
rect 29043 14909 29055 14943
rect 28997 14903 29055 14909
rect 27801 14875 27859 14881
rect 27801 14872 27813 14875
rect 26252 14844 27292 14872
rect 27448 14844 27813 14872
rect 25958 14804 25964 14816
rect 25792 14776 25964 14804
rect 25958 14764 25964 14776
rect 26016 14804 26022 14816
rect 26252 14804 26280 14844
rect 27448 14816 27476 14844
rect 27801 14841 27813 14844
rect 27847 14841 27859 14875
rect 27801 14835 27859 14841
rect 27985 14875 28043 14881
rect 27985 14841 27997 14875
rect 28031 14841 28043 14875
rect 27985 14835 28043 14841
rect 28169 14875 28227 14881
rect 28169 14841 28181 14875
rect 28215 14872 28227 14875
rect 29012 14872 29040 14903
rect 29086 14900 29092 14952
rect 29144 14940 29150 14952
rect 29288 14949 29316 14980
rect 29454 14968 29460 14980
rect 29512 15008 29518 15020
rect 29512 14980 30052 15008
rect 29512 14968 29518 14980
rect 29181 14943 29239 14949
rect 29181 14940 29193 14943
rect 29144 14912 29193 14940
rect 29144 14900 29150 14912
rect 29181 14909 29193 14912
rect 29227 14909 29239 14943
rect 29181 14903 29239 14909
rect 29273 14943 29331 14949
rect 29273 14909 29285 14943
rect 29319 14909 29331 14943
rect 29273 14903 29331 14909
rect 29365 14943 29423 14949
rect 29365 14909 29377 14943
rect 29411 14937 29423 14943
rect 29546 14940 29552 14952
rect 29472 14937 29552 14940
rect 29411 14912 29552 14937
rect 29411 14909 29500 14912
rect 29365 14903 29423 14909
rect 28215 14844 29040 14872
rect 29196 14872 29224 14903
rect 29546 14900 29552 14912
rect 29604 14900 29610 14952
rect 29730 14900 29736 14952
rect 29788 14900 29794 14952
rect 30024 14949 30052 14980
rect 29917 14943 29975 14949
rect 29917 14909 29929 14943
rect 29963 14909 29975 14943
rect 29917 14903 29975 14909
rect 30009 14943 30067 14949
rect 30009 14909 30021 14943
rect 30055 14909 30067 14943
rect 30009 14903 30067 14909
rect 30101 14943 30159 14949
rect 30101 14909 30113 14943
rect 30147 14940 30159 14943
rect 30742 14940 30748 14952
rect 30147 14912 30748 14940
rect 30147 14909 30159 14912
rect 30101 14903 30159 14909
rect 29932 14872 29960 14903
rect 30742 14900 30748 14912
rect 30800 14900 30806 14952
rect 29196 14844 29960 14872
rect 28215 14841 28227 14844
rect 28169 14835 28227 14841
rect 26016 14776 26280 14804
rect 26016 14764 26022 14776
rect 26602 14764 26608 14816
rect 26660 14804 26666 14816
rect 26881 14807 26939 14813
rect 26881 14804 26893 14807
rect 26660 14776 26893 14804
rect 26660 14764 26666 14776
rect 26881 14773 26893 14776
rect 26927 14773 26939 14807
rect 26881 14767 26939 14773
rect 27430 14764 27436 14816
rect 27488 14764 27494 14816
rect 28000 14804 28028 14835
rect 28902 14804 28908 14816
rect 28000 14776 28908 14804
rect 28902 14764 28908 14776
rect 28960 14764 28966 14816
rect 29638 14764 29644 14816
rect 29696 14764 29702 14816
rect 29932 14804 29960 14844
rect 30098 14804 30104 14816
rect 29932 14776 30104 14804
rect 30098 14764 30104 14776
rect 30156 14764 30162 14816
rect 552 14714 31648 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 12096 14714
rect 12148 14662 12160 14714
rect 12212 14662 12224 14714
rect 12276 14662 12288 14714
rect 12340 14662 12352 14714
rect 12404 14662 19870 14714
rect 19922 14662 19934 14714
rect 19986 14662 19998 14714
rect 20050 14662 20062 14714
rect 20114 14662 20126 14714
rect 20178 14662 27644 14714
rect 27696 14662 27708 14714
rect 27760 14662 27772 14714
rect 27824 14662 27836 14714
rect 27888 14662 27900 14714
rect 27952 14662 31648 14714
rect 552 14640 31648 14662
rect 2869 14603 2927 14609
rect 2869 14569 2881 14603
rect 2915 14600 2927 14603
rect 2915 14572 4108 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 4080 14544 4108 14572
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 4856 14572 5089 14600
rect 4856 14560 4862 14572
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 5350 14560 5356 14612
rect 5408 14600 5414 14612
rect 6273 14603 6331 14609
rect 6273 14600 6285 14603
rect 5408 14572 6285 14600
rect 5408 14560 5414 14572
rect 6273 14569 6285 14572
rect 6319 14569 6331 14603
rect 6273 14563 6331 14569
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 7055 14572 12296 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 1578 14492 1584 14544
rect 1636 14532 1642 14544
rect 1734 14535 1792 14541
rect 1734 14532 1746 14535
rect 1636 14504 1746 14532
rect 1636 14492 1642 14504
rect 1734 14501 1746 14504
rect 1780 14501 1792 14535
rect 1734 14495 1792 14501
rect 2958 14492 2964 14544
rect 3016 14532 3022 14544
rect 3418 14532 3424 14544
rect 3016 14504 3424 14532
rect 3016 14492 3022 14504
rect 1486 14424 1492 14476
rect 1544 14424 1550 14476
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 3160 14473 3188 14504
rect 3418 14492 3424 14504
rect 3476 14532 3482 14544
rect 3970 14532 3976 14544
rect 3476 14504 3976 14532
rect 3476 14492 3482 14504
rect 3970 14492 3976 14504
rect 4028 14492 4034 14544
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 4120 14504 8432 14532
rect 4120 14492 4126 14504
rect 3053 14467 3111 14473
rect 3053 14464 3065 14467
rect 2832 14436 3065 14464
rect 2832 14424 2838 14436
rect 3053 14433 3065 14436
rect 3099 14433 3111 14467
rect 3053 14427 3111 14433
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 7098 14464 7104 14476
rect 3145 14427 3203 14433
rect 4080 14436 7104 14464
rect 3068 14396 3096 14427
rect 4080 14408 4108 14436
rect 3510 14396 3516 14408
rect 3068 14368 3516 14396
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 6362 14356 6368 14408
rect 6420 14356 6426 14408
rect 6472 14405 6500 14436
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 7300 14405 7328 14504
rect 8404 14473 8432 14504
rect 9030 14492 9036 14544
rect 9088 14532 9094 14544
rect 9462 14535 9520 14541
rect 9462 14532 9474 14535
rect 9088 14504 9474 14532
rect 9088 14492 9094 14504
rect 9462 14501 9474 14504
rect 9508 14501 9520 14535
rect 9462 14495 9520 14501
rect 11606 14492 11612 14544
rect 11664 14532 11670 14544
rect 12268 14541 12296 14572
rect 12894 14560 12900 14612
rect 12952 14600 12958 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 12952 14572 13277 14600
rect 12952 14560 12958 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14884 14572 15117 14600
rect 14884 14560 14890 14572
rect 15105 14569 15117 14572
rect 15151 14600 15163 14603
rect 17497 14603 17555 14609
rect 15151 14572 15332 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 12069 14535 12127 14541
rect 12069 14532 12081 14535
rect 11664 14504 12081 14532
rect 11664 14492 11670 14504
rect 12069 14501 12081 14504
rect 12115 14501 12127 14535
rect 12069 14495 12127 14501
rect 12253 14535 12311 14541
rect 12253 14501 12265 14535
rect 12299 14532 12311 14535
rect 12299 14504 12664 14532
rect 12299 14501 12311 14504
rect 12253 14495 12311 14501
rect 12636 14476 12664 14504
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 13970 14535 14028 14541
rect 13970 14532 13982 14535
rect 13412 14504 13982 14532
rect 13412 14492 13418 14504
rect 13970 14501 13982 14504
rect 14016 14501 14028 14535
rect 15304 14532 15332 14572
rect 17497 14569 17509 14603
rect 17543 14600 17555 14603
rect 17586 14600 17592 14612
rect 17543 14572 17592 14600
rect 17543 14569 17555 14572
rect 17497 14563 17555 14569
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 17678 14560 17684 14612
rect 17736 14600 17742 14612
rect 18785 14603 18843 14609
rect 17736 14572 18184 14600
rect 17736 14560 17742 14572
rect 15304 14504 16804 14532
rect 13970 14495 14028 14501
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 8389 14467 8447 14473
rect 7423 14436 7972 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 7944 14408 7972 14436
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 8846 14424 8852 14476
rect 8904 14464 8910 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 8904 14436 9229 14464
rect 8904 14424 8910 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 11790 14464 11796 14476
rect 9217 14427 9275 14433
rect 9324 14436 11796 14464
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6604 14368 6837 14396
rect 6604 14356 6610 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 3050 14288 3056 14340
rect 3108 14288 3114 14340
rect 4893 14331 4951 14337
rect 4893 14297 4905 14331
rect 4939 14328 4951 14331
rect 4982 14328 4988 14340
rect 4939 14300 4988 14328
rect 4939 14297 4951 14300
rect 4893 14291 4951 14297
rect 4982 14288 4988 14300
rect 5040 14288 5046 14340
rect 5350 14288 5356 14340
rect 5408 14328 5414 14340
rect 5445 14331 5503 14337
rect 5445 14328 5457 14331
rect 5408 14300 5457 14328
rect 5408 14288 5414 14300
rect 5445 14297 5457 14300
rect 5491 14297 5503 14331
rect 6840 14328 6868 14359
rect 7852 14328 7880 14359
rect 7926 14356 7932 14408
rect 7984 14356 7990 14408
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14396 8263 14399
rect 9324 14396 9352 14436
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 12483 14436 12541 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12529 14433 12541 14436
rect 12575 14433 12587 14467
rect 12529 14427 12587 14433
rect 8251 14368 9352 14396
rect 11517 14399 11575 14405
rect 8251 14365 8263 14368
rect 8205 14359 8263 14365
rect 11517 14365 11529 14399
rect 11563 14365 11575 14399
rect 12452 14396 12480 14427
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12676 14436 12725 14464
rect 12676 14424 12682 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 12713 14427 12771 14433
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13449 14467 13507 14473
rect 13449 14464 13461 14467
rect 13044 14436 13461 14464
rect 13044 14424 13050 14436
rect 13449 14433 13461 14436
rect 13495 14433 13507 14467
rect 13449 14427 13507 14433
rect 13630 14424 13636 14476
rect 13688 14424 13694 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 14550 14464 14556 14476
rect 13872 14436 14556 14464
rect 13872 14424 13878 14436
rect 14550 14424 14556 14436
rect 14608 14464 14614 14476
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 14608 14436 15209 14464
rect 14608 14424 14614 14436
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 15351 14467 15409 14473
rect 15351 14433 15363 14467
rect 15397 14464 15409 14467
rect 15746 14464 15752 14476
rect 15397 14436 15752 14464
rect 15397 14433 15409 14436
rect 15351 14427 15409 14433
rect 13078 14396 13084 14408
rect 12452 14368 13084 14396
rect 11517 14359 11575 14365
rect 6840 14300 7880 14328
rect 5445 14291 5503 14297
rect 10502 14288 10508 14340
rect 10560 14328 10566 14340
rect 10597 14331 10655 14337
rect 10597 14328 10609 14331
rect 10560 14300 10609 14328
rect 10560 14288 10566 14300
rect 10597 14297 10609 14300
rect 10643 14328 10655 14331
rect 11532 14328 11560 14359
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13722 14356 13728 14408
rect 13780 14356 13786 14408
rect 10643 14300 11560 14328
rect 10643 14297 10655 14300
rect 10597 14291 10655 14297
rect 12526 14288 12532 14340
rect 12584 14288 12590 14340
rect 15212 14328 15240 14427
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 16776 14473 16804 14504
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14433 16819 14467
rect 16761 14427 16819 14433
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17218 14464 17224 14476
rect 17175 14436 17224 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14396 15623 14399
rect 16574 14396 16580 14408
rect 15611 14368 16580 14396
rect 15611 14365 15623 14368
rect 15565 14359 15623 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 17144 14396 17172 14427
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 17494 14424 17500 14476
rect 17552 14464 17558 14476
rect 17681 14467 17739 14473
rect 17681 14464 17693 14467
rect 17552 14436 17693 14464
rect 17552 14424 17558 14436
rect 17681 14433 17693 14436
rect 17727 14464 17739 14467
rect 17954 14464 17960 14476
rect 17727 14436 17960 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 18156 14473 18184 14572
rect 18785 14569 18797 14603
rect 18831 14600 18843 14603
rect 19702 14600 19708 14612
rect 18831 14572 19708 14600
rect 18831 14569 18843 14572
rect 18785 14563 18843 14569
rect 19702 14560 19708 14572
rect 19760 14600 19766 14612
rect 20993 14603 21051 14609
rect 19760 14572 20668 14600
rect 19760 14560 19766 14572
rect 18506 14492 18512 14544
rect 18564 14532 18570 14544
rect 19610 14532 19616 14544
rect 18564 14504 19616 14532
rect 18564 14492 18570 14504
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 19797 14535 19855 14541
rect 19797 14501 19809 14535
rect 19843 14532 19855 14535
rect 19886 14532 19892 14544
rect 19843 14504 19892 14532
rect 19843 14501 19855 14504
rect 19797 14495 19855 14501
rect 19886 14492 19892 14504
rect 19944 14492 19950 14544
rect 20530 14492 20536 14544
rect 20588 14492 20594 14544
rect 18141 14467 18199 14473
rect 18141 14433 18153 14467
rect 18187 14433 18199 14467
rect 18141 14427 18199 14433
rect 16684 14368 17172 14396
rect 16684 14328 16712 14368
rect 17770 14356 17776 14408
rect 17828 14356 17834 14408
rect 18156 14396 18184 14427
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 18288 14436 18429 14464
rect 18288 14424 18294 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 18598 14424 18604 14476
rect 18656 14424 18662 14476
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14464 20039 14467
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 20027 14436 20085 14464
rect 20027 14433 20039 14436
rect 19981 14427 20039 14433
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 18506 14396 18512 14408
rect 18156 14368 18512 14396
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 20088 14396 20116 14427
rect 20254 14424 20260 14476
rect 20312 14424 20318 14476
rect 20548 14464 20576 14492
rect 20364 14436 20576 14464
rect 20364 14396 20392 14436
rect 20088 14368 20392 14396
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14365 20591 14399
rect 20640 14396 20668 14572
rect 20993 14569 21005 14603
rect 21039 14600 21051 14603
rect 21542 14600 21548 14612
rect 21039 14572 21548 14600
rect 21039 14569 21051 14572
rect 20993 14563 21051 14569
rect 21542 14560 21548 14572
rect 21600 14560 21606 14612
rect 21652 14572 23060 14600
rect 21082 14492 21088 14544
rect 21140 14532 21146 14544
rect 21652 14532 21680 14572
rect 22557 14535 22615 14541
rect 22557 14532 22569 14535
rect 21140 14504 21680 14532
rect 21836 14504 22569 14532
rect 21140 14492 21146 14504
rect 20714 14424 20720 14476
rect 20772 14424 20778 14476
rect 21358 14424 21364 14476
rect 21416 14464 21422 14476
rect 21836 14473 21864 14504
rect 22557 14501 22569 14504
rect 22603 14501 22615 14535
rect 22557 14495 22615 14501
rect 22738 14492 22744 14544
rect 22796 14492 22802 14544
rect 23032 14532 23060 14572
rect 23474 14560 23480 14612
rect 23532 14600 23538 14612
rect 23753 14603 23811 14609
rect 23753 14600 23765 14603
rect 23532 14572 23765 14600
rect 23532 14560 23538 14572
rect 23753 14569 23765 14572
rect 23799 14600 23811 14603
rect 23799 14572 23980 14600
rect 23799 14569 23811 14572
rect 23753 14563 23811 14569
rect 23845 14535 23903 14541
rect 23845 14532 23857 14535
rect 23032 14504 23857 14532
rect 21821 14467 21879 14473
rect 21821 14464 21833 14467
rect 21416 14436 21833 14464
rect 21416 14424 21422 14436
rect 21821 14433 21833 14436
rect 21867 14433 21879 14467
rect 21821 14427 21879 14433
rect 21910 14424 21916 14476
rect 21968 14424 21974 14476
rect 22005 14467 22063 14473
rect 22005 14433 22017 14467
rect 22051 14464 22063 14467
rect 22094 14464 22100 14476
rect 22051 14436 22100 14464
rect 22051 14433 22063 14436
rect 22005 14427 22063 14433
rect 22094 14424 22100 14436
rect 22152 14424 22158 14476
rect 22189 14467 22247 14473
rect 22189 14433 22201 14467
rect 22235 14433 22247 14467
rect 22189 14427 22247 14433
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20640 14368 21097 14396
rect 20533 14359 20591 14365
rect 21085 14365 21097 14368
rect 21131 14396 21143 14399
rect 21545 14399 21603 14405
rect 21545 14396 21557 14399
rect 21131 14368 21557 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 21545 14365 21557 14368
rect 21591 14396 21603 14399
rect 22204 14396 22232 14427
rect 22278 14424 22284 14476
rect 22336 14464 22342 14476
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 22336 14436 22385 14464
rect 22336 14424 22342 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 22462 14424 22468 14476
rect 22520 14424 22526 14476
rect 22646 14424 22652 14476
rect 22704 14424 22710 14476
rect 23032 14473 23060 14504
rect 23845 14501 23857 14504
rect 23891 14501 23903 14535
rect 23952 14532 23980 14572
rect 24026 14560 24032 14612
rect 24084 14600 24090 14612
rect 24213 14603 24271 14609
rect 24213 14600 24225 14603
rect 24084 14572 24225 14600
rect 24084 14560 24090 14572
rect 24213 14569 24225 14572
rect 24259 14569 24271 14603
rect 26237 14603 26295 14609
rect 26237 14600 26249 14603
rect 24213 14563 24271 14569
rect 25056 14572 26249 14600
rect 25056 14532 25084 14572
rect 26237 14569 26249 14572
rect 26283 14600 26295 14603
rect 26694 14600 26700 14612
rect 26283 14572 26700 14600
rect 26283 14569 26295 14572
rect 26237 14563 26295 14569
rect 26694 14560 26700 14572
rect 26752 14600 26758 14612
rect 26881 14603 26939 14609
rect 26881 14600 26893 14603
rect 26752 14572 26893 14600
rect 26752 14560 26758 14572
rect 26881 14569 26893 14572
rect 26927 14569 26939 14603
rect 26881 14563 26939 14569
rect 27341 14603 27399 14609
rect 27341 14569 27353 14603
rect 27387 14600 27399 14603
rect 27522 14600 27528 14612
rect 27387 14572 27528 14600
rect 27387 14569 27399 14572
rect 27341 14563 27399 14569
rect 27522 14560 27528 14572
rect 27580 14560 27586 14612
rect 28902 14560 28908 14612
rect 28960 14600 28966 14612
rect 29457 14603 29515 14609
rect 29457 14600 29469 14603
rect 28960 14572 29469 14600
rect 28960 14560 28966 14572
rect 29457 14569 29469 14572
rect 29503 14569 29515 14603
rect 29457 14563 29515 14569
rect 29546 14560 29552 14612
rect 29604 14560 29610 14612
rect 29917 14603 29975 14609
rect 29917 14569 29929 14603
rect 29963 14600 29975 14603
rect 29963 14572 31064 14600
rect 29963 14569 29975 14572
rect 29917 14563 29975 14569
rect 23952 14504 25084 14532
rect 25124 14535 25182 14541
rect 23845 14495 23903 14501
rect 25124 14501 25136 14535
rect 25170 14532 25182 14535
rect 25314 14532 25320 14544
rect 25170 14504 25320 14532
rect 25170 14501 25182 14504
rect 25124 14495 25182 14501
rect 25314 14492 25320 14504
rect 25372 14492 25378 14544
rect 29555 14532 29583 14560
rect 27540 14504 29583 14532
rect 23017 14467 23075 14473
rect 23017 14433 23029 14467
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 23109 14467 23167 14473
rect 23109 14433 23121 14467
rect 23155 14433 23167 14467
rect 23109 14427 23167 14433
rect 23201 14467 23259 14473
rect 23201 14433 23213 14467
rect 23247 14464 23259 14467
rect 23290 14464 23296 14476
rect 23247 14436 23296 14464
rect 23247 14433 23259 14436
rect 23201 14427 23259 14433
rect 21591 14368 22232 14396
rect 23124 14396 23152 14427
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 23382 14424 23388 14476
rect 23440 14424 23446 14476
rect 24118 14464 24124 14476
rect 23492 14436 24124 14464
rect 23492 14396 23520 14436
rect 24118 14424 24124 14436
rect 24176 14424 24182 14476
rect 24302 14424 24308 14476
rect 24360 14464 24366 14476
rect 24397 14467 24455 14473
rect 24397 14464 24409 14467
rect 24360 14436 24409 14464
rect 24360 14424 24366 14436
rect 24397 14433 24409 14436
rect 24443 14433 24455 14467
rect 24762 14464 24768 14476
rect 24397 14427 24455 14433
rect 24596 14436 24768 14464
rect 23124 14368 23520 14396
rect 23661 14399 23719 14405
rect 21591 14365 21603 14368
rect 21545 14359 21603 14365
rect 23661 14365 23673 14399
rect 23707 14396 23719 14399
rect 24596 14396 24624 14436
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 24854 14424 24860 14476
rect 24912 14424 24918 14476
rect 27540 14473 27568 14504
rect 29638 14492 29644 14544
rect 29696 14532 29702 14544
rect 29696 14504 30788 14532
rect 29696 14492 29702 14504
rect 26973 14467 27031 14473
rect 26973 14433 26985 14467
rect 27019 14464 27031 14467
rect 27525 14467 27583 14473
rect 27525 14464 27537 14467
rect 27019 14436 27537 14464
rect 27019 14433 27031 14436
rect 26973 14427 27031 14433
rect 27525 14433 27537 14436
rect 27571 14433 27583 14467
rect 27525 14427 27583 14433
rect 27709 14467 27767 14473
rect 27709 14433 27721 14467
rect 27755 14433 27767 14467
rect 27709 14427 27767 14433
rect 23707 14368 24624 14396
rect 23707 14365 23719 14368
rect 23661 14359 23719 14365
rect 15212 14300 16712 14328
rect 16945 14331 17003 14337
rect 16945 14297 16957 14331
rect 16991 14328 17003 14331
rect 17402 14328 17408 14340
rect 16991 14300 17408 14328
rect 16991 14297 17003 14300
rect 16945 14291 17003 14297
rect 17402 14288 17408 14300
rect 17460 14328 17466 14340
rect 20548 14328 20576 14359
rect 26142 14356 26148 14408
rect 26200 14396 26206 14408
rect 27065 14399 27123 14405
rect 27065 14396 27077 14399
rect 26200 14368 27077 14396
rect 26200 14356 26206 14368
rect 27065 14365 27077 14368
rect 27111 14365 27123 14399
rect 27065 14359 27123 14365
rect 27430 14356 27436 14408
rect 27488 14396 27494 14408
rect 27724 14396 27752 14427
rect 27982 14424 27988 14476
rect 28040 14424 28046 14476
rect 28169 14467 28227 14473
rect 28169 14464 28181 14467
rect 28092 14436 28181 14464
rect 27488 14368 27752 14396
rect 27488 14356 27494 14368
rect 21910 14328 21916 14340
rect 17460 14300 21916 14328
rect 17460 14288 17466 14300
rect 21910 14288 21916 14300
rect 21968 14288 21974 14340
rect 26786 14288 26792 14340
rect 26844 14328 26850 14340
rect 28092 14328 28120 14436
rect 28169 14433 28181 14436
rect 28215 14433 28227 14467
rect 28169 14427 28227 14433
rect 28353 14467 28411 14473
rect 28353 14433 28365 14467
rect 28399 14433 28411 14467
rect 28353 14427 28411 14433
rect 26844 14300 28120 14328
rect 28368 14328 28396 14427
rect 28442 14424 28448 14476
rect 28500 14424 28506 14476
rect 28537 14467 28595 14473
rect 28537 14433 28549 14467
rect 28583 14464 28595 14467
rect 29178 14464 29184 14476
rect 28583 14436 29184 14464
rect 28583 14433 28595 14436
rect 28537 14427 28595 14433
rect 29178 14424 29184 14436
rect 29236 14424 29242 14476
rect 29822 14424 29828 14476
rect 29880 14464 29886 14476
rect 30193 14467 30251 14473
rect 30193 14464 30205 14467
rect 29880 14436 30205 14464
rect 29880 14424 29886 14436
rect 30193 14433 30205 14436
rect 30239 14433 30251 14467
rect 30193 14427 30251 14433
rect 30282 14424 30288 14476
rect 30340 14424 30346 14476
rect 30466 14424 30472 14476
rect 30524 14424 30530 14476
rect 30558 14424 30564 14476
rect 30616 14464 30622 14476
rect 30760 14473 30788 14504
rect 30653 14467 30711 14473
rect 30653 14464 30665 14467
rect 30616 14436 30665 14464
rect 30616 14424 30622 14436
rect 30653 14433 30665 14436
rect 30699 14433 30711 14467
rect 30653 14427 30711 14433
rect 30745 14467 30803 14473
rect 30745 14433 30757 14467
rect 30791 14433 30803 14467
rect 30745 14427 30803 14433
rect 30926 14424 30932 14476
rect 30984 14424 30990 14476
rect 31036 14473 31064 14572
rect 31021 14467 31079 14473
rect 31021 14433 31033 14467
rect 31067 14433 31079 14467
rect 31021 14427 31079 14433
rect 29270 14356 29276 14408
rect 29328 14356 29334 14408
rect 31205 14331 31263 14337
rect 31205 14328 31217 14331
rect 28368 14300 31217 14328
rect 26844 14288 26850 14300
rect 5074 14220 5080 14272
rect 5132 14220 5138 14272
rect 5902 14220 5908 14272
rect 5960 14220 5966 14272
rect 10962 14220 10968 14272
rect 11020 14220 11026 14272
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 17092 14232 17325 14260
rect 17092 14220 17098 14232
rect 17313 14229 17325 14232
rect 17359 14260 17371 14263
rect 17681 14263 17739 14269
rect 17681 14260 17693 14263
rect 17359 14232 17693 14260
rect 17359 14229 17371 14232
rect 17313 14223 17371 14229
rect 17681 14229 17693 14232
rect 17727 14260 17739 14263
rect 18598 14260 18604 14272
rect 17727 14232 18604 14260
rect 17727 14229 17739 14232
rect 17681 14223 17739 14229
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 20438 14220 20444 14272
rect 20496 14260 20502 14272
rect 20898 14260 20904 14272
rect 20496 14232 20904 14260
rect 20496 14220 20502 14232
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 21266 14220 21272 14272
rect 21324 14220 21330 14272
rect 21726 14220 21732 14272
rect 21784 14220 21790 14272
rect 24673 14263 24731 14269
rect 24673 14229 24685 14263
rect 24719 14260 24731 14263
rect 24854 14260 24860 14272
rect 24719 14232 24860 14260
rect 24719 14229 24731 14232
rect 24673 14223 24731 14229
rect 24854 14220 24860 14232
rect 24912 14260 24918 14272
rect 26142 14260 26148 14272
rect 24912 14232 26148 14260
rect 24912 14220 24918 14232
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 26513 14263 26571 14269
rect 26513 14229 26525 14263
rect 26559 14260 26571 14263
rect 26694 14260 26700 14272
rect 26559 14232 26700 14260
rect 26559 14229 26571 14232
rect 26513 14223 26571 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 27893 14263 27951 14269
rect 27893 14229 27905 14263
rect 27939 14260 27951 14263
rect 27982 14260 27988 14272
rect 27939 14232 27988 14260
rect 27939 14229 27951 14232
rect 27893 14223 27951 14229
rect 27982 14220 27988 14232
rect 28040 14220 28046 14272
rect 28092 14260 28120 14300
rect 31205 14297 31217 14300
rect 31251 14297 31263 14331
rect 31205 14291 31263 14297
rect 28626 14260 28632 14272
rect 28092 14232 28632 14260
rect 28626 14220 28632 14232
rect 28684 14220 28690 14272
rect 28813 14263 28871 14269
rect 28813 14229 28825 14263
rect 28859 14260 28871 14263
rect 28994 14260 29000 14272
rect 28859 14232 29000 14260
rect 28859 14229 28871 14232
rect 28813 14223 28871 14229
rect 28994 14220 29000 14232
rect 29052 14220 29058 14272
rect 29086 14220 29092 14272
rect 29144 14260 29150 14272
rect 30009 14263 30067 14269
rect 30009 14260 30021 14263
rect 29144 14232 30021 14260
rect 29144 14220 29150 14232
rect 30009 14229 30021 14232
rect 30055 14229 30067 14263
rect 30009 14223 30067 14229
rect 552 14170 31648 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 11436 14170
rect 11488 14118 11500 14170
rect 11552 14118 11564 14170
rect 11616 14118 11628 14170
rect 11680 14118 11692 14170
rect 11744 14118 19210 14170
rect 19262 14118 19274 14170
rect 19326 14118 19338 14170
rect 19390 14118 19402 14170
rect 19454 14118 19466 14170
rect 19518 14118 26984 14170
rect 27036 14118 27048 14170
rect 27100 14118 27112 14170
rect 27164 14118 27176 14170
rect 27228 14118 27240 14170
rect 27292 14118 31648 14170
rect 552 14096 31648 14118
rect 6270 14056 6276 14068
rect 4356 14028 6276 14056
rect 3050 13948 3056 14000
rect 3108 13948 3114 14000
rect 3068 13920 3096 13948
rect 4062 13920 4068 13932
rect 3068 13892 4068 13920
rect 4062 13880 4068 13892
rect 4120 13920 4126 13932
rect 4120 13892 4200 13920
rect 4120 13880 4126 13892
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 1360 13824 2605 13852
rect 1360 13812 1366 13824
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 2608 13784 2636 13815
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 3053 13855 3111 13861
rect 3053 13821 3065 13855
rect 3099 13852 3111 13855
rect 3697 13855 3755 13861
rect 3697 13852 3709 13855
rect 3099 13824 3709 13852
rect 3099 13821 3111 13824
rect 3053 13815 3111 13821
rect 3697 13821 3709 13824
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 3878 13812 3884 13864
rect 3936 13812 3942 13864
rect 4172 13861 4200 13892
rect 4356 13861 4384 14028
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 7009 14059 7067 14065
rect 7009 14056 7021 14059
rect 6420 14028 7021 14056
rect 6420 14016 6426 14028
rect 7009 14025 7021 14028
rect 7055 14025 7067 14059
rect 7009 14019 7067 14025
rect 5534 13988 5540 14000
rect 4724 13960 5540 13988
rect 4724 13861 4752 13960
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 7024 13988 7052 14019
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 9548 14028 9965 14056
rect 9548 14016 9554 14028
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 9953 14019 10011 14025
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 12526 14056 12532 14068
rect 10652 14028 12532 14056
rect 10652 14016 10658 14028
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 13909 14059 13967 14065
rect 13909 14056 13921 14059
rect 13780 14028 13921 14056
rect 13780 14016 13786 14028
rect 13909 14025 13921 14028
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 15010 14016 15016 14068
rect 15068 14016 15074 14068
rect 15197 14059 15255 14065
rect 15197 14025 15209 14059
rect 15243 14025 15255 14059
rect 15197 14019 15255 14025
rect 11238 13988 11244 14000
rect 7024 13960 11244 13988
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 14918 13948 14924 14000
rect 14976 13988 14982 14000
rect 15212 13988 15240 14019
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 16356 14028 18000 14056
rect 16356 14016 16362 14028
rect 16482 13988 16488 14000
rect 14976 13960 16488 13988
rect 14976 13948 14982 13960
rect 16482 13948 16488 13960
rect 16540 13948 16546 14000
rect 17494 13948 17500 14000
rect 17552 13948 17558 14000
rect 17589 13991 17647 13997
rect 17589 13957 17601 13991
rect 17635 13988 17647 13991
rect 17862 13988 17868 14000
rect 17635 13960 17868 13988
rect 17635 13957 17647 13960
rect 17589 13951 17647 13957
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 17972 13988 18000 14028
rect 18138 14016 18144 14068
rect 18196 14016 18202 14068
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 21266 14056 21272 14068
rect 20119 14028 21272 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 22462 14056 22468 14068
rect 21376 14028 22468 14056
rect 17972 13960 19840 13988
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13920 4859 13923
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 4847 13892 5641 13920
rect 4847 13889 4859 13892
rect 4801 13883 4859 13889
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7156 13892 7757 13920
rect 7156 13880 7162 13892
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 9490 13920 9496 13932
rect 7745 13883 7803 13889
rect 8036 13892 9496 13920
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13821 4399 13855
rect 4341 13815 4399 13821
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13821 4767 13855
rect 4709 13815 4767 13821
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5199 13855 5257 13861
rect 5199 13852 5211 13855
rect 5132 13824 5211 13852
rect 5132 13812 5138 13824
rect 5199 13821 5211 13824
rect 5245 13821 5257 13855
rect 5199 13815 5257 13821
rect 5350 13812 5356 13864
rect 5408 13812 5414 13864
rect 5902 13861 5908 13864
rect 5896 13852 5908 13861
rect 5863 13824 5908 13852
rect 5896 13815 5908 13824
rect 5902 13812 5908 13815
rect 5960 13812 5966 13864
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 8036 13852 8064 13892
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 10962 13920 10968 13932
rect 10152 13892 10968 13920
rect 6328 13824 8064 13852
rect 6328 13812 6334 13824
rect 8938 13812 8944 13864
rect 8996 13852 9002 13864
rect 9306 13852 9312 13864
rect 8996 13824 9312 13852
rect 8996 13812 9002 13824
rect 9306 13812 9312 13824
rect 9364 13852 9370 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 9364 13824 9689 13852
rect 9364 13812 9370 13824
rect 9677 13821 9689 13824
rect 9723 13852 9735 13855
rect 9950 13852 9956 13864
rect 9723 13824 9956 13852
rect 9723 13821 9735 13824
rect 9677 13815 9735 13821
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10152 13861 10180 13892
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 14642 13880 14648 13932
rect 14700 13920 14706 13932
rect 15381 13923 15439 13929
rect 14700 13892 15332 13920
rect 14700 13880 14706 13892
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 10594 13852 10600 13864
rect 10367 13824 10600 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10735 13824 11100 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 5442 13784 5448 13796
rect 2608 13756 5448 13784
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 6788 13756 7573 13784
rect 6788 13744 6794 13756
rect 7561 13753 7573 13756
rect 7607 13753 7619 13787
rect 7561 13747 7619 13753
rect 9490 13744 9496 13796
rect 9548 13744 9554 13796
rect 9861 13787 9919 13793
rect 9861 13753 9873 13787
rect 9907 13784 9919 13787
rect 10042 13784 10048 13796
rect 9907 13756 10048 13784
rect 9907 13753 9919 13756
rect 9861 13747 9919 13753
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 11072 13784 11100 13824
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 11204 13824 11253 13852
rect 11204 13812 11210 13824
rect 11241 13821 11253 13824
rect 11287 13852 11299 13855
rect 11974 13852 11980 13864
rect 11287 13824 11980 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 11974 13812 11980 13824
rect 12032 13852 12038 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 12032 13824 14013 13852
rect 12032 13812 12038 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 14792 13824 15209 13852
rect 14792 13812 14798 13824
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15304 13852 15332 13892
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 15427 13892 16405 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 16393 13889 16405 13892
rect 16439 13920 16451 13923
rect 17770 13920 17776 13932
rect 16439 13892 17776 13920
rect 16439 13889 16451 13892
rect 16393 13883 16451 13889
rect 17770 13880 17776 13892
rect 17828 13880 17834 13932
rect 19426 13920 19432 13932
rect 17880 13892 19432 13920
rect 16298 13852 16304 13864
rect 15304 13824 16304 13852
rect 15197 13815 15255 13821
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 16540 13824 17540 13852
rect 16540 13812 16546 13824
rect 11882 13784 11888 13796
rect 11072 13756 11888 13784
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 15470 13744 15476 13796
rect 15528 13744 15534 13796
rect 17034 13744 17040 13796
rect 17092 13784 17098 13796
rect 17129 13787 17187 13793
rect 17129 13784 17141 13787
rect 17092 13756 17141 13784
rect 17092 13744 17098 13756
rect 17129 13753 17141 13756
rect 17175 13753 17187 13787
rect 17512 13784 17540 13824
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 17681 13855 17739 13861
rect 17681 13852 17693 13855
rect 17644 13824 17693 13852
rect 17644 13812 17650 13824
rect 17681 13821 17693 13824
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 17880 13796 17908 13892
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 19812 13920 19840 13960
rect 19886 13948 19892 14000
rect 19944 13988 19950 14000
rect 20349 13991 20407 13997
rect 20349 13988 20361 13991
rect 19944 13960 20361 13988
rect 19944 13948 19950 13960
rect 20349 13957 20361 13960
rect 20395 13957 20407 13991
rect 20349 13951 20407 13957
rect 20530 13948 20536 14000
rect 20588 13948 20594 14000
rect 20901 13991 20959 13997
rect 20901 13957 20913 13991
rect 20947 13988 20959 13991
rect 21082 13988 21088 14000
rect 20947 13960 21088 13988
rect 20947 13957 20959 13960
rect 20901 13951 20959 13957
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 21376 13988 21404 14028
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 23750 14016 23756 14068
rect 23808 14056 23814 14068
rect 23808 14028 25184 14056
rect 23808 14016 23814 14028
rect 21192 13960 21404 13988
rect 25156 13988 25184 14028
rect 25222 14016 25228 14068
rect 25280 14056 25286 14068
rect 25682 14056 25688 14068
rect 25280 14028 25688 14056
rect 25280 14016 25286 14028
rect 25682 14016 25688 14028
rect 25740 14016 25746 14068
rect 27985 14059 28043 14065
rect 27985 14056 27997 14059
rect 27080 14028 27997 14056
rect 26786 13988 26792 14000
rect 25156 13960 26792 13988
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 19812 13892 20821 13920
rect 20809 13889 20821 13892
rect 20855 13920 20867 13923
rect 21192 13920 21220 13960
rect 20855 13892 21220 13920
rect 22281 13923 22339 13929
rect 20855 13889 20867 13892
rect 20809 13883 20867 13889
rect 22281 13889 22293 13923
rect 22327 13920 22339 13923
rect 22465 13923 22523 13929
rect 22465 13920 22477 13923
rect 22327 13892 22477 13920
rect 22327 13889 22339 13892
rect 22281 13883 22339 13889
rect 22465 13889 22477 13892
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 23017 13923 23075 13929
rect 23017 13889 23029 13923
rect 23063 13920 23075 13923
rect 23063 13892 23980 13920
rect 23063 13889 23075 13892
rect 23017 13883 23075 13889
rect 18046 13812 18052 13864
rect 18104 13812 18110 13864
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13821 18199 13855
rect 18141 13815 18199 13821
rect 17862 13784 17868 13796
rect 17512 13756 17868 13784
rect 17129 13747 17187 13753
rect 17862 13744 17868 13756
rect 17920 13744 17926 13796
rect 18156 13784 18184 13815
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 22014 13855 22072 13861
rect 22014 13852 22026 13855
rect 20312 13824 22026 13852
rect 20312 13812 20318 13824
rect 22014 13821 22026 13824
rect 22060 13821 22072 13855
rect 22014 13815 22072 13821
rect 22370 13812 22376 13864
rect 22428 13812 22434 13864
rect 23293 13855 23351 13861
rect 23293 13821 23305 13855
rect 23339 13821 23351 13855
rect 23293 13815 23351 13821
rect 18064 13756 18184 13784
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 2501 13719 2559 13725
rect 2501 13716 2513 13719
rect 2372 13688 2513 13716
rect 2372 13676 2378 13688
rect 2501 13685 2513 13688
rect 2547 13685 2559 13719
rect 2501 13679 2559 13685
rect 2958 13676 2964 13728
rect 3016 13676 3022 13728
rect 4985 13719 5043 13725
rect 4985 13685 4997 13719
rect 5031 13716 5043 13719
rect 5166 13716 5172 13728
rect 5031 13688 5172 13716
rect 5031 13685 5043 13688
rect 4985 13679 5043 13685
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 7190 13676 7196 13728
rect 7248 13676 7254 13728
rect 7650 13676 7656 13728
rect 7708 13676 7714 13728
rect 10318 13676 10324 13728
rect 10376 13716 10382 13728
rect 10505 13719 10563 13725
rect 10505 13716 10517 13719
rect 10376 13688 10517 13716
rect 10376 13676 10382 13688
rect 10505 13685 10517 13688
rect 10551 13685 10563 13719
rect 10505 13679 10563 13685
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 11112 13688 11161 13716
rect 11112 13676 11118 13688
rect 11149 13685 11161 13688
rect 11195 13685 11207 13719
rect 11149 13679 11207 13685
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 17310 13716 17316 13728
rect 16816 13688 17316 13716
rect 16816 13676 16822 13688
rect 17310 13676 17316 13688
rect 17368 13716 17374 13728
rect 18064 13716 18092 13756
rect 19610 13744 19616 13796
rect 19668 13784 19674 13796
rect 19889 13787 19947 13793
rect 19889 13784 19901 13787
rect 19668 13756 19901 13784
rect 19668 13744 19674 13756
rect 19889 13753 19901 13756
rect 19935 13784 19947 13787
rect 19978 13784 19984 13796
rect 19935 13756 19984 13784
rect 19935 13753 19947 13756
rect 19889 13747 19947 13753
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 20105 13787 20163 13793
rect 20105 13753 20117 13787
rect 20151 13784 20163 13787
rect 20990 13784 20996 13796
rect 20151 13756 20996 13784
rect 20151 13753 20163 13756
rect 20105 13747 20163 13753
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 23308 13784 23336 13815
rect 23382 13812 23388 13864
rect 23440 13812 23446 13864
rect 23477 13855 23535 13861
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 23566 13852 23572 13864
rect 23523 13824 23572 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 23566 13812 23572 13824
rect 23624 13812 23630 13864
rect 23661 13855 23719 13861
rect 23661 13821 23673 13855
rect 23707 13852 23719 13855
rect 23750 13852 23756 13864
rect 23707 13824 23756 13852
rect 23707 13821 23719 13824
rect 23661 13815 23719 13821
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 23842 13812 23848 13864
rect 23900 13812 23906 13864
rect 23952 13852 23980 13892
rect 25406 13880 25412 13932
rect 25464 13920 25470 13932
rect 25961 13923 26019 13929
rect 25464 13892 25820 13920
rect 25464 13880 25470 13892
rect 24101 13855 24159 13861
rect 24101 13852 24113 13855
rect 23952 13824 24113 13852
rect 24101 13821 24113 13824
rect 24147 13821 24159 13855
rect 24101 13815 24159 13821
rect 25682 13812 25688 13864
rect 25740 13812 25746 13864
rect 25792 13852 25820 13892
rect 25961 13889 25973 13923
rect 26007 13920 26019 13923
rect 26142 13920 26148 13932
rect 26007 13892 26148 13920
rect 26007 13889 26019 13892
rect 25961 13883 26019 13889
rect 26142 13880 26148 13892
rect 26200 13880 26206 13932
rect 26712 13861 26740 13960
rect 26786 13948 26792 13960
rect 26844 13948 26850 14000
rect 26697 13855 26755 13861
rect 25792 13824 26648 13852
rect 24302 13784 24308 13796
rect 23308 13756 24308 13784
rect 24302 13744 24308 13756
rect 24360 13744 24366 13796
rect 26510 13784 26516 13796
rect 24412 13756 26516 13784
rect 17368 13688 18092 13716
rect 17368 13676 17374 13688
rect 18322 13676 18328 13728
rect 18380 13676 18386 13728
rect 20254 13676 20260 13728
rect 20312 13676 20318 13728
rect 20806 13676 20812 13728
rect 20864 13716 20870 13728
rect 24412 13716 24440 13756
rect 26510 13744 26516 13756
rect 26568 13744 26574 13796
rect 26620 13784 26648 13824
rect 26697 13821 26709 13855
rect 26743 13821 26755 13855
rect 26697 13815 26755 13821
rect 26878 13812 26884 13864
rect 26936 13812 26942 13864
rect 26970 13812 26976 13864
rect 27028 13812 27034 13864
rect 27080 13861 27108 14028
rect 27985 14025 27997 14028
rect 28031 14025 28043 14059
rect 27985 14019 28043 14025
rect 28166 14016 28172 14068
rect 28224 14056 28230 14068
rect 28224 14028 29500 14056
rect 28224 14016 28230 14028
rect 29362 13988 29368 14000
rect 27733 13960 29368 13988
rect 27341 13923 27399 13929
rect 27341 13889 27353 13923
rect 27387 13920 27399 13923
rect 27614 13920 27620 13932
rect 27387 13892 27620 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 27614 13880 27620 13892
rect 27672 13880 27678 13932
rect 27065 13855 27123 13861
rect 27065 13821 27077 13855
rect 27111 13821 27123 13855
rect 27065 13815 27123 13821
rect 27430 13784 27436 13796
rect 26620 13756 27436 13784
rect 27430 13744 27436 13756
rect 27488 13784 27494 13796
rect 27733 13793 27761 13960
rect 29362 13948 29368 13960
rect 29420 13948 29426 14000
rect 29472 13988 29500 14028
rect 29822 14016 29828 14068
rect 29880 14016 29886 14068
rect 30466 14016 30472 14068
rect 30524 14056 30530 14068
rect 30561 14059 30619 14065
rect 30561 14056 30573 14059
rect 30524 14028 30573 14056
rect 30524 14016 30530 14028
rect 30561 14025 30573 14028
rect 30607 14025 30619 14059
rect 30561 14019 30619 14025
rect 29472 13960 30236 13988
rect 27893 13923 27951 13929
rect 27893 13889 27905 13923
rect 27939 13920 27951 13923
rect 27939 13892 28948 13920
rect 27939 13889 27951 13892
rect 27893 13883 27951 13889
rect 28537 13855 28595 13861
rect 28537 13821 28549 13855
rect 28583 13821 28595 13855
rect 28920 13852 28948 13892
rect 29270 13880 29276 13932
rect 29328 13880 29334 13932
rect 29917 13855 29975 13861
rect 29917 13852 29929 13855
rect 28920 13824 29929 13852
rect 28537 13815 28595 13821
rect 29917 13821 29929 13824
rect 29963 13821 29975 13855
rect 29917 13815 29975 13821
rect 27525 13787 27583 13793
rect 27525 13784 27537 13787
rect 27488 13756 27537 13784
rect 27488 13744 27494 13756
rect 27525 13753 27537 13756
rect 27571 13753 27583 13787
rect 27525 13747 27583 13753
rect 27709 13787 27767 13793
rect 27709 13753 27721 13787
rect 27755 13753 27767 13787
rect 27709 13747 27767 13753
rect 28552 13784 28580 13815
rect 30098 13812 30104 13864
rect 30156 13812 30162 13864
rect 30208 13861 30236 13960
rect 30193 13855 30251 13861
rect 30193 13821 30205 13855
rect 30239 13821 30251 13855
rect 30193 13815 30251 13821
rect 30285 13855 30343 13861
rect 30285 13821 30297 13855
rect 30331 13821 30343 13855
rect 30285 13815 30343 13821
rect 29457 13787 29515 13793
rect 29457 13784 29469 13787
rect 28552 13756 29469 13784
rect 20864 13688 24440 13716
rect 20864 13676 20870 13688
rect 25314 13676 25320 13728
rect 25372 13676 25378 13728
rect 25777 13719 25835 13725
rect 25777 13685 25789 13719
rect 25823 13716 25835 13719
rect 25866 13716 25872 13728
rect 25823 13688 25872 13716
rect 25823 13685 25835 13688
rect 25777 13679 25835 13685
rect 25866 13676 25872 13688
rect 25924 13716 25930 13728
rect 28552 13716 28580 13756
rect 29457 13753 29469 13756
rect 29503 13784 29515 13787
rect 30300 13784 30328 13815
rect 29503 13756 30328 13784
rect 29503 13753 29515 13756
rect 29457 13747 29515 13753
rect 28718 13716 28724 13728
rect 25924 13688 28724 13716
rect 25924 13676 25930 13688
rect 28718 13676 28724 13688
rect 28776 13676 28782 13728
rect 29362 13676 29368 13728
rect 29420 13716 29426 13728
rect 30742 13716 30748 13728
rect 29420 13688 30748 13716
rect 29420 13676 29426 13688
rect 30742 13676 30748 13688
rect 30800 13676 30806 13728
rect 552 13626 31648 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 12096 13626
rect 12148 13574 12160 13626
rect 12212 13574 12224 13626
rect 12276 13574 12288 13626
rect 12340 13574 12352 13626
rect 12404 13574 19870 13626
rect 19922 13574 19934 13626
rect 19986 13574 19998 13626
rect 20050 13574 20062 13626
rect 20114 13574 20126 13626
rect 20178 13574 27644 13626
rect 27696 13574 27708 13626
rect 27760 13574 27772 13626
rect 27824 13574 27836 13626
rect 27888 13574 27900 13626
rect 27952 13574 31648 13626
rect 552 13552 31648 13574
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3510 13512 3516 13524
rect 2924 13484 3516 13512
rect 2924 13472 2930 13484
rect 3510 13472 3516 13484
rect 3568 13512 3574 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3568 13484 3801 13512
rect 3568 13472 3574 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 4065 13515 4123 13521
rect 4065 13481 4077 13515
rect 4111 13512 4123 13515
rect 4890 13512 4896 13524
rect 4111 13484 4896 13512
rect 4111 13481 4123 13484
rect 4065 13475 4123 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 7469 13515 7527 13521
rect 7469 13481 7481 13515
rect 7515 13512 7527 13515
rect 7650 13512 7656 13524
rect 7515 13484 7656 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 7760 13484 9674 13512
rect 2584 13447 2642 13453
rect 2584 13413 2596 13447
rect 2630 13444 2642 13447
rect 2958 13444 2964 13456
rect 2630 13416 2964 13444
rect 2630 13413 2642 13416
rect 2584 13407 2642 13413
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 3602 13404 3608 13456
rect 3660 13444 3666 13456
rect 3973 13447 4031 13453
rect 3973 13444 3985 13447
rect 3660 13416 3985 13444
rect 3660 13404 3666 13416
rect 3973 13413 3985 13416
rect 4019 13413 4031 13447
rect 4341 13447 4399 13453
rect 4341 13444 4353 13447
rect 3973 13407 4031 13413
rect 4080 13416 4353 13444
rect 2314 13336 2320 13388
rect 2372 13336 2378 13388
rect 3418 13336 3424 13388
rect 3476 13376 3482 13388
rect 4080 13376 4108 13416
rect 4341 13413 4353 13416
rect 4387 13413 4399 13447
rect 4908 13444 4936 13472
rect 7760 13444 7788 13484
rect 4908 13416 7788 13444
rect 4341 13407 4399 13413
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 9646 13444 9674 13484
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12345 13515 12403 13521
rect 12345 13512 12357 13515
rect 11940 13484 12357 13512
rect 11940 13472 11946 13484
rect 12345 13481 12357 13484
rect 12391 13481 12403 13515
rect 12345 13475 12403 13481
rect 12894 13472 12900 13524
rect 12952 13472 12958 13524
rect 13630 13472 13636 13524
rect 13688 13472 13694 13524
rect 14461 13515 14519 13521
rect 14461 13481 14473 13515
rect 14507 13512 14519 13515
rect 16666 13512 16672 13524
rect 14507 13484 16672 13512
rect 14507 13481 14519 13484
rect 14461 13475 14519 13481
rect 10597 13447 10655 13453
rect 8260 13416 8340 13444
rect 9646 13416 10272 13444
rect 8260 13404 8266 13416
rect 3476 13348 4108 13376
rect 4157 13379 4215 13385
rect 3476 13336 3482 13348
rect 4157 13345 4169 13379
rect 4203 13345 4215 13379
rect 4157 13339 4215 13345
rect 3878 13308 3884 13320
rect 3712 13280 3884 13308
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 3712 13181 3740 13280
rect 3878 13268 3884 13280
rect 3936 13308 3942 13320
rect 4172 13308 4200 13339
rect 5442 13336 5448 13388
rect 5500 13336 5506 13388
rect 6080 13379 6138 13385
rect 6080 13345 6092 13379
rect 6126 13376 6138 13379
rect 7190 13376 7196 13388
rect 6126 13348 7196 13376
rect 6126 13345 6138 13348
rect 6080 13339 6138 13345
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 8312 13383 8340 13416
rect 8297 13377 8355 13383
rect 8297 13343 8309 13377
rect 8343 13343 8355 13377
rect 8297 13337 8355 13343
rect 9306 13336 9312 13388
rect 9364 13336 9370 13388
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 3936 13280 4200 13308
rect 5537 13311 5595 13317
rect 3936 13268 3942 13280
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5583 13280 5825 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 8021 13311 8079 13317
rect 8021 13308 8033 13311
rect 5813 13271 5871 13277
rect 7024 13280 8033 13308
rect 3697 13175 3755 13181
rect 3697 13172 3709 13175
rect 3476 13144 3709 13172
rect 3476 13132 3482 13144
rect 3697 13141 3709 13144
rect 3743 13141 3755 13175
rect 7024 13172 7052 13280
rect 8021 13277 8033 13280
rect 8067 13308 8079 13311
rect 9398 13308 9404 13320
rect 8067 13280 9404 13308
rect 8067 13277 8079 13280
rect 8021 13271 8079 13277
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 9508 13240 9536 13339
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9732 13348 9965 13376
rect 9732 13336 9738 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 10042 13336 10048 13388
rect 10100 13376 10106 13388
rect 10244 13385 10272 13416
rect 10597 13413 10609 13447
rect 10643 13444 10655 13447
rect 11210 13447 11268 13453
rect 11210 13444 11222 13447
rect 10643 13416 11222 13444
rect 10643 13413 10655 13416
rect 10597 13407 10655 13413
rect 11210 13413 11222 13416
rect 11256 13413 11268 13447
rect 11210 13407 11268 13413
rect 13173 13447 13231 13453
rect 13173 13413 13185 13447
rect 13219 13444 13231 13447
rect 13648 13444 13676 13472
rect 13219 13416 13676 13444
rect 13219 13413 13231 13416
rect 13173 13407 13231 13413
rect 13722 13404 13728 13456
rect 13780 13444 13786 13456
rect 14476 13444 14504 13475
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 20438 13512 20444 13524
rect 18187 13484 20444 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 23842 13472 23848 13524
rect 23900 13512 23906 13524
rect 24121 13515 24179 13521
rect 24121 13512 24133 13515
rect 23900 13484 24133 13512
rect 23900 13472 23906 13484
rect 24121 13481 24133 13484
rect 24167 13481 24179 13515
rect 24121 13475 24179 13481
rect 28718 13472 28724 13524
rect 28776 13472 28782 13524
rect 29178 13472 29184 13524
rect 29236 13512 29242 13524
rect 29733 13515 29791 13521
rect 29733 13512 29745 13515
rect 29236 13484 29745 13512
rect 29236 13472 29242 13484
rect 29733 13481 29745 13484
rect 29779 13481 29791 13515
rect 29733 13475 29791 13481
rect 14734 13444 14740 13456
rect 13780 13416 14504 13444
rect 14568 13416 14740 13444
rect 13780 13404 13786 13416
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 10100 13348 10149 13376
rect 10100 13336 10106 13348
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 7156 13212 9536 13240
rect 7156 13200 7162 13212
rect 7193 13175 7251 13181
rect 7193 13172 7205 13175
rect 7024 13144 7205 13172
rect 3697 13135 3755 13141
rect 7193 13141 7205 13144
rect 7239 13141 7251 13175
rect 7193 13135 7251 13141
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 8389 13175 8447 13181
rect 8389 13172 8401 13175
rect 8352 13144 8401 13172
rect 8352 13132 8358 13144
rect 8389 13141 8401 13144
rect 8435 13141 8447 13175
rect 8389 13135 8447 13141
rect 8846 13132 8852 13184
rect 8904 13172 8910 13184
rect 9125 13175 9183 13181
rect 9125 13172 9137 13175
rect 8904 13144 9137 13172
rect 8904 13132 8910 13144
rect 9125 13141 9137 13144
rect 9171 13141 9183 13175
rect 10244 13172 10272 13339
rect 10318 13336 10324 13388
rect 10376 13336 10382 13388
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 11054 13376 11060 13388
rect 11011 13348 11060 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 11848 13348 12725 13376
rect 11848 13336 11854 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 13354 13336 13360 13388
rect 13412 13336 13418 13388
rect 13446 13336 13452 13388
rect 13504 13376 13510 13388
rect 14016 13385 14044 13416
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13504 13348 13645 13376
rect 13504 13336 13510 13348
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13345 13875 13379
rect 13817 13339 13875 13345
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13345 13967 13379
rect 13909 13339 13967 13345
rect 14001 13379 14059 13385
rect 14001 13345 14013 13379
rect 14047 13345 14059 13379
rect 14568 13376 14596 13416
rect 14734 13404 14740 13416
rect 14792 13444 14798 13456
rect 14792 13416 15240 13444
rect 14792 13404 14798 13416
rect 15212 13385 15240 13416
rect 24302 13404 24308 13456
rect 24360 13404 24366 13456
rect 25038 13404 25044 13456
rect 25096 13404 25102 13456
rect 25406 13404 25412 13456
rect 25464 13444 25470 13456
rect 25685 13447 25743 13453
rect 25685 13444 25697 13447
rect 25464 13416 25697 13444
rect 25464 13404 25470 13416
rect 25685 13413 25697 13416
rect 25731 13413 25743 13447
rect 25685 13407 25743 13413
rect 25866 13404 25872 13456
rect 25924 13404 25930 13456
rect 26050 13404 26056 13456
rect 26108 13404 26114 13456
rect 26694 13404 26700 13456
rect 26752 13444 26758 13456
rect 26752 13416 26924 13444
rect 26752 13404 26758 13416
rect 14001 13339 14059 13345
rect 14200 13348 14596 13376
rect 14645 13379 14703 13385
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 12584 13280 13093 13308
rect 12584 13268 12590 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 13832 13308 13860 13339
rect 13587 13280 13860 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 13170 13240 13176 13252
rect 12636 13212 13176 13240
rect 12636 13172 12664 13212
rect 13170 13200 13176 13212
rect 13228 13240 13234 13252
rect 13924 13240 13952 13339
rect 13228 13212 13952 13240
rect 13228 13200 13234 13212
rect 10244 13144 12664 13172
rect 9125 13135 9183 13141
rect 12710 13132 12716 13184
rect 12768 13132 12774 13184
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 14200 13172 14228 13348
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13345 15255 13379
rect 15197 13339 15255 13345
rect 14660 13308 14688 13339
rect 15378 13336 15384 13388
rect 15436 13336 15442 13388
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13376 16727 13379
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 16715 13348 17049 13376
rect 16715 13345 16727 13348
rect 16669 13339 16727 13345
rect 17037 13345 17049 13348
rect 17083 13376 17095 13379
rect 17126 13376 17132 13388
rect 17083 13348 17132 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13376 17739 13379
rect 17954 13376 17960 13388
rect 17727 13348 17960 13376
rect 17727 13345 17739 13348
rect 17681 13339 17739 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 18601 13379 18659 13385
rect 18601 13345 18613 13379
rect 18647 13376 18659 13379
rect 19610 13376 19616 13388
rect 18647 13348 19616 13376
rect 18647 13345 18659 13348
rect 18601 13339 18659 13345
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 21453 13379 21511 13385
rect 21453 13345 21465 13379
rect 21499 13376 21511 13379
rect 21910 13376 21916 13388
rect 21499 13348 21916 13376
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22186 13336 22192 13388
rect 22244 13376 22250 13388
rect 23937 13379 23995 13385
rect 23937 13376 23949 13379
rect 22244 13348 23949 13376
rect 22244 13336 22250 13348
rect 23937 13345 23949 13348
rect 23983 13345 23995 13379
rect 23937 13339 23995 13345
rect 24213 13379 24271 13385
rect 24213 13345 24225 13379
rect 24259 13376 24271 13379
rect 24578 13376 24584 13388
rect 24259 13348 24584 13376
rect 24259 13345 24271 13348
rect 24213 13339 24271 13345
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 24949 13379 25007 13385
rect 24949 13345 24961 13379
rect 24995 13376 25007 13379
rect 25130 13376 25136 13388
rect 24995 13348 25136 13376
rect 24995 13345 25007 13348
rect 24949 13339 25007 13345
rect 25130 13336 25136 13348
rect 25188 13336 25194 13388
rect 25222 13336 25228 13388
rect 25280 13336 25286 13388
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13345 25375 13379
rect 25317 13339 25375 13345
rect 16482 13308 16488 13320
rect 14660 13280 16488 13308
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 18230 13308 18236 13320
rect 17819 13280 18236 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19058 13308 19064 13320
rect 18923 13280 19064 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19702 13268 19708 13320
rect 19760 13308 19766 13320
rect 20530 13308 20536 13320
rect 19760 13280 20536 13308
rect 19760 13268 19766 13280
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 21821 13311 21879 13317
rect 21821 13277 21833 13311
rect 21867 13308 21879 13311
rect 22554 13308 22560 13320
rect 21867 13280 22560 13308
rect 21867 13277 21879 13280
rect 21821 13271 21879 13277
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 25332 13308 25360 13339
rect 25498 13336 25504 13388
rect 25556 13336 25562 13388
rect 25590 13336 25596 13388
rect 25648 13336 25654 13388
rect 26418 13336 26424 13388
rect 26476 13376 26482 13388
rect 26513 13379 26571 13385
rect 26513 13376 26525 13379
rect 26476 13348 26525 13376
rect 26476 13336 26482 13348
rect 26513 13345 26525 13348
rect 26559 13345 26571 13379
rect 26513 13339 26571 13345
rect 26602 13336 26608 13388
rect 26660 13336 26666 13388
rect 26896 13385 26924 13416
rect 26970 13404 26976 13456
rect 27028 13444 27034 13456
rect 27065 13447 27123 13453
rect 27065 13444 27077 13447
rect 27028 13416 27077 13444
rect 27028 13404 27034 13416
rect 27065 13413 27077 13416
rect 27111 13413 27123 13447
rect 27982 13444 27988 13456
rect 27065 13407 27123 13413
rect 27356 13416 27988 13444
rect 27356 13385 27384 13416
rect 27982 13404 27988 13416
rect 28040 13404 28046 13456
rect 28166 13404 28172 13456
rect 28224 13444 28230 13456
rect 28224 13416 29224 13444
rect 28224 13404 28230 13416
rect 27614 13385 27620 13388
rect 26789 13379 26847 13385
rect 26789 13345 26801 13379
rect 26835 13345 26847 13379
rect 26789 13339 26847 13345
rect 26881 13379 26939 13385
rect 26881 13345 26893 13379
rect 26927 13345 26939 13379
rect 26881 13339 26939 13345
rect 27341 13379 27399 13385
rect 27341 13345 27353 13379
rect 27387 13345 27399 13379
rect 27608 13376 27620 13385
rect 27575 13348 27620 13376
rect 27341 13339 27399 13345
rect 27608 13339 27620 13348
rect 26804 13308 26832 13339
rect 27614 13336 27620 13339
rect 27672 13336 27678 13388
rect 28626 13336 28632 13388
rect 28684 13376 28690 13388
rect 28905 13379 28963 13385
rect 28905 13376 28917 13379
rect 28684 13348 28917 13376
rect 28684 13336 28690 13348
rect 28905 13345 28917 13348
rect 28951 13345 28963 13379
rect 28905 13339 28963 13345
rect 29086 13336 29092 13388
rect 29144 13336 29150 13388
rect 29196 13385 29224 13416
rect 29181 13379 29239 13385
rect 29181 13345 29193 13379
rect 29227 13345 29239 13379
rect 29181 13339 29239 13345
rect 29273 13379 29331 13385
rect 29273 13345 29285 13379
rect 29319 13376 29331 13379
rect 30469 13379 30527 13385
rect 30469 13376 30481 13379
rect 29319 13348 30481 13376
rect 29319 13345 29331 13348
rect 29273 13339 29331 13345
rect 30469 13345 30481 13348
rect 30515 13345 30527 13379
rect 30469 13339 30527 13345
rect 24228 13280 26832 13308
rect 30377 13311 30435 13317
rect 18325 13243 18383 13249
rect 18325 13209 18337 13243
rect 18371 13240 18383 13243
rect 18785 13243 18843 13249
rect 18785 13240 18797 13243
rect 18371 13212 18797 13240
rect 18371 13209 18383 13212
rect 18325 13203 18383 13209
rect 18785 13209 18797 13212
rect 18831 13209 18843 13243
rect 21744 13240 21772 13268
rect 24228 13252 24256 13280
rect 30377 13277 30389 13311
rect 30423 13308 30435 13311
rect 30742 13308 30748 13320
rect 30423 13280 30748 13308
rect 30423 13277 30435 13280
rect 30377 13271 30435 13277
rect 30742 13268 30748 13280
rect 30800 13268 30806 13320
rect 31018 13268 31024 13320
rect 31076 13268 31082 13320
rect 22370 13240 22376 13252
rect 21744 13212 22376 13240
rect 18785 13203 18843 13209
rect 22370 13200 22376 13212
rect 22428 13240 22434 13252
rect 22646 13240 22652 13252
rect 22428 13212 22652 13240
rect 22428 13200 22434 13212
rect 22646 13200 22652 13212
rect 22704 13200 22710 13252
rect 23753 13243 23811 13249
rect 23753 13209 23765 13243
rect 23799 13240 23811 13243
rect 24210 13240 24216 13252
rect 23799 13212 24216 13240
rect 23799 13209 23811 13212
rect 23753 13203 23811 13209
rect 24210 13200 24216 13212
rect 24268 13200 24274 13252
rect 13412 13144 14228 13172
rect 14277 13175 14335 13181
rect 13412 13132 13418 13144
rect 14277 13141 14289 13175
rect 14323 13172 14335 13175
rect 14366 13172 14372 13184
rect 14323 13144 14372 13172
rect 14323 13141 14335 13144
rect 14277 13135 14335 13141
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15562 13172 15568 13184
rect 15335 13144 15568 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 16574 13132 16580 13184
rect 16632 13132 16638 13184
rect 17126 13132 17132 13184
rect 17184 13132 17190 13184
rect 17497 13175 17555 13181
rect 17497 13141 17509 13175
rect 17543 13172 17555 13175
rect 17586 13172 17592 13184
rect 17543 13144 17592 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 17770 13132 17776 13184
rect 17828 13172 17834 13184
rect 18141 13175 18199 13181
rect 18141 13172 18153 13175
rect 17828 13144 18153 13172
rect 17828 13132 17834 13144
rect 18141 13141 18153 13144
rect 18187 13141 18199 13175
rect 18141 13135 18199 13141
rect 18414 13132 18420 13184
rect 18472 13132 18478 13184
rect 18598 13132 18604 13184
rect 18656 13172 18662 13184
rect 22830 13172 22836 13184
rect 18656 13144 22836 13172
rect 18656 13132 18662 13144
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 29546 13132 29552 13184
rect 29604 13132 29610 13184
rect 552 13082 31648 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 11436 13082
rect 11488 13030 11500 13082
rect 11552 13030 11564 13082
rect 11616 13030 11628 13082
rect 11680 13030 11692 13082
rect 11744 13030 19210 13082
rect 19262 13030 19274 13082
rect 19326 13030 19338 13082
rect 19390 13030 19402 13082
rect 19454 13030 19466 13082
rect 19518 13030 26984 13082
rect 27036 13030 27048 13082
rect 27100 13030 27112 13082
rect 27164 13030 27176 13082
rect 27228 13030 27240 13082
rect 27292 13030 31648 13082
rect 552 13008 31648 13030
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 9364 12940 9505 12968
rect 9364 12928 9370 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 9493 12931 9551 12937
rect 12897 12971 12955 12977
rect 12897 12937 12909 12971
rect 12943 12968 12955 12971
rect 15102 12968 15108 12980
rect 12943 12940 15108 12968
rect 12943 12937 12955 12940
rect 12897 12931 12955 12937
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 15562 12928 15568 12980
rect 15620 12928 15626 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 18049 12971 18107 12977
rect 18049 12968 18061 12971
rect 16080 12940 18061 12968
rect 16080 12928 16086 12940
rect 18049 12937 18061 12940
rect 18095 12968 18107 12971
rect 18230 12968 18236 12980
rect 18095 12940 18236 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 18322 12928 18328 12980
rect 18380 12968 18386 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 18380 12940 18889 12968
rect 18380 12928 18386 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 18877 12931 18935 12937
rect 19058 12928 19064 12980
rect 19116 12928 19122 12980
rect 29638 12928 29644 12980
rect 29696 12968 29702 12980
rect 30653 12971 30711 12977
rect 30653 12968 30665 12971
rect 29696 12940 30665 12968
rect 29696 12928 29702 12940
rect 30653 12937 30665 12940
rect 30699 12968 30711 12971
rect 31018 12968 31024 12980
rect 30699 12940 31024 12968
rect 30699 12937 30711 12940
rect 30653 12931 30711 12937
rect 31018 12928 31024 12940
rect 31076 12928 31082 12980
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3053 12903 3111 12909
rect 3053 12900 3065 12903
rect 2924 12872 3065 12900
rect 2924 12860 2930 12872
rect 3053 12869 3065 12872
rect 3099 12900 3111 12903
rect 13814 12900 13820 12912
rect 3099 12872 3372 12900
rect 3099 12869 3111 12872
rect 3053 12863 3111 12869
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 3344 12773 3372 12872
rect 8680 12872 13820 12900
rect 8202 12832 8208 12844
rect 7024 12804 8208 12832
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12764 1547 12767
rect 1673 12767 1731 12773
rect 1673 12764 1685 12767
rect 1535 12736 1685 12764
rect 1535 12733 1547 12736
rect 1489 12727 1547 12733
rect 1673 12733 1685 12736
rect 1719 12733 1731 12767
rect 1673 12727 1731 12733
rect 3329 12767 3387 12773
rect 3329 12733 3341 12767
rect 3375 12764 3387 12767
rect 4525 12767 4583 12773
rect 4525 12764 4537 12767
rect 3375 12736 4537 12764
rect 3375 12733 3387 12736
rect 3329 12727 3387 12733
rect 4525 12733 4537 12736
rect 4571 12733 4583 12767
rect 4525 12727 4583 12733
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 7024 12773 7052 12804
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 7009 12767 7067 12773
rect 7009 12764 7021 12767
rect 5500 12736 7021 12764
rect 5500 12724 5506 12736
rect 7009 12733 7021 12736
rect 7055 12733 7067 12767
rect 7009 12727 7067 12733
rect 7098 12724 7104 12776
rect 7156 12724 7162 12776
rect 8110 12724 8116 12776
rect 8168 12724 8174 12776
rect 8680 12773 8708 12872
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 15473 12903 15531 12909
rect 15473 12869 15485 12903
rect 15519 12900 15531 12903
rect 16301 12903 16359 12909
rect 15519 12872 16160 12900
rect 15519 12869 15531 12872
rect 15473 12863 15531 12869
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 9456 12804 11192 12832
rect 9456 12792 9462 12804
rect 8665 12767 8723 12773
rect 8665 12733 8677 12767
rect 8711 12733 8723 12767
rect 8665 12727 8723 12733
rect 8757 12767 8815 12773
rect 8757 12733 8769 12767
rect 8803 12733 8815 12767
rect 8757 12727 8815 12733
rect 1946 12705 1952 12708
rect 1940 12659 1952 12705
rect 1946 12656 1952 12659
rect 2004 12656 2010 12708
rect 2958 12656 2964 12708
rect 3016 12696 3022 12708
rect 3973 12699 4031 12705
rect 3973 12696 3985 12699
rect 3016 12668 3985 12696
rect 3016 12656 3022 12668
rect 3973 12665 3985 12668
rect 4019 12665 4031 12699
rect 3973 12659 4031 12665
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 7331 12668 7573 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7561 12665 7573 12668
rect 7607 12665 7619 12699
rect 8772 12696 8800 12727
rect 8846 12724 8852 12776
rect 8904 12724 8910 12776
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12764 9091 12767
rect 9306 12764 9312 12776
rect 9079 12736 9312 12764
rect 9079 12733 9091 12736
rect 9033 12727 9091 12733
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 10042 12724 10048 12776
rect 10100 12724 10106 12776
rect 11164 12764 11192 12804
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11296 12804 11560 12832
rect 11296 12792 11302 12804
rect 11532 12773 11560 12804
rect 12084 12804 12480 12832
rect 11363 12767 11421 12773
rect 11363 12764 11375 12767
rect 11164 12736 11375 12764
rect 11363 12733 11375 12736
rect 11409 12733 11421 12767
rect 11363 12727 11421 12733
rect 11517 12767 11575 12773
rect 11517 12733 11529 12767
rect 11563 12764 11575 12767
rect 11974 12764 11980 12776
rect 11563 12736 11980 12764
rect 11563 12733 11575 12736
rect 11517 12727 11575 12733
rect 9122 12696 9128 12708
rect 8772 12668 9128 12696
rect 7561 12659 7619 12665
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 11378 12696 11406 12727
rect 11974 12724 11980 12736
rect 12032 12764 12038 12776
rect 12084 12773 12112 12804
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 12032 12736 12081 12764
rect 12032 12724 12038 12736
rect 12069 12733 12081 12736
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12733 12311 12767
rect 12452 12764 12480 12804
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 12952 12804 13737 12832
rect 12952 12792 12958 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 16022 12832 16028 12844
rect 13725 12795 13783 12801
rect 15764 12804 16028 12832
rect 12526 12764 12532 12776
rect 12452 12736 12532 12764
rect 12253 12727 12311 12733
rect 11698 12696 11704 12708
rect 11378 12668 11704 12696
rect 11698 12656 11704 12668
rect 11756 12696 11762 12708
rect 12268 12696 12296 12727
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 12618 12724 12624 12776
rect 12676 12724 12682 12776
rect 12710 12724 12716 12776
rect 12768 12764 12774 12776
rect 13262 12764 13268 12776
rect 12768 12736 13268 12764
rect 12768 12724 12774 12736
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13504 12736 13645 12764
rect 13504 12724 13510 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13740 12764 13768 12795
rect 13909 12767 13967 12773
rect 13740 12736 13860 12764
rect 13633 12727 13691 12733
rect 12728 12696 12756 12724
rect 13078 12696 13084 12708
rect 11756 12668 12756 12696
rect 12820 12668 13084 12696
rect 11756 12656 11762 12668
rect 3878 12588 3884 12640
rect 3936 12588 3942 12640
rect 6914 12588 6920 12640
rect 6972 12588 6978 12640
rect 7469 12631 7527 12637
rect 7469 12597 7481 12631
rect 7515 12628 7527 12631
rect 8018 12628 8024 12640
rect 7515 12600 8024 12628
rect 7515 12597 7527 12600
rect 7469 12591 7527 12597
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8389 12631 8447 12637
rect 8389 12597 8401 12631
rect 8435 12628 8447 12631
rect 8478 12628 8484 12640
rect 8435 12600 8484 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 11149 12631 11207 12637
rect 11149 12597 11161 12631
rect 11195 12628 11207 12631
rect 11238 12628 11244 12640
rect 11195 12600 11244 12628
rect 11195 12597 11207 12600
rect 11149 12591 11207 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12820 12628 12848 12668
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 13541 12699 13599 12705
rect 13541 12665 13553 12699
rect 13587 12696 13599 12699
rect 13722 12696 13728 12708
rect 13587 12668 13728 12696
rect 13587 12665 13599 12668
rect 13541 12659 13599 12665
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 13832 12696 13860 12736
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 13998 12764 14004 12776
rect 13955 12736 14004 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14090 12724 14096 12776
rect 14148 12724 14154 12776
rect 14366 12773 14372 12776
rect 14360 12764 14372 12773
rect 14327 12736 14372 12764
rect 14360 12727 14372 12736
rect 14366 12724 14372 12727
rect 14424 12724 14430 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 15764 12773 15792 12804
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16132 12773 16160 12872
rect 16301 12869 16313 12903
rect 16347 12900 16359 12903
rect 16482 12900 16488 12912
rect 16347 12872 16488 12900
rect 16347 12869 16359 12872
rect 16301 12863 16359 12869
rect 15565 12767 15623 12773
rect 15565 12764 15577 12767
rect 15528 12736 15577 12764
rect 15528 12724 15534 12736
rect 15565 12733 15577 12736
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 15749 12767 15807 12773
rect 15749 12733 15761 12767
rect 15795 12733 15807 12767
rect 15749 12727 15807 12733
rect 15841 12767 15899 12773
rect 15841 12733 15853 12767
rect 15887 12733 15899 12767
rect 15841 12727 15899 12733
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12733 16175 12767
rect 16117 12727 16175 12733
rect 15764 12696 15792 12727
rect 13832 12668 14136 12696
rect 12299 12600 12848 12628
rect 13817 12631 13875 12637
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 13998 12628 14004 12640
rect 13863 12600 14004 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 14108 12628 14136 12668
rect 15396 12668 15792 12696
rect 15856 12696 15884 12727
rect 16316 12696 16344 12863
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 17494 12909 17500 12912
rect 17451 12903 17500 12909
rect 17451 12869 17463 12903
rect 17497 12869 17500 12903
rect 17451 12863 17500 12869
rect 17494 12860 17500 12863
rect 17552 12860 17558 12912
rect 17589 12903 17647 12909
rect 17589 12869 17601 12903
rect 17635 12900 17647 12903
rect 17865 12903 17923 12909
rect 17865 12900 17877 12903
rect 17635 12872 17877 12900
rect 17635 12869 17647 12872
rect 17589 12863 17647 12869
rect 17865 12869 17877 12872
rect 17911 12869 17923 12903
rect 17865 12863 17923 12869
rect 18138 12860 18144 12912
rect 18196 12900 18202 12912
rect 20346 12900 20352 12912
rect 18196 12872 20352 12900
rect 18196 12860 18202 12872
rect 20346 12860 20352 12872
rect 20404 12860 20410 12912
rect 26053 12903 26111 12909
rect 26053 12869 26065 12903
rect 26099 12900 26111 12903
rect 26694 12900 26700 12912
rect 26099 12872 26700 12900
rect 26099 12869 26111 12872
rect 26053 12863 26111 12869
rect 26694 12860 26700 12872
rect 26752 12860 26758 12912
rect 28721 12835 28779 12841
rect 17604 12804 18736 12832
rect 17604 12776 17632 12804
rect 17218 12724 17224 12776
rect 17276 12724 17282 12776
rect 17310 12724 17316 12776
rect 17368 12724 17374 12776
rect 17586 12724 17592 12776
rect 17644 12724 17650 12776
rect 17773 12767 17831 12773
rect 17773 12733 17785 12767
rect 17819 12764 17831 12767
rect 17862 12764 17868 12776
rect 17819 12736 17868 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18046 12724 18052 12776
rect 18104 12724 18110 12776
rect 18138 12724 18144 12776
rect 18196 12724 18202 12776
rect 15856 12668 16344 12696
rect 17681 12699 17739 12705
rect 15396 12628 15424 12668
rect 17681 12665 17693 12699
rect 17727 12696 17739 12699
rect 17727 12668 18368 12696
rect 17727 12665 17739 12668
rect 17681 12659 17739 12665
rect 14108 12600 15424 12628
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 16025 12631 16083 12637
rect 16025 12628 16037 12631
rect 15528 12600 16037 12628
rect 15528 12588 15534 12600
rect 16025 12597 16037 12600
rect 16071 12597 16083 12631
rect 16025 12591 16083 12597
rect 16577 12631 16635 12637
rect 16577 12597 16589 12631
rect 16623 12628 16635 12631
rect 16666 12628 16672 12640
rect 16623 12600 16672 12628
rect 16623 12597 16635 12600
rect 16577 12591 16635 12597
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 18340 12628 18368 12668
rect 18506 12656 18512 12708
rect 18564 12656 18570 12708
rect 18708 12705 18736 12804
rect 28721 12801 28733 12835
rect 28767 12832 28779 12835
rect 29273 12835 29331 12841
rect 29273 12832 29285 12835
rect 28767 12804 29285 12832
rect 28767 12801 28779 12804
rect 28721 12795 28779 12801
rect 29273 12801 29285 12804
rect 29319 12801 29331 12835
rect 29273 12795 29331 12801
rect 25958 12724 25964 12776
rect 26016 12724 26022 12776
rect 26142 12724 26148 12776
rect 26200 12724 26206 12776
rect 26326 12724 26332 12776
rect 26384 12764 26390 12776
rect 26421 12767 26479 12773
rect 26421 12764 26433 12767
rect 26384 12736 26433 12764
rect 26384 12724 26390 12736
rect 26421 12733 26433 12736
rect 26467 12733 26479 12767
rect 26421 12727 26479 12733
rect 26697 12767 26755 12773
rect 26697 12733 26709 12767
rect 26743 12733 26755 12767
rect 26697 12727 26755 12733
rect 18693 12699 18751 12705
rect 18693 12665 18705 12699
rect 18739 12665 18751 12699
rect 18693 12659 18751 12665
rect 24854 12656 24860 12708
rect 24912 12696 24918 12708
rect 26712 12696 26740 12727
rect 28074 12724 28080 12776
rect 28132 12764 28138 12776
rect 29546 12773 29552 12776
rect 28629 12767 28687 12773
rect 28629 12764 28641 12767
rect 28132 12736 28641 12764
rect 28132 12724 28138 12736
rect 28629 12733 28641 12736
rect 28675 12764 28687 12767
rect 28997 12767 29055 12773
rect 28997 12764 29009 12767
rect 28675 12736 29009 12764
rect 28675 12733 28687 12736
rect 28629 12727 28687 12733
rect 28997 12733 29009 12736
rect 29043 12733 29055 12767
rect 29540 12764 29552 12773
rect 29507 12736 29552 12764
rect 28997 12727 29055 12733
rect 29540 12727 29552 12736
rect 29546 12724 29552 12727
rect 29604 12724 29610 12776
rect 24912 12668 26740 12696
rect 24912 12656 24918 12668
rect 18893 12631 18951 12637
rect 18893 12628 18905 12631
rect 18340 12600 18905 12628
rect 18893 12597 18905 12600
rect 18939 12597 18951 12631
rect 18893 12591 18951 12597
rect 26326 12588 26332 12640
rect 26384 12588 26390 12640
rect 26418 12588 26424 12640
rect 26476 12628 26482 12640
rect 26605 12631 26663 12637
rect 26605 12628 26617 12631
rect 26476 12600 26617 12628
rect 26476 12588 26482 12600
rect 26605 12597 26617 12600
rect 26651 12597 26663 12631
rect 26605 12591 26663 12597
rect 29086 12588 29092 12640
rect 29144 12588 29150 12640
rect 552 12538 31648 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 12096 12538
rect 12148 12486 12160 12538
rect 12212 12486 12224 12538
rect 12276 12486 12288 12538
rect 12340 12486 12352 12538
rect 12404 12486 19870 12538
rect 19922 12486 19934 12538
rect 19986 12486 19998 12538
rect 20050 12486 20062 12538
rect 20114 12486 20126 12538
rect 20178 12486 27644 12538
rect 27696 12486 27708 12538
rect 27760 12486 27772 12538
rect 27824 12486 27836 12538
rect 27888 12486 27900 12538
rect 27952 12486 31648 12538
rect 552 12464 31648 12486
rect 2976 12396 3372 12424
rect 2853 12359 2911 12365
rect 2853 12356 2865 12359
rect 2240 12328 2865 12356
rect 1946 12180 1952 12232
rect 2004 12180 2010 12232
rect 2240 12229 2268 12328
rect 2853 12325 2865 12328
rect 2899 12356 2911 12359
rect 2976 12356 3004 12396
rect 2899 12328 3004 12356
rect 3053 12359 3111 12365
rect 2899 12325 2911 12328
rect 2853 12319 2911 12325
rect 3053 12325 3065 12359
rect 3099 12356 3111 12359
rect 3344 12356 3372 12396
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 3936 12396 4077 12424
rect 3936 12384 3942 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 6914 12424 6920 12436
rect 4065 12387 4123 12393
rect 6748 12396 6920 12424
rect 3510 12356 3516 12368
rect 3099 12328 3280 12356
rect 3344 12328 3516 12356
rect 3099 12325 3111 12328
rect 3053 12319 3111 12325
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2958 12288 2964 12300
rect 2363 12260 2964 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 3252 12232 3280 12328
rect 3510 12316 3516 12328
rect 3568 12356 3574 12368
rect 3568 12328 4200 12356
rect 3568 12316 3574 12328
rect 4172 12297 4200 12328
rect 4264 12328 5396 12356
rect 3789 12291 3847 12297
rect 3789 12257 3801 12291
rect 3835 12288 3847 12291
rect 3881 12291 3939 12297
rect 3881 12288 3893 12291
rect 3835 12260 3893 12288
rect 3835 12257 3847 12260
rect 3789 12251 3847 12257
rect 3881 12257 3893 12260
rect 3927 12257 3939 12291
rect 3881 12251 3939 12257
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 4062 12220 4068 12232
rect 3476 12192 4068 12220
rect 3476 12180 3482 12192
rect 4062 12180 4068 12192
rect 4120 12220 4126 12232
rect 4264 12220 4292 12328
rect 5258 12297 5264 12300
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 5231 12291 5264 12297
rect 5231 12257 5243 12291
rect 5231 12251 5264 12257
rect 4120 12192 4292 12220
rect 4120 12180 4126 12192
rect 4982 12180 4988 12232
rect 5040 12220 5046 12232
rect 5092 12220 5120 12251
rect 5258 12248 5264 12251
rect 5316 12248 5322 12300
rect 5368 12288 5396 12328
rect 6027 12291 6085 12297
rect 6027 12288 6039 12291
rect 5368 12260 6039 12288
rect 6027 12257 6039 12260
rect 6073 12257 6085 12291
rect 6027 12251 6085 12257
rect 6178 12248 6184 12300
rect 6236 12248 6242 12300
rect 6748 12297 6776 12396
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 8110 12384 8116 12436
rect 8168 12384 8174 12436
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 9769 12427 9827 12433
rect 9769 12424 9781 12427
rect 9548 12396 9781 12424
rect 9548 12384 9554 12396
rect 9769 12393 9781 12396
rect 9815 12393 9827 12427
rect 9769 12387 9827 12393
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11204 12396 12434 12424
rect 11204 12384 11210 12396
rect 8128 12356 8156 12384
rect 8478 12365 8484 12368
rect 8472 12356 8484 12365
rect 6840 12328 8156 12356
rect 8439 12328 8484 12356
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12257 6791 12291
rect 6733 12251 6791 12257
rect 6840 12220 6868 12328
rect 8472 12319 8484 12328
rect 8478 12316 8484 12319
rect 8536 12316 8542 12368
rect 10042 12356 10048 12368
rect 9600 12328 10048 12356
rect 7000 12291 7058 12297
rect 7000 12257 7012 12291
rect 7046 12288 7058 12291
rect 7558 12288 7564 12300
rect 7046 12260 7564 12288
rect 7046 12257 7058 12260
rect 7000 12251 7058 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 8294 12288 8300 12300
rect 8251 12260 8300 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 5040 12192 6868 12220
rect 5040 12180 5046 12192
rect 5442 12112 5448 12164
rect 5500 12152 5506 12164
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 5500 12124 5825 12152
rect 5500 12112 5506 12124
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 2682 12044 2688 12096
rect 2740 12044 2746 12096
rect 2866 12044 2872 12096
rect 2924 12044 2930 12096
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 3881 12087 3939 12093
rect 3881 12084 3893 12087
rect 3476 12056 3893 12084
rect 3476 12044 3482 12056
rect 3881 12053 3893 12056
rect 3927 12053 3939 12087
rect 3881 12047 3939 12053
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 5534 12084 5540 12096
rect 5307 12056 5540 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 9600 12093 9628 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 11054 12316 11060 12368
rect 11112 12356 11118 12368
rect 11977 12359 12035 12365
rect 11977 12356 11989 12359
rect 11112 12328 11989 12356
rect 11112 12316 11118 12328
rect 11977 12325 11989 12328
rect 12023 12325 12035 12359
rect 12406 12356 12434 12396
rect 13630 12384 13636 12436
rect 13688 12384 13694 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 14148 12396 14289 12424
rect 14148 12384 14154 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 14366 12384 14372 12436
rect 14424 12424 14430 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 14424 12396 14473 12424
rect 14424 12384 14430 12396
rect 14461 12393 14473 12396
rect 14507 12424 14519 12427
rect 15562 12424 15568 12436
rect 14507 12396 15568 12424
rect 14507 12393 14519 12396
rect 14461 12387 14519 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17402 12424 17408 12436
rect 17276 12396 17408 12424
rect 17276 12384 17282 12396
rect 17402 12384 17408 12396
rect 17460 12424 17466 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17460 12396 17509 12424
rect 17460 12384 17466 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 17497 12387 17555 12393
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 19153 12427 19211 12433
rect 19153 12424 19165 12427
rect 18012 12396 19165 12424
rect 18012 12384 18018 12396
rect 19153 12393 19165 12396
rect 19199 12393 19211 12427
rect 19153 12387 19211 12393
rect 15746 12356 15752 12368
rect 12406 12328 14412 12356
rect 11977 12319 12035 12325
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 10597 12291 10655 12297
rect 10597 12257 10609 12291
rect 10643 12257 10655 12291
rect 10597 12251 10655 12257
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11149 12291 11207 12297
rect 11149 12288 11161 12291
rect 10827 12260 11161 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11149 12257 11161 12260
rect 11195 12288 11207 12291
rect 11238 12288 11244 12300
rect 11195 12260 11244 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 9876 12152 9904 12251
rect 10612 12220 10640 12251
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 11348 12220 11376 12251
rect 11698 12248 11704 12300
rect 11756 12248 11762 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 12066 12288 12072 12300
rect 11848 12260 12072 12288
rect 11848 12248 11854 12260
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 12216 12260 12449 12288
rect 12216 12248 12222 12260
rect 12437 12257 12449 12260
rect 12483 12288 12495 12291
rect 12713 12291 12771 12297
rect 12713 12288 12725 12291
rect 12483 12260 12725 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 12713 12257 12725 12260
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 12894 12248 12900 12300
rect 12952 12248 12958 12300
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 14384 12297 14412 12328
rect 14844 12328 15752 12356
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 13320 12260 13461 12288
rect 13320 12248 13326 12260
rect 13449 12257 13461 12260
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 14369 12291 14427 12297
rect 14369 12257 14381 12291
rect 14415 12257 14427 12291
rect 14369 12251 14427 12257
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 14844 12297 14872 12328
rect 15746 12316 15752 12328
rect 15804 12356 15810 12368
rect 16574 12356 16580 12368
rect 15804 12328 15973 12356
rect 15804 12316 15810 12328
rect 14675 12291 14733 12297
rect 14675 12288 14687 12291
rect 14608 12260 14687 12288
rect 14608 12248 14614 12260
rect 14675 12257 14687 12260
rect 14721 12257 14733 12291
rect 14675 12251 14733 12257
rect 14829 12291 14887 12297
rect 14829 12257 14841 12291
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15565 12291 15623 12297
rect 15565 12288 15577 12291
rect 15344 12260 15577 12288
rect 15344 12248 15350 12260
rect 15565 12257 15577 12260
rect 15611 12288 15623 12291
rect 15654 12288 15660 12300
rect 15611 12260 15660 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15304 12220 15332 12248
rect 10612 12192 12572 12220
rect 12544 12164 12572 12192
rect 12636 12192 15332 12220
rect 9876 12124 11560 12152
rect 9585 12087 9643 12093
rect 9585 12084 9597 12087
rect 6236 12056 9597 12084
rect 6236 12044 6242 12056
rect 9585 12053 9597 12056
rect 9631 12053 9643 12087
rect 9585 12047 9643 12053
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 10781 12087 10839 12093
rect 10781 12084 10793 12087
rect 9916 12056 10793 12084
rect 9916 12044 9922 12056
rect 10781 12053 10793 12056
rect 10827 12053 10839 12087
rect 10781 12047 10839 12053
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 11425 12087 11483 12093
rect 11425 12084 11437 12087
rect 11296 12056 11437 12084
rect 11296 12044 11302 12056
rect 11425 12053 11437 12056
rect 11471 12053 11483 12087
rect 11532 12084 11560 12124
rect 12526 12112 12532 12164
rect 12584 12112 12590 12164
rect 12636 12084 12664 12192
rect 15378 12112 15384 12164
rect 15436 12152 15442 12164
rect 15746 12152 15752 12164
rect 15436 12124 15752 12152
rect 15436 12112 15442 12124
rect 15746 12112 15752 12124
rect 15804 12112 15810 12164
rect 11532 12056 12664 12084
rect 11425 12047 11483 12053
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 15838 12084 15844 12096
rect 13872 12056 15844 12084
rect 13872 12044 13878 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 15945 12084 15973 12328
rect 16132 12328 16580 12356
rect 16132 12297 16160 12328
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 18040 12359 18098 12365
rect 18040 12325 18052 12359
rect 18086 12356 18098 12359
rect 18414 12356 18420 12368
rect 18086 12328 18420 12356
rect 18086 12325 18098 12328
rect 18040 12319 18098 12325
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 19168 12356 19196 12387
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19668 12396 19809 12424
rect 19668 12384 19674 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 25593 12427 25651 12433
rect 19797 12387 19855 12393
rect 22066 12396 22850 12424
rect 19168 12328 20208 12356
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 16206 12248 16212 12300
rect 16264 12288 16270 12300
rect 16373 12291 16431 12297
rect 16373 12288 16385 12291
rect 16264 12260 16385 12288
rect 16264 12248 16270 12260
rect 16373 12257 16385 12260
rect 16419 12257 16431 12291
rect 16373 12251 16431 12257
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17184 12260 17785 12288
rect 17184 12248 17190 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 17773 12251 17831 12257
rect 19058 12248 19064 12300
rect 19116 12288 19122 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19116 12260 19441 12288
rect 19116 12248 19122 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19702 12248 19708 12300
rect 19760 12248 19766 12300
rect 20180 12297 20208 12328
rect 20530 12316 20536 12368
rect 20588 12356 20594 12368
rect 22066 12365 22094 12396
rect 22051 12359 22109 12365
rect 22051 12356 22063 12359
rect 20588 12328 22063 12356
rect 20588 12316 20594 12328
rect 22051 12325 22063 12328
rect 22097 12325 22109 12359
rect 22051 12319 22109 12325
rect 22186 12316 22192 12368
rect 22244 12316 22250 12368
rect 22462 12356 22468 12368
rect 22296 12328 22468 12356
rect 22296 12297 22324 12328
rect 22462 12316 22468 12328
rect 22520 12316 22526 12368
rect 22554 12316 22560 12368
rect 22612 12316 22618 12368
rect 22822 12365 22850 12396
rect 25593 12393 25605 12427
rect 25639 12424 25651 12427
rect 25958 12424 25964 12436
rect 25639 12396 25964 12424
rect 25639 12393 25651 12396
rect 25593 12387 25651 12393
rect 25958 12384 25964 12396
rect 26016 12384 26022 12436
rect 27893 12427 27951 12433
rect 27893 12424 27905 12427
rect 26436 12396 27905 12424
rect 22807 12359 22865 12365
rect 22807 12325 22819 12359
rect 22853 12356 22865 12359
rect 25682 12356 25688 12368
rect 22853 12328 25688 12356
rect 22853 12325 22865 12328
rect 22807 12319 22865 12325
rect 25682 12316 25688 12328
rect 25740 12356 25746 12368
rect 26079 12359 26137 12365
rect 26079 12356 26091 12359
rect 25740 12328 26091 12356
rect 25740 12316 25746 12328
rect 26079 12325 26091 12328
rect 26125 12325 26137 12359
rect 26079 12319 26137 12325
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12288 20223 12291
rect 22281 12291 22339 12297
rect 20211 12260 22232 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 18932 12192 19625 12220
rect 18932 12180 18938 12192
rect 19613 12189 19625 12192
rect 19659 12220 19671 12223
rect 19886 12220 19892 12232
rect 19659 12192 19892 12220
rect 19659 12189 19671 12192
rect 19613 12183 19671 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 19996 12220 20024 12251
rect 22204 12232 22232 12260
rect 22281 12257 22293 12291
rect 22327 12257 22339 12291
rect 22572 12288 22600 12316
rect 22397 12287 22600 12288
rect 22281 12251 22339 12257
rect 22372 12281 22600 12287
rect 22372 12247 22384 12281
rect 22418 12260 22600 12281
rect 22649 12291 22707 12297
rect 22418 12247 22430 12260
rect 22649 12257 22661 12291
rect 22695 12288 22707 12291
rect 22925 12291 22983 12297
rect 22695 12260 22784 12288
rect 22695 12257 22707 12260
rect 22649 12251 22707 12257
rect 22372 12241 22430 12247
rect 22756 12232 22784 12260
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 20530 12220 20536 12232
rect 19996 12192 20536 12220
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 19245 12155 19303 12161
rect 19245 12152 19257 12155
rect 19024 12124 19257 12152
rect 19024 12112 19030 12124
rect 19245 12121 19257 12124
rect 19291 12121 19303 12155
rect 19245 12115 19303 12121
rect 20254 12112 20260 12164
rect 20312 12152 20318 12164
rect 20349 12155 20407 12161
rect 20349 12152 20361 12155
rect 20312 12124 20361 12152
rect 20312 12112 20318 12124
rect 20349 12121 20361 12124
rect 20395 12152 20407 12155
rect 20438 12152 20444 12164
rect 20395 12124 20444 12152
rect 20395 12121 20407 12124
rect 20349 12115 20407 12121
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 21928 12152 21956 12183
rect 22186 12180 22192 12232
rect 22244 12180 22250 12232
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 22830 12180 22836 12232
rect 22888 12220 22894 12232
rect 22940 12220 22968 12251
rect 23014 12248 23020 12300
rect 23072 12248 23078 12300
rect 23106 12248 23112 12300
rect 23164 12288 23170 12300
rect 24026 12288 24032 12300
rect 23164 12260 24032 12288
rect 23164 12248 23170 12260
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 25314 12288 25320 12300
rect 25271 12260 25320 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 25498 12248 25504 12300
rect 25556 12288 25562 12300
rect 25777 12291 25835 12297
rect 25777 12288 25789 12291
rect 25556 12260 25789 12288
rect 25556 12248 25562 12260
rect 25777 12257 25789 12260
rect 25823 12257 25835 12291
rect 25777 12251 25835 12257
rect 25866 12248 25872 12300
rect 25924 12248 25930 12300
rect 25958 12248 25964 12300
rect 26016 12248 26022 12300
rect 26237 12291 26295 12297
rect 26237 12257 26249 12291
rect 26283 12288 26295 12291
rect 26326 12288 26332 12300
rect 26283 12260 26332 12288
rect 26283 12257 26295 12260
rect 26237 12251 26295 12257
rect 26326 12248 26332 12260
rect 26384 12248 26390 12300
rect 26436 12297 26464 12396
rect 27893 12393 27905 12396
rect 27939 12424 27951 12427
rect 28626 12424 28632 12436
rect 27939 12396 28632 12424
rect 27939 12393 27951 12396
rect 27893 12387 27951 12393
rect 28626 12384 28632 12396
rect 28684 12384 28690 12436
rect 30742 12384 30748 12436
rect 30800 12384 30806 12436
rect 26510 12316 26516 12368
rect 26568 12356 26574 12368
rect 26568 12328 26740 12356
rect 26568 12316 26574 12328
rect 26421 12291 26479 12297
rect 26421 12257 26433 12291
rect 26467 12257 26479 12291
rect 26421 12251 26479 12257
rect 22888 12192 22968 12220
rect 25409 12223 25467 12229
rect 22888 12180 22894 12192
rect 25409 12189 25421 12223
rect 25455 12220 25467 12223
rect 26142 12220 26148 12232
rect 25455 12192 26148 12220
rect 25455 12189 25467 12192
rect 25409 12183 25467 12189
rect 26142 12180 26148 12192
rect 26200 12220 26206 12232
rect 26436 12220 26464 12251
rect 26602 12248 26608 12300
rect 26660 12248 26666 12300
rect 26712 12297 26740 12328
rect 28994 12316 29000 12368
rect 29052 12356 29058 12368
rect 29610 12359 29668 12365
rect 29610 12356 29622 12359
rect 29052 12328 29622 12356
rect 29052 12316 29058 12328
rect 29610 12325 29622 12328
rect 29656 12325 29668 12359
rect 29610 12319 29668 12325
rect 26697 12291 26755 12297
rect 26697 12257 26709 12291
rect 26743 12257 26755 12291
rect 26697 12251 26755 12257
rect 26789 12291 26847 12297
rect 26789 12257 26801 12291
rect 26835 12257 26847 12291
rect 26789 12251 26847 12257
rect 26200 12192 26464 12220
rect 26804 12220 26832 12251
rect 26878 12248 26884 12300
rect 26936 12288 26942 12300
rect 27249 12291 27307 12297
rect 27249 12288 27261 12291
rect 26936 12260 27261 12288
rect 26936 12248 26942 12260
rect 27249 12257 27261 12260
rect 27295 12257 27307 12291
rect 27249 12251 27307 12257
rect 27430 12248 27436 12300
rect 27488 12288 27494 12300
rect 27801 12291 27859 12297
rect 27801 12288 27813 12291
rect 27488 12260 27813 12288
rect 27488 12248 27494 12260
rect 27801 12257 27813 12260
rect 27847 12257 27859 12291
rect 27801 12251 27859 12257
rect 29086 12248 29092 12300
rect 29144 12288 29150 12300
rect 29365 12291 29423 12297
rect 29365 12288 29377 12291
rect 29144 12260 29377 12288
rect 29144 12248 29150 12260
rect 29365 12257 29377 12260
rect 29411 12257 29423 12291
rect 29365 12251 29423 12257
rect 27525 12223 27583 12229
rect 27525 12220 27537 12223
rect 26804 12192 27537 12220
rect 26200 12180 26206 12192
rect 20640 12124 21956 12152
rect 16114 12084 16120 12096
rect 15945 12056 16120 12084
rect 16114 12044 16120 12056
rect 16172 12084 16178 12096
rect 20640 12084 20668 12124
rect 25866 12112 25872 12164
rect 25924 12152 25930 12164
rect 26786 12152 26792 12164
rect 25924 12124 26792 12152
rect 25924 12112 25930 12124
rect 26786 12112 26792 12124
rect 26844 12112 26850 12164
rect 16172 12056 20668 12084
rect 16172 12044 16178 12056
rect 21450 12044 21456 12096
rect 21508 12084 21514 12096
rect 22557 12087 22615 12093
rect 22557 12084 22569 12087
rect 21508 12056 22569 12084
rect 21508 12044 21514 12056
rect 22557 12053 22569 12056
rect 22603 12053 22615 12087
rect 22557 12047 22615 12053
rect 23293 12087 23351 12093
rect 23293 12053 23305 12087
rect 23339 12084 23351 12087
rect 23382 12084 23388 12096
rect 23339 12056 23388 12084
rect 23339 12053 23351 12056
rect 23293 12047 23351 12053
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 25038 12044 25044 12096
rect 25096 12044 25102 12096
rect 25774 12044 25780 12096
rect 25832 12084 25838 12096
rect 25958 12084 25964 12096
rect 25832 12056 25964 12084
rect 25832 12044 25838 12056
rect 25958 12044 25964 12056
rect 26016 12084 26022 12096
rect 26896 12084 26924 12192
rect 27525 12189 27537 12192
rect 27571 12189 27583 12223
rect 27525 12183 27583 12189
rect 27065 12155 27123 12161
rect 27065 12121 27077 12155
rect 27111 12152 27123 12155
rect 27706 12152 27712 12164
rect 27111 12124 27712 12152
rect 27111 12121 27123 12124
rect 27065 12115 27123 12121
rect 27706 12112 27712 12124
rect 27764 12112 27770 12164
rect 26016 12056 26924 12084
rect 26016 12044 26022 12056
rect 552 11994 31648 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 11436 11994
rect 11488 11942 11500 11994
rect 11552 11942 11564 11994
rect 11616 11942 11628 11994
rect 11680 11942 11692 11994
rect 11744 11942 19210 11994
rect 19262 11942 19274 11994
rect 19326 11942 19338 11994
rect 19390 11942 19402 11994
rect 19454 11942 19466 11994
rect 19518 11942 26984 11994
rect 27036 11942 27048 11994
rect 27100 11942 27112 11994
rect 27164 11942 27176 11994
rect 27228 11942 27240 11994
rect 27292 11942 31648 11994
rect 552 11920 31648 11942
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3234 11880 3240 11892
rect 3099 11852 3240 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3234 11840 3240 11852
rect 3292 11880 3298 11892
rect 4157 11883 4215 11889
rect 4157 11880 4169 11883
rect 3292 11852 4169 11880
rect 3292 11840 3298 11852
rect 4157 11849 4169 11852
rect 4203 11880 4215 11883
rect 4246 11880 4252 11892
rect 4203 11852 4252 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 5350 11880 5356 11892
rect 4663 11852 5356 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 7558 11840 7564 11892
rect 7616 11840 7622 11892
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 16577 11883 16635 11889
rect 16577 11880 16589 11883
rect 12492 11852 16589 11880
rect 12492 11840 12498 11852
rect 16577 11849 16589 11852
rect 16623 11880 16635 11883
rect 19794 11880 19800 11892
rect 16623 11852 19800 11880
rect 16623 11849 16635 11852
rect 16577 11843 16635 11849
rect 19794 11840 19800 11852
rect 19852 11880 19858 11892
rect 21266 11880 21272 11892
rect 19852 11852 21272 11880
rect 19852 11840 19858 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 22646 11840 22652 11892
rect 22704 11880 22710 11892
rect 23109 11883 23167 11889
rect 23109 11880 23121 11883
rect 22704 11852 23121 11880
rect 22704 11840 22710 11852
rect 23109 11849 23121 11852
rect 23155 11849 23167 11883
rect 23109 11843 23167 11849
rect 26605 11883 26663 11889
rect 26605 11849 26617 11883
rect 26651 11880 26663 11883
rect 26878 11880 26884 11892
rect 26651 11852 26884 11880
rect 26651 11849 26663 11852
rect 26605 11843 26663 11849
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 27982 11880 27988 11892
rect 27080 11852 27988 11880
rect 4982 11772 4988 11824
rect 5040 11772 5046 11824
rect 5258 11812 5264 11824
rect 5092 11784 5264 11812
rect 2866 11704 2872 11756
rect 2924 11744 2930 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 2924 11716 3985 11744
rect 2924 11704 2930 11716
rect 3973 11713 3985 11716
rect 4019 11744 4031 11747
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 4019 11716 4721 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4709 11713 4721 11716
rect 4755 11744 4767 11747
rect 5092 11744 5120 11784
rect 5258 11772 5264 11784
rect 5316 11772 5322 11824
rect 16025 11815 16083 11821
rect 16025 11781 16037 11815
rect 16071 11812 16083 11815
rect 16206 11812 16212 11824
rect 16071 11784 16212 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 17126 11772 17132 11824
rect 17184 11812 17190 11824
rect 18138 11812 18144 11824
rect 17184 11784 18144 11812
rect 17184 11772 17190 11784
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 20530 11772 20536 11824
rect 20588 11772 20594 11824
rect 26050 11772 26056 11824
rect 26108 11812 26114 11824
rect 27080 11812 27108 11852
rect 27982 11840 27988 11852
rect 28040 11880 28046 11892
rect 28261 11883 28319 11889
rect 28261 11880 28273 11883
rect 28040 11852 28273 11880
rect 28040 11840 28046 11852
rect 28261 11849 28273 11852
rect 28307 11849 28319 11883
rect 28261 11843 28319 11849
rect 26108 11784 27108 11812
rect 26108 11772 26114 11784
rect 4755 11716 5120 11744
rect 5169 11747 5227 11753
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 8846 11744 8852 11756
rect 5169 11707 5227 11713
rect 7852 11716 8852 11744
rect 1305 11679 1363 11685
rect 1305 11645 1317 11679
rect 1351 11676 1363 11679
rect 1394 11676 1400 11688
rect 1351 11648 1400 11676
rect 1351 11645 1363 11648
rect 1305 11639 1363 11645
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 1489 11679 1547 11685
rect 1489 11645 1501 11679
rect 1535 11676 1547 11679
rect 1673 11679 1731 11685
rect 1673 11676 1685 11679
rect 1535 11648 1685 11676
rect 1535 11645 1547 11648
rect 1489 11639 1547 11645
rect 1673 11645 1685 11648
rect 1719 11645 1731 11679
rect 1673 11639 1731 11645
rect 2682 11636 2688 11688
rect 2740 11676 2746 11688
rect 3237 11679 3295 11685
rect 3237 11676 3249 11679
rect 2740 11648 3249 11676
rect 2740 11636 2746 11648
rect 3237 11645 3249 11648
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 3418 11636 3424 11688
rect 3476 11636 3482 11688
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11676 3939 11679
rect 4062 11676 4068 11688
rect 3927 11648 4068 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4154 11636 4160 11688
rect 4212 11636 4218 11688
rect 4433 11679 4491 11685
rect 4433 11676 4445 11679
rect 4356 11648 4445 11676
rect 1940 11611 1998 11617
rect 1940 11577 1952 11611
rect 1986 11608 1998 11611
rect 3329 11611 3387 11617
rect 3329 11608 3341 11611
rect 1986 11580 3341 11608
rect 1986 11577 1998 11580
rect 1940 11571 1998 11577
rect 3329 11577 3341 11580
rect 3375 11577 3387 11611
rect 3329 11571 3387 11577
rect 1210 11500 1216 11552
rect 1268 11500 1274 11552
rect 4356 11549 4384 11648
rect 4433 11645 4445 11648
rect 4479 11645 4491 11679
rect 4433 11639 4491 11645
rect 4614 11636 4620 11688
rect 4672 11636 4678 11688
rect 5184 11676 5212 11707
rect 5442 11685 5448 11688
rect 5261 11679 5319 11685
rect 5261 11676 5273 11679
rect 5184 11648 5273 11676
rect 5261 11645 5273 11648
rect 5307 11645 5319 11679
rect 5261 11639 5319 11645
rect 5409 11679 5448 11685
rect 5409 11645 5421 11679
rect 5409 11639 5448 11645
rect 5442 11636 5448 11639
rect 5500 11636 5506 11688
rect 5534 11636 5540 11688
rect 5592 11636 5598 11688
rect 5718 11636 5724 11688
rect 5776 11685 5782 11688
rect 7852 11685 7880 11716
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 12066 11744 12072 11756
rect 11256 11716 12072 11744
rect 5776 11676 5784 11685
rect 7837 11679 7895 11685
rect 5776 11648 5821 11676
rect 5776 11639 5784 11648
rect 7837 11645 7849 11679
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 5776 11636 5782 11639
rect 5629 11611 5687 11617
rect 5629 11577 5641 11611
rect 5675 11608 5687 11611
rect 7944 11608 7972 11639
rect 8018 11636 8024 11688
rect 8076 11636 8082 11688
rect 8202 11636 8208 11688
rect 8260 11636 8266 11688
rect 9122 11676 9128 11688
rect 8312 11648 9128 11676
rect 8312 11608 8340 11648
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 9999 11648 10149 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10137 11645 10149 11648
rect 10183 11645 10195 11679
rect 10137 11639 10195 11645
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 11146 11676 11152 11688
rect 10275 11648 11152 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11256 11685 11284 11716
rect 12066 11704 12072 11716
rect 12124 11744 12130 11756
rect 12124 11716 12434 11744
rect 12124 11704 12130 11716
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11425 11679 11483 11685
rect 11425 11676 11437 11679
rect 11388 11648 11437 11676
rect 11388 11636 11394 11648
rect 11425 11645 11437 11648
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11645 11759 11679
rect 12406 11676 12434 11716
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 16666 11744 16672 11756
rect 15611 11716 16672 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 17678 11704 17684 11756
rect 17736 11744 17742 11756
rect 17862 11744 17868 11756
rect 17736 11716 17868 11744
rect 17736 11704 17742 11716
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 21269 11747 21327 11753
rect 21269 11744 21281 11747
rect 19944 11716 21281 11744
rect 19944 11704 19950 11716
rect 21269 11713 21281 11716
rect 21315 11744 21327 11747
rect 21315 11716 21864 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12406 11648 12633 11676
rect 11701 11639 11759 11645
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 5675 11580 6040 11608
rect 7944 11580 8340 11608
rect 5675 11577 5687 11580
rect 5629 11571 5687 11577
rect 4341 11543 4399 11549
rect 4341 11509 4353 11543
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 5902 11500 5908 11552
rect 5960 11500 5966 11552
rect 6012 11540 6040 11580
rect 8754 11568 8760 11620
rect 8812 11608 8818 11620
rect 9686 11611 9744 11617
rect 9686 11608 9698 11611
rect 8812 11580 9698 11608
rect 8812 11568 8818 11580
rect 9686 11577 9698 11580
rect 9732 11577 9744 11611
rect 11716 11608 11744 11639
rect 13078 11636 13084 11688
rect 13136 11636 13142 11688
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 18138 11676 18144 11688
rect 13403 11648 18144 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11645 18383 11679
rect 18325 11639 18383 11645
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 18463 11648 18889 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 11716 11580 12434 11608
rect 9686 11571 9744 11577
rect 6086 11540 6092 11552
rect 6012 11512 6092 11540
rect 6086 11500 6092 11512
rect 6144 11540 6150 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 6144 11512 8585 11540
rect 6144 11500 6150 11512
rect 8573 11509 8585 11512
rect 8619 11540 8631 11543
rect 9306 11540 9312 11552
rect 8619 11512 9312 11540
rect 8619 11509 8631 11512
rect 8573 11503 8631 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11848 11512 11897 11540
rect 11848 11500 11854 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 12406 11540 12434 11580
rect 17862 11568 17868 11620
rect 17920 11568 17926 11620
rect 18340 11608 18368 11639
rect 18966 11636 18972 11688
rect 19024 11676 19030 11688
rect 19133 11679 19191 11685
rect 19133 11676 19145 11679
rect 19024 11648 19145 11676
rect 19024 11636 19030 11648
rect 19133 11645 19145 11648
rect 19179 11645 19191 11679
rect 19133 11639 19191 11645
rect 20346 11636 20352 11688
rect 20404 11636 20410 11688
rect 21450 11636 21456 11688
rect 21508 11636 21514 11688
rect 21726 11636 21732 11688
rect 21784 11636 21790 11688
rect 21836 11676 21864 11716
rect 23290 11704 23296 11756
rect 23348 11744 23354 11756
rect 23569 11747 23627 11753
rect 23569 11744 23581 11747
rect 23348 11716 23581 11744
rect 23348 11704 23354 11716
rect 23569 11713 23581 11716
rect 23615 11713 23627 11747
rect 24854 11744 24860 11756
rect 23569 11707 23627 11713
rect 24688 11716 24860 11744
rect 21836 11648 22094 11676
rect 18782 11608 18788 11620
rect 18340 11580 18788 11608
rect 18782 11568 18788 11580
rect 18840 11568 18846 11620
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 20990 11608 20996 11620
rect 20220 11580 20996 11608
rect 20220 11568 20226 11580
rect 20990 11568 20996 11580
rect 21048 11568 21054 11620
rect 21637 11611 21695 11617
rect 21637 11577 21649 11611
rect 21683 11608 21695 11611
rect 21974 11611 22032 11617
rect 21974 11608 21986 11611
rect 21683 11580 21986 11608
rect 21683 11577 21695 11580
rect 21637 11571 21695 11577
rect 21974 11577 21986 11580
rect 22020 11577 22032 11611
rect 21974 11571 22032 11577
rect 12618 11540 12624 11552
rect 12406 11512 12624 11540
rect 11885 11503 11943 11509
rect 12618 11500 12624 11512
rect 12676 11540 12682 11552
rect 15194 11540 15200 11552
rect 12676 11512 15200 11540
rect 12676 11500 12682 11512
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 15657 11543 15715 11549
rect 15657 11509 15669 11543
rect 15703 11540 15715 11543
rect 15838 11540 15844 11552
rect 15703 11512 15844 11540
rect 15703 11509 15715 11512
rect 15657 11503 15715 11509
rect 15838 11500 15844 11512
rect 15896 11540 15902 11552
rect 16022 11540 16028 11552
rect 15896 11512 16028 11540
rect 15896 11500 15902 11512
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 20257 11543 20315 11549
rect 20257 11540 20269 11543
rect 19760 11512 20269 11540
rect 19760 11500 19766 11512
rect 20257 11509 20269 11512
rect 20303 11509 20315 11543
rect 22066 11540 22094 11648
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 23014 11676 23020 11688
rect 22520 11648 23020 11676
rect 22520 11636 22526 11648
rect 23014 11636 23020 11648
rect 23072 11636 23078 11688
rect 23382 11636 23388 11688
rect 23440 11636 23446 11688
rect 23658 11636 23664 11688
rect 23716 11676 23722 11688
rect 24688 11685 24716 11716
rect 24854 11704 24860 11716
rect 24912 11704 24918 11756
rect 23845 11679 23903 11685
rect 23845 11676 23857 11679
rect 23716 11648 23857 11676
rect 23716 11636 23722 11648
rect 23845 11645 23857 11648
rect 23891 11645 23903 11679
rect 23845 11639 23903 11645
rect 24673 11679 24731 11685
rect 24673 11645 24685 11679
rect 24719 11645 24731 11679
rect 24673 11639 24731 11645
rect 24765 11679 24823 11685
rect 24765 11645 24777 11679
rect 24811 11676 24823 11679
rect 24949 11679 25007 11685
rect 24949 11676 24961 11679
rect 24811 11648 24961 11676
rect 24811 11645 24823 11648
rect 24765 11639 24823 11645
rect 24949 11645 24961 11648
rect 24995 11645 25007 11679
rect 24949 11639 25007 11645
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 25205 11679 25263 11685
rect 25205 11676 25217 11679
rect 25096 11648 25217 11676
rect 25096 11636 25102 11648
rect 25205 11645 25217 11648
rect 25251 11645 25263 11679
rect 25205 11639 25263 11645
rect 27706 11636 27712 11688
rect 27764 11685 27770 11688
rect 27764 11676 27776 11685
rect 27985 11679 28043 11685
rect 27764 11648 27809 11676
rect 27764 11639 27776 11648
rect 27985 11645 27997 11679
rect 28031 11676 28043 11679
rect 28537 11679 28595 11685
rect 28537 11676 28549 11679
rect 28031 11648 28549 11676
rect 28031 11645 28043 11648
rect 27985 11639 28043 11645
rect 28537 11645 28549 11648
rect 28583 11645 28595 11679
rect 28537 11639 28595 11645
rect 28629 11679 28687 11685
rect 28629 11645 28641 11679
rect 28675 11676 28687 11679
rect 28994 11676 29000 11688
rect 28675 11648 29000 11676
rect 28675 11645 28687 11648
rect 28629 11639 28687 11645
rect 27764 11636 27770 11639
rect 28994 11636 29000 11648
rect 29052 11676 29058 11688
rect 29641 11679 29699 11685
rect 29641 11676 29653 11679
rect 29052 11648 29653 11676
rect 29052 11636 29058 11648
rect 29641 11645 29653 11648
rect 29687 11676 29699 11679
rect 30282 11676 30288 11688
rect 29687 11648 30288 11676
rect 29687 11645 29699 11648
rect 29641 11639 29699 11645
rect 30282 11636 30288 11648
rect 30340 11636 30346 11688
rect 30561 11679 30619 11685
rect 30561 11645 30573 11679
rect 30607 11676 30619 11679
rect 30834 11676 30840 11688
rect 30607 11648 30840 11676
rect 30607 11645 30619 11648
rect 30561 11639 30619 11645
rect 30834 11636 30840 11648
rect 30892 11636 30898 11688
rect 22186 11568 22192 11620
rect 22244 11608 22250 11620
rect 28169 11611 28227 11617
rect 28169 11608 28181 11611
rect 22244 11580 28181 11608
rect 22244 11568 22250 11580
rect 28169 11577 28181 11580
rect 28215 11577 28227 11611
rect 28169 11571 28227 11577
rect 23106 11540 23112 11552
rect 22066 11512 23112 11540
rect 20257 11503 20315 11509
rect 23106 11500 23112 11512
rect 23164 11500 23170 11552
rect 23198 11500 23204 11552
rect 23256 11500 23262 11552
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 23937 11543 23995 11549
rect 23937 11540 23949 11543
rect 23532 11512 23949 11540
rect 23532 11500 23538 11512
rect 23937 11509 23949 11512
rect 23983 11509 23995 11543
rect 23937 11503 23995 11509
rect 25590 11500 25596 11552
rect 25648 11540 25654 11552
rect 26329 11543 26387 11549
rect 26329 11540 26341 11543
rect 25648 11512 26341 11540
rect 25648 11500 25654 11512
rect 26329 11509 26341 11512
rect 26375 11509 26387 11543
rect 26329 11503 26387 11509
rect 29362 11500 29368 11552
rect 29420 11540 29426 11552
rect 29549 11543 29607 11549
rect 29549 11540 29561 11543
rect 29420 11512 29561 11540
rect 29420 11500 29426 11512
rect 29549 11509 29561 11512
rect 29595 11509 29607 11543
rect 29549 11503 29607 11509
rect 29914 11500 29920 11552
rect 29972 11500 29978 11552
rect 552 11450 31648 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 12096 11450
rect 12148 11398 12160 11450
rect 12212 11398 12224 11450
rect 12276 11398 12288 11450
rect 12340 11398 12352 11450
rect 12404 11398 19870 11450
rect 19922 11398 19934 11450
rect 19986 11398 19998 11450
rect 20050 11398 20062 11450
rect 20114 11398 20126 11450
rect 20178 11398 27644 11450
rect 27696 11398 27708 11450
rect 27760 11398 27772 11450
rect 27824 11398 27836 11450
rect 27888 11398 27900 11450
rect 27952 11398 31648 11450
rect 552 11376 31648 11398
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 5537 11339 5595 11345
rect 4304 11308 4752 11336
rect 4304 11296 4310 11308
rect 2682 11228 2688 11280
rect 2740 11268 2746 11280
rect 2740 11240 4292 11268
rect 2740 11228 2746 11240
rect 1210 11160 1216 11212
rect 1268 11200 1274 11212
rect 1857 11203 1915 11209
rect 1857 11200 1869 11203
rect 1268 11172 1869 11200
rect 1268 11160 1274 11172
rect 1857 11169 1869 11172
rect 1903 11169 1915 11203
rect 1857 11163 1915 11169
rect 2124 11203 2182 11209
rect 2124 11169 2136 11203
rect 2170 11200 2182 11203
rect 2406 11200 2412 11212
rect 2170 11172 2412 11200
rect 2170 11169 2182 11172
rect 2124 11163 2182 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 4264 11209 4292 11240
rect 4724 11209 4752 11308
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 5902 11336 5908 11348
rect 5583 11308 5908 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 5902 11296 5908 11308
rect 5960 11296 5966 11348
rect 8754 11296 8760 11348
rect 8812 11296 8818 11348
rect 10042 11336 10048 11348
rect 9048 11308 10048 11336
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11169 4307 11203
rect 4249 11163 4307 11169
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11169 4767 11203
rect 4709 11163 4767 11169
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5534 11200 5540 11212
rect 5399 11172 5540 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 5813 11203 5871 11209
rect 5813 11200 5825 11203
rect 5675 11172 5825 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5813 11169 5825 11172
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 5997 11203 6055 11209
rect 5997 11169 6009 11203
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 3881 11135 3939 11141
rect 3881 11132 3893 11135
rect 3436 11104 3893 11132
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 3329 11067 3387 11073
rect 3329 11064 3341 11067
rect 2924 11036 3341 11064
rect 2924 11024 2930 11036
rect 3329 11033 3341 11036
rect 3375 11033 3387 11067
rect 3329 11027 3387 11033
rect 3237 10999 3295 11005
rect 3237 10965 3249 10999
rect 3283 10996 3295 10999
rect 3436 10996 3464 11104
rect 3881 11101 3893 11104
rect 3927 11132 3939 11135
rect 4154 11132 4160 11144
rect 3927 11104 4160 11132
rect 3927 11101 3939 11104
rect 3881 11095 3939 11101
rect 4154 11092 4160 11104
rect 4212 11132 4218 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4212 11104 4445 11132
rect 4212 11092 4218 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 5718 11132 5724 11144
rect 4847 11104 5724 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 5718 11092 5724 11104
rect 5776 11132 5782 11144
rect 6012 11132 6040 11163
rect 6086 11160 6092 11212
rect 6144 11160 6150 11212
rect 6362 11160 6368 11212
rect 6420 11160 6426 11212
rect 9048 11209 9076 11308
rect 10042 11296 10048 11308
rect 10100 11336 10106 11348
rect 14918 11336 14924 11348
rect 10100 11308 14924 11336
rect 10100 11296 10106 11308
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 15562 11296 15568 11348
rect 15620 11296 15626 11348
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19153 11339 19211 11345
rect 19153 11336 19165 11339
rect 19116 11308 19165 11336
rect 19116 11296 19122 11308
rect 19153 11305 19165 11308
rect 19199 11305 19211 11339
rect 19518 11336 19524 11348
rect 19153 11299 19211 11305
rect 19352 11308 19524 11336
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 9677 11271 9735 11277
rect 9677 11268 9689 11271
rect 9364 11240 9689 11268
rect 9364 11228 9370 11240
rect 9677 11237 9689 11240
rect 9723 11237 9735 11271
rect 9677 11231 9735 11237
rect 12406 11240 17264 11268
rect 9033 11203 9091 11209
rect 9033 11169 9045 11203
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9122 11160 9128 11212
rect 9180 11160 9186 11212
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11169 9275 11203
rect 9217 11163 9275 11169
rect 5776 11104 6040 11132
rect 5776 11092 5782 11104
rect 6270 11092 6276 11144
rect 6328 11092 6334 11144
rect 9232 11132 9260 11163
rect 9398 11160 9404 11212
rect 9456 11160 9462 11212
rect 9858 11160 9864 11212
rect 9916 11160 9922 11212
rect 9493 11135 9551 11141
rect 9493 11132 9505 11135
rect 9232 11104 9505 11132
rect 9493 11101 9505 11104
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 5169 11067 5227 11073
rect 5169 11064 5181 11067
rect 4948 11036 5181 11064
rect 4948 11024 4954 11036
rect 5169 11033 5181 11036
rect 5215 11033 5227 11067
rect 5169 11027 5227 11033
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 12406 11064 12434 11240
rect 15838 11160 15844 11212
rect 15896 11160 15902 11212
rect 16390 11160 16396 11212
rect 16448 11160 16454 11212
rect 15746 11132 15752 11144
rect 5316 11036 12434 11064
rect 15212 11104 15752 11132
rect 5316 11024 5322 11036
rect 3283 10968 3464 10996
rect 3283 10965 3295 10968
rect 3237 10959 3295 10965
rect 4062 10956 4068 11008
rect 4120 10956 4126 11008
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 9950 10996 9956 11008
rect 4856 10968 9956 10996
rect 4856 10956 4862 10968
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 15212 10996 15240 11104
rect 15746 11092 15752 11104
rect 15804 11132 15810 11144
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 15804 11104 16221 11132
rect 15804 11092 15810 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 17236 11132 17264 11240
rect 19352 11209 19380 11308
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 20530 11296 20536 11348
rect 20588 11296 20594 11348
rect 21726 11296 21732 11348
rect 21784 11336 21790 11348
rect 21913 11339 21971 11345
rect 21913 11336 21925 11339
rect 21784 11308 21925 11336
rect 21784 11296 21790 11308
rect 21913 11305 21925 11308
rect 21959 11305 21971 11339
rect 21913 11299 21971 11305
rect 25314 11296 25320 11348
rect 25372 11296 25378 11348
rect 25866 11296 25872 11348
rect 25924 11296 25930 11348
rect 26237 11339 26295 11345
rect 26237 11305 26249 11339
rect 26283 11336 26295 11339
rect 26602 11336 26608 11348
rect 26283 11308 26608 11336
rect 26283 11305 26295 11308
rect 26237 11299 26295 11305
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 27338 11296 27344 11348
rect 27396 11336 27402 11348
rect 27801 11339 27859 11345
rect 27801 11336 27813 11339
rect 27396 11308 27813 11336
rect 27396 11296 27402 11308
rect 27801 11305 27813 11308
rect 27847 11305 27859 11339
rect 29914 11336 29920 11348
rect 27801 11299 27859 11305
rect 29012 11308 29920 11336
rect 19659 11271 19717 11277
rect 19659 11237 19671 11271
rect 19705 11268 19717 11271
rect 20548 11268 20576 11296
rect 19705 11240 20576 11268
rect 19705 11237 19717 11240
rect 19659 11231 19717 11237
rect 23198 11228 23204 11280
rect 23256 11277 23262 11280
rect 23256 11268 23268 11277
rect 25685 11271 25743 11277
rect 23256 11240 23301 11268
rect 23256 11231 23268 11240
rect 25685 11237 25697 11271
rect 25731 11268 25743 11271
rect 25884 11268 25912 11296
rect 26694 11277 26700 11280
rect 26688 11268 26700 11277
rect 25731 11240 25912 11268
rect 26068 11240 26556 11268
rect 26655 11240 26700 11268
rect 25731 11237 25743 11240
rect 25685 11231 25743 11237
rect 23256 11228 23262 11231
rect 26068 11212 26096 11240
rect 19337 11203 19395 11209
rect 19337 11169 19349 11203
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 19426 11160 19432 11212
rect 19484 11160 19490 11212
rect 19521 11203 19579 11209
rect 19521 11169 19533 11203
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 19797 11203 19855 11209
rect 19797 11169 19809 11203
rect 19843 11200 19855 11203
rect 19978 11200 19984 11212
rect 19843 11172 19984 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 19536 11132 19564 11163
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20070 11160 20076 11212
rect 20128 11160 20134 11212
rect 20162 11160 20168 11212
rect 20220 11160 20226 11212
rect 20254 11160 20260 11212
rect 20312 11160 20318 11212
rect 20346 11160 20352 11212
rect 20404 11209 20410 11212
rect 20404 11203 20433 11209
rect 20421 11169 20433 11203
rect 20404 11163 20433 11169
rect 20404 11160 20410 11163
rect 21174 11160 21180 11212
rect 21232 11200 21238 11212
rect 22005 11203 22063 11209
rect 22005 11200 22017 11203
rect 21232 11172 22017 11200
rect 21232 11160 21238 11172
rect 22005 11169 22017 11172
rect 22051 11169 22063 11203
rect 22005 11163 22063 11169
rect 23474 11160 23480 11212
rect 23532 11160 23538 11212
rect 24026 11160 24032 11212
rect 24084 11200 24090 11212
rect 25498 11200 25504 11212
rect 24084 11172 25504 11200
rect 24084 11160 24090 11172
rect 25498 11160 25504 11172
rect 25556 11160 25562 11212
rect 25590 11160 25596 11212
rect 25648 11160 25654 11212
rect 25774 11160 25780 11212
rect 25832 11209 25838 11212
rect 25832 11203 25861 11209
rect 25849 11169 25861 11203
rect 25832 11163 25861 11169
rect 25832 11160 25838 11163
rect 25958 11160 25964 11212
rect 26016 11160 26022 11212
rect 26050 11160 26056 11212
rect 26108 11160 26114 11212
rect 26234 11160 26240 11212
rect 26292 11160 26298 11212
rect 26418 11160 26424 11212
rect 26476 11160 26482 11212
rect 26528 11200 26556 11240
rect 26688 11231 26700 11240
rect 26694 11228 26700 11231
rect 26752 11228 26758 11280
rect 26528 11172 28580 11200
rect 20272 11132 20300 11160
rect 17236 11104 19334 11132
rect 19536 11104 20300 11132
rect 16209 11095 16267 11101
rect 19306 11076 19334 11104
rect 20530 11092 20536 11144
rect 20588 11092 20594 11144
rect 28552 11132 28580 11172
rect 28626 11160 28632 11212
rect 28684 11160 28690 11212
rect 28810 11160 28816 11212
rect 28868 11160 28874 11212
rect 29012 11209 29040 11308
rect 29914 11296 29920 11308
rect 29972 11296 29978 11348
rect 29273 11271 29331 11277
rect 29273 11237 29285 11271
rect 29319 11268 29331 11271
rect 29610 11271 29668 11277
rect 29610 11268 29622 11271
rect 29319 11240 29622 11268
rect 29319 11237 29331 11240
rect 29273 11231 29331 11237
rect 29610 11237 29622 11240
rect 29656 11237 29668 11271
rect 29610 11231 29668 11237
rect 28905 11203 28963 11209
rect 28905 11169 28917 11203
rect 28951 11169 28963 11203
rect 28905 11163 28963 11169
rect 28997 11203 29055 11209
rect 28997 11169 29009 11203
rect 29043 11169 29055 11203
rect 28997 11163 29055 11169
rect 28920 11132 28948 11163
rect 29362 11160 29368 11212
rect 29420 11160 29426 11212
rect 29086 11132 29092 11144
rect 28552 11104 29092 11132
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 19306 11036 19340 11076
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 20898 11064 20904 11076
rect 20220 11036 20904 11064
rect 20220 11024 20226 11036
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 22097 11067 22155 11073
rect 22097 11033 22109 11067
rect 22143 11064 22155 11067
rect 22462 11064 22468 11076
rect 22143 11036 22468 11064
rect 22143 11033 22155 11036
rect 22097 11027 22155 11033
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 29178 11064 29184 11076
rect 28966 11036 29184 11064
rect 14332 10968 15240 10996
rect 14332 10956 14338 10968
rect 16574 10956 16580 11008
rect 16632 10956 16638 11008
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 17586 10996 17592 11008
rect 16908 10968 17592 10996
rect 16908 10956 16914 10968
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 19610 10956 19616 11008
rect 19668 10996 19674 11008
rect 19889 10999 19947 11005
rect 19889 10996 19901 10999
rect 19668 10968 19901 10996
rect 19668 10956 19674 10968
rect 19889 10965 19901 10968
rect 19935 10965 19947 10999
rect 19889 10959 19947 10965
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 28966 10996 28994 11036
rect 29178 11024 29184 11036
rect 29236 11024 29242 11076
rect 30745 11067 30803 11073
rect 30745 11033 30757 11067
rect 30791 11064 30803 11067
rect 30834 11064 30840 11076
rect 30791 11036 30840 11064
rect 30791 11033 30803 11036
rect 30745 11027 30803 11033
rect 30834 11024 30840 11036
rect 30892 11024 30898 11076
rect 20036 10968 28994 10996
rect 20036 10956 20042 10968
rect 552 10906 31648 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 11436 10906
rect 11488 10854 11500 10906
rect 11552 10854 11564 10906
rect 11616 10854 11628 10906
rect 11680 10854 11692 10906
rect 11744 10854 19210 10906
rect 19262 10854 19274 10906
rect 19326 10854 19338 10906
rect 19390 10854 19402 10906
rect 19454 10854 19466 10906
rect 19518 10854 26984 10906
rect 27036 10854 27048 10906
rect 27100 10854 27112 10906
rect 27164 10854 27176 10906
rect 27228 10854 27240 10906
rect 27292 10854 31648 10906
rect 552 10832 31648 10854
rect 2406 10752 2412 10804
rect 2464 10752 2470 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5592 10764 5641 10792
rect 5592 10752 5598 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 9858 10792 9864 10804
rect 5629 10755 5687 10761
rect 7852 10764 9864 10792
rect 2774 10724 2780 10736
rect 2240 10696 2780 10724
rect 2240 10597 2268 10696
rect 2774 10684 2780 10696
rect 2832 10724 2838 10736
rect 3326 10724 3332 10736
rect 2832 10696 3332 10724
rect 2832 10684 2838 10696
rect 3326 10684 3332 10696
rect 3384 10724 3390 10736
rect 4062 10724 4068 10736
rect 3384 10696 4068 10724
rect 3384 10684 3390 10696
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 7852 10668 7880 10764
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10008 10764 15792 10792
rect 10008 10752 10014 10764
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 9122 10724 9128 10736
rect 8812 10696 9128 10724
rect 8812 10684 8818 10696
rect 9122 10684 9128 10696
rect 9180 10684 9186 10736
rect 15764 10724 15792 10764
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15896 10764 16037 10792
rect 15896 10752 15902 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 16482 10792 16488 10804
rect 16025 10755 16083 10761
rect 16132 10764 16488 10792
rect 16132 10724 16160 10764
rect 16482 10752 16488 10764
rect 16540 10792 16546 10804
rect 16540 10764 20852 10792
rect 16540 10752 16546 10764
rect 15764 10696 16160 10724
rect 20824 10724 20852 10764
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 22428 10764 26740 10792
rect 22428 10752 22434 10764
rect 26421 10727 26479 10733
rect 26421 10724 26433 10727
rect 20824 10696 26433 10724
rect 26421 10693 26433 10696
rect 26467 10724 26479 10727
rect 26510 10724 26516 10736
rect 26467 10696 26516 10724
rect 26467 10693 26479 10696
rect 26421 10687 26479 10693
rect 26510 10684 26516 10696
rect 26568 10684 26574 10736
rect 26712 10724 26740 10764
rect 26786 10752 26792 10804
rect 26844 10792 26850 10804
rect 26881 10795 26939 10801
rect 26881 10792 26893 10795
rect 26844 10764 26893 10792
rect 26844 10752 26850 10764
rect 26881 10761 26893 10764
rect 26927 10761 26939 10795
rect 26881 10755 26939 10761
rect 28810 10752 28816 10804
rect 28868 10792 28874 10804
rect 29181 10795 29239 10801
rect 29181 10792 29193 10795
rect 28868 10764 29193 10792
rect 28868 10752 28874 10764
rect 29181 10761 29193 10764
rect 29227 10761 29239 10795
rect 29181 10755 29239 10761
rect 27154 10724 27160 10736
rect 26712 10696 27160 10724
rect 27154 10684 27160 10696
rect 27212 10724 27218 10736
rect 28074 10724 28080 10736
rect 27212 10696 28080 10724
rect 27212 10684 27218 10696
rect 28074 10684 28080 10696
rect 28132 10684 28138 10736
rect 30834 10724 30840 10736
rect 29012 10696 30840 10724
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2424 10628 2697 10656
rect 2424 10597 2452 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 6270 10656 6276 10668
rect 4571 10628 6276 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 2590 10548 2596 10600
rect 2648 10548 2654 10600
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 2866 10588 2872 10600
rect 2823 10560 2872 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3200 10560 3433 10588
rect 3200 10548 3206 10560
rect 3421 10557 3433 10560
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 6012 10597 6040 10628
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7834 10656 7840 10668
rect 7156 10628 7840 10656
rect 7156 10616 7162 10628
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 18877 10659 18935 10665
rect 8588 10628 11100 10656
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 4212 10560 4445 10588
rect 4212 10548 4218 10560
rect 4433 10557 4445 10560
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6362 10588 6368 10600
rect 6227 10560 6368 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 5828 10520 5856 10551
rect 6362 10548 6368 10560
rect 6420 10588 6426 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 6420 10560 8033 10588
rect 6420 10548 6426 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8588 10588 8616 10628
rect 8021 10551 8079 10557
rect 8128 10560 8616 10588
rect 3344 10492 5856 10520
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 3344 10461 3372 10492
rect 3329 10455 3387 10461
rect 3329 10452 3341 10455
rect 2188 10424 3341 10452
rect 2188 10412 2194 10424
rect 3329 10421 3341 10424
rect 3375 10421 3387 10455
rect 5828 10452 5856 10492
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 6086 10520 6092 10532
rect 5951 10492 6092 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 6086 10480 6092 10492
rect 6144 10520 6150 10532
rect 6144 10492 7788 10520
rect 6144 10480 6150 10492
rect 5994 10452 6000 10464
rect 5828 10424 6000 10452
rect 3329 10415 3387 10421
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 7760 10452 7788 10492
rect 7834 10480 7840 10532
rect 7892 10480 7898 10532
rect 8128 10452 8156 10560
rect 8662 10548 8668 10600
rect 8720 10548 8726 10600
rect 8754 10548 8760 10600
rect 8812 10548 8818 10600
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 8205 10523 8263 10529
rect 8205 10489 8217 10523
rect 8251 10520 8263 10523
rect 8864 10520 8892 10551
rect 9030 10548 9036 10600
rect 9088 10548 9094 10600
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 9916 10560 10241 10588
rect 9916 10548 9922 10560
rect 10229 10557 10241 10560
rect 10275 10588 10287 10591
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10275 10560 10885 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 8251 10492 8892 10520
rect 9048 10520 9076 10548
rect 9490 10520 9496 10532
rect 9048 10492 9496 10520
rect 8251 10489 8263 10492
rect 8205 10483 8263 10489
rect 9490 10480 9496 10492
rect 9548 10480 9554 10532
rect 10410 10480 10416 10532
rect 10468 10480 10474 10532
rect 11072 10529 11100 10628
rect 16040 10628 16252 10656
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12759 10560 12909 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 12897 10557 12909 10560
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 13722 10588 13728 10600
rect 13035 10560 13728 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 14274 10548 14280 10600
rect 14332 10548 14338 10600
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 11057 10523 11115 10529
rect 11057 10489 11069 10523
rect 11103 10520 11115 10523
rect 11103 10492 11376 10520
rect 11103 10489 11115 10492
rect 11057 10483 11115 10489
rect 7760 10424 8156 10452
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 8754 10412 8760 10464
rect 8812 10452 8818 10464
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 8812 10424 9229 10452
rect 8812 10412 8818 10424
rect 9217 10421 9229 10424
rect 9263 10421 9275 10455
rect 9217 10415 9275 10421
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 11238 10412 11244 10464
rect 11296 10412 11302 10464
rect 11348 10461 11376 10492
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12446 10523 12504 10529
rect 12446 10520 12458 10523
rect 12032 10492 12458 10520
rect 12032 10480 12038 10492
rect 12446 10489 12458 10492
rect 12492 10489 12504 10523
rect 12446 10483 12504 10489
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 13446 10520 13452 10532
rect 13136 10492 13452 10520
rect 13136 10480 13142 10492
rect 13446 10480 13452 10492
rect 13504 10520 13510 10532
rect 14384 10520 14412 10551
rect 14642 10548 14648 10600
rect 14700 10548 14706 10600
rect 15194 10548 15200 10600
rect 15252 10588 15258 10600
rect 16040 10588 16068 10628
rect 15252 10560 16068 10588
rect 15252 10548 15258 10560
rect 16114 10548 16120 10600
rect 16172 10548 16178 10600
rect 16224 10588 16252 10628
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 18923 10628 19533 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 24210 10616 24216 10668
rect 24268 10656 24274 10668
rect 24489 10659 24547 10665
rect 24489 10656 24501 10659
rect 24268 10628 24501 10656
rect 24268 10616 24274 10628
rect 24489 10625 24501 10628
rect 24535 10625 24547 10659
rect 24489 10619 24547 10625
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 24912 10628 25636 10656
rect 24912 10616 24918 10628
rect 17678 10588 17684 10600
rect 16224 10560 17684 10588
rect 17678 10548 17684 10560
rect 17736 10588 17742 10600
rect 17736 10560 18000 10588
rect 17736 10548 17742 10560
rect 13504 10492 14412 10520
rect 14912 10523 14970 10529
rect 13504 10480 13510 10492
rect 14912 10489 14924 10523
rect 14958 10520 14970 10523
rect 16384 10523 16442 10529
rect 14958 10492 16344 10520
rect 14958 10489 14970 10492
rect 14912 10483 14970 10489
rect 11333 10455 11391 10461
rect 11333 10421 11345 10455
rect 11379 10421 11391 10455
rect 11333 10415 11391 10421
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 13228 10424 13645 10452
rect 13228 10412 13234 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 13633 10415 13691 10421
rect 14550 10412 14556 10464
rect 14608 10412 14614 10464
rect 16316 10452 16344 10492
rect 16384 10489 16396 10523
rect 16430 10520 16442 10523
rect 16574 10520 16580 10532
rect 16430 10492 16580 10520
rect 16430 10489 16442 10492
rect 16384 10483 16442 10489
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 16758 10480 16764 10532
rect 16816 10520 16822 10532
rect 17972 10520 18000 10560
rect 18782 10548 18788 10600
rect 18840 10548 18846 10600
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19061 10591 19119 10597
rect 19061 10588 19073 10591
rect 19024 10560 19073 10588
rect 19024 10548 19030 10560
rect 19061 10557 19073 10560
rect 19107 10557 19119 10591
rect 19061 10551 19119 10557
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10588 19303 10591
rect 19610 10588 19616 10600
rect 19291 10560 19616 10588
rect 19291 10557 19303 10560
rect 19245 10551 19303 10557
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 21174 10548 21180 10600
rect 21232 10548 21238 10600
rect 24026 10548 24032 10600
rect 24084 10548 24090 10600
rect 25130 10548 25136 10600
rect 25188 10588 25194 10600
rect 25608 10597 25636 10628
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 25188 10560 25237 10588
rect 25188 10548 25194 10560
rect 25225 10557 25237 10560
rect 25271 10557 25283 10591
rect 25225 10551 25283 10557
rect 25593 10591 25651 10597
rect 25593 10557 25605 10591
rect 25639 10557 25651 10591
rect 25593 10551 25651 10557
rect 26326 10548 26332 10600
rect 26384 10588 26390 10600
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26384 10560 26985 10588
rect 26384 10548 26390 10560
rect 26973 10557 26985 10560
rect 27019 10588 27031 10591
rect 27338 10588 27344 10600
rect 27019 10560 27344 10588
rect 27019 10557 27031 10560
rect 26973 10551 27031 10557
rect 27338 10548 27344 10560
rect 27396 10548 27402 10600
rect 29012 10588 29040 10696
rect 30834 10684 30840 10696
rect 30892 10684 30898 10736
rect 29178 10616 29184 10668
rect 29236 10656 29242 10668
rect 29236 10628 29868 10656
rect 29236 10616 29242 10628
rect 28920 10560 29040 10588
rect 18322 10520 18328 10532
rect 16816 10492 17540 10520
rect 17972 10492 18328 10520
rect 16816 10480 16822 10492
rect 17512 10464 17540 10492
rect 18322 10480 18328 10492
rect 18380 10480 18386 10532
rect 19429 10523 19487 10529
rect 19429 10489 19441 10523
rect 19475 10520 19487 10523
rect 19766 10523 19824 10529
rect 19766 10520 19778 10523
rect 19475 10492 19778 10520
rect 19475 10489 19487 10492
rect 19429 10483 19487 10489
rect 19766 10489 19778 10492
rect 19812 10489 19824 10523
rect 19766 10483 19824 10489
rect 24121 10523 24179 10529
rect 24121 10489 24133 10523
rect 24167 10489 24179 10523
rect 24121 10483 24179 10489
rect 24213 10523 24271 10529
rect 24213 10489 24225 10523
rect 24259 10489 24271 10523
rect 24213 10483 24271 10489
rect 24351 10523 24409 10529
rect 24351 10489 24363 10523
rect 24397 10520 24409 10523
rect 25774 10520 25780 10532
rect 24397 10492 25780 10520
rect 24397 10489 24409 10492
rect 24351 10483 24409 10489
rect 17218 10452 17224 10464
rect 16316 10424 17224 10452
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 17494 10412 17500 10464
rect 17552 10412 17558 10464
rect 18340 10452 18368 10480
rect 19886 10452 19892 10464
rect 18340 10424 19892 10452
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 21082 10412 21088 10464
rect 21140 10412 21146 10464
rect 23845 10455 23903 10461
rect 23845 10421 23857 10455
rect 23891 10452 23903 10455
rect 23934 10452 23940 10464
rect 23891 10424 23940 10452
rect 23891 10421 23903 10424
rect 23845 10415 23903 10421
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 24026 10412 24032 10464
rect 24084 10452 24090 10464
rect 24136 10452 24164 10483
rect 24084 10424 24164 10452
rect 24228 10452 24256 10483
rect 25774 10480 25780 10492
rect 25832 10520 25838 10532
rect 26234 10520 26240 10532
rect 25832 10492 26240 10520
rect 25832 10480 25838 10492
rect 26234 10480 26240 10492
rect 26292 10480 26298 10532
rect 26605 10523 26663 10529
rect 26605 10489 26617 10523
rect 26651 10520 26663 10523
rect 28920 10520 28948 10560
rect 29086 10548 29092 10600
rect 29144 10548 29150 10600
rect 29270 10548 29276 10600
rect 29328 10588 29334 10600
rect 29840 10597 29868 10628
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29328 10560 29745 10588
rect 29328 10548 29334 10560
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 29825 10591 29883 10597
rect 29825 10557 29837 10591
rect 29871 10557 29883 10591
rect 29825 10551 29883 10557
rect 29917 10591 29975 10597
rect 29917 10557 29929 10591
rect 29963 10557 29975 10591
rect 29917 10551 29975 10557
rect 29932 10520 29960 10551
rect 30098 10548 30104 10600
rect 30156 10548 30162 10600
rect 30282 10548 30288 10600
rect 30340 10588 30346 10600
rect 30745 10591 30803 10597
rect 30745 10588 30757 10591
rect 30340 10560 30757 10588
rect 30340 10548 30346 10560
rect 30745 10557 30757 10560
rect 30791 10557 30803 10591
rect 30745 10551 30803 10557
rect 26651 10492 28948 10520
rect 29840 10492 29960 10520
rect 26651 10489 26663 10492
rect 26605 10483 26663 10489
rect 24673 10455 24731 10461
rect 24673 10452 24685 10455
rect 24228 10424 24685 10452
rect 24084 10412 24090 10424
rect 24673 10421 24685 10424
rect 24719 10421 24731 10455
rect 24673 10415 24731 10421
rect 25498 10412 25504 10464
rect 25556 10412 25562 10464
rect 26694 10412 26700 10464
rect 26752 10452 26758 10464
rect 27982 10452 27988 10464
rect 26752 10424 27988 10452
rect 26752 10412 26758 10424
rect 27982 10412 27988 10424
rect 28040 10412 28046 10464
rect 28626 10412 28632 10464
rect 28684 10452 28690 10464
rect 29840 10452 29868 10492
rect 28684 10424 29868 10452
rect 28684 10412 28690 10424
rect 30006 10412 30012 10464
rect 30064 10412 30070 10464
rect 30742 10412 30748 10464
rect 30800 10452 30806 10464
rect 30837 10455 30895 10461
rect 30837 10452 30849 10455
rect 30800 10424 30849 10452
rect 30800 10412 30806 10424
rect 30837 10421 30849 10424
rect 30883 10421 30895 10455
rect 30837 10415 30895 10421
rect 552 10362 31648 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 12096 10362
rect 12148 10310 12160 10362
rect 12212 10310 12224 10362
rect 12276 10310 12288 10362
rect 12340 10310 12352 10362
rect 12404 10310 19870 10362
rect 19922 10310 19934 10362
rect 19986 10310 19998 10362
rect 20050 10310 20062 10362
rect 20114 10310 20126 10362
rect 20178 10310 27644 10362
rect 27696 10310 27708 10362
rect 27760 10310 27772 10362
rect 27824 10310 27836 10362
rect 27888 10310 27900 10362
rect 27952 10310 31648 10362
rect 552 10288 31648 10310
rect 2774 10248 2780 10260
rect 2746 10208 2780 10248
rect 2832 10208 2838 10260
rect 3142 10208 3148 10260
rect 3200 10208 3206 10260
rect 5074 10208 5080 10260
rect 5132 10208 5138 10260
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 7377 10251 7435 10257
rect 7377 10248 7389 10251
rect 6420 10220 7389 10248
rect 6420 10208 6426 10220
rect 7377 10217 7389 10220
rect 7423 10217 7435 10251
rect 7377 10211 7435 10217
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 8202 10248 8208 10260
rect 7984 10220 8208 10248
rect 7984 10208 7990 10220
rect 8202 10208 8208 10220
rect 8260 10248 8266 10260
rect 9030 10248 9036 10260
rect 8260 10220 9036 10248
rect 8260 10208 8266 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9122 10208 9128 10260
rect 9180 10248 9186 10260
rect 11882 10248 11888 10260
rect 9180 10220 9260 10248
rect 9180 10208 9186 10220
rect 2746 10180 2774 10208
rect 2608 10152 2774 10180
rect 2130 10072 2136 10124
rect 2188 10072 2194 10124
rect 2608 10121 2636 10152
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 5353 10183 5411 10189
rect 3568 10152 4660 10180
rect 3568 10140 3574 10152
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10081 2651 10115
rect 2593 10075 2651 10081
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 2774 10112 2780 10124
rect 2731 10084 2780 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2608 10044 2636 10075
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 4632 10121 4660 10152
rect 5353 10149 5365 10183
rect 5399 10180 5411 10183
rect 6822 10180 6828 10192
rect 5399 10152 6828 10180
rect 5399 10149 5411 10152
rect 5353 10143 5411 10149
rect 6822 10140 6828 10152
rect 6880 10140 6886 10192
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 8490 10183 8548 10189
rect 8490 10180 8502 10183
rect 8444 10152 8502 10180
rect 8444 10140 8450 10152
rect 8490 10149 8502 10152
rect 8536 10149 8548 10183
rect 8490 10143 8548 10149
rect 9232 10180 9260 10220
rect 10428 10220 11888 10248
rect 9232 10152 9812 10180
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 3881 10115 3939 10121
rect 3881 10112 3893 10115
rect 2915 10084 3893 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3881 10081 3893 10084
rect 3927 10081 3939 10115
rect 3881 10075 3939 10081
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10081 4675 10115
rect 4617 10075 4675 10081
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 4982 10112 4988 10124
rect 4847 10084 4988 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 2271 10016 2636 10044
rect 2792 10044 2820 10072
rect 3697 10047 3755 10053
rect 3697 10044 3709 10047
rect 2792 10016 3709 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 3697 10013 3709 10016
rect 3743 10013 3755 10047
rect 3697 10007 3755 10013
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4304 10016 4445 10044
rect 4304 10004 4310 10016
rect 4433 10013 4445 10016
rect 4479 10044 4491 10047
rect 5074 10044 5080 10056
rect 4479 10016 5080 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5276 10044 5304 10075
rect 5442 10072 5448 10124
rect 5500 10072 5506 10124
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 5902 10112 5908 10124
rect 5675 10084 5908 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 5994 10072 6000 10124
rect 6052 10072 6058 10124
rect 6086 10072 6092 10124
rect 6144 10072 6150 10124
rect 6362 10072 6368 10124
rect 6420 10072 6426 10124
rect 8754 10072 8760 10124
rect 8812 10072 8818 10124
rect 8938 10072 8944 10124
rect 8996 10112 9002 10124
rect 9232 10121 9260 10152
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8996 10084 9137 10112
rect 8996 10072 9002 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9398 10112 9404 10124
rect 9355 10084 9404 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 5718 10044 5724 10056
rect 5276 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 9140 10044 9168 10075
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9490 10072 9496 10124
rect 9548 10072 9554 10124
rect 9674 10044 9680 10056
rect 9140 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 9784 10044 9812 10152
rect 10428 10121 10456 10220
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 11974 10208 11980 10260
rect 12032 10208 12038 10260
rect 14642 10208 14648 10260
rect 14700 10248 14706 10260
rect 14829 10251 14887 10257
rect 14829 10248 14841 10251
rect 14700 10220 14841 10248
rect 14700 10208 14706 10220
rect 14829 10217 14841 10220
rect 14875 10217 14887 10251
rect 14829 10211 14887 10217
rect 15841 10251 15899 10257
rect 15841 10217 15853 10251
rect 15887 10248 15899 10251
rect 15930 10248 15936 10260
rect 15887 10220 15936 10248
rect 15887 10217 15899 10220
rect 15841 10211 15899 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 16172 10220 16313 10248
rect 16172 10208 16178 10220
rect 16301 10217 16313 10220
rect 16347 10217 16359 10251
rect 16301 10211 16359 10217
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16485 10251 16543 10257
rect 16485 10248 16497 10251
rect 16448 10220 16497 10248
rect 16448 10208 16454 10220
rect 16485 10217 16497 10220
rect 16531 10217 16543 10251
rect 16485 10211 16543 10217
rect 17218 10208 17224 10260
rect 17276 10208 17282 10260
rect 20346 10248 20352 10260
rect 19306 10220 20352 10248
rect 11146 10180 11152 10192
rect 10520 10152 11152 10180
rect 10520 10121 10548 10152
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 11238 10140 11244 10192
rect 11296 10180 11302 10192
rect 11296 10152 11560 10180
rect 11296 10140 11302 10152
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10520 10044 10548 10075
rect 10594 10072 10600 10124
rect 10652 10072 10658 10124
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10112 10839 10115
rect 11330 10112 11336 10124
rect 10827 10084 11336 10112
rect 10827 10081 10839 10084
rect 10781 10075 10839 10081
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 11532 10121 11560 10152
rect 13630 10140 13636 10192
rect 13688 10180 13694 10192
rect 13688 10152 15056 10180
rect 13688 10140 13694 10152
rect 15028 10124 15056 10152
rect 16040 10152 16436 10180
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 11609 10115 11667 10121
rect 11609 10081 11621 10115
rect 11655 10081 11667 10115
rect 11609 10075 11667 10081
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10112 11759 10115
rect 13078 10112 13084 10124
rect 11747 10084 13084 10112
rect 11747 10081 11759 10084
rect 11701 10075 11759 10081
rect 9784 10016 10548 10044
rect 11422 10004 11428 10056
rect 11480 10044 11486 10056
rect 11624 10044 11652 10075
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13170 10072 13176 10124
rect 13228 10072 13234 10124
rect 13446 10121 13452 10124
rect 13440 10075 13452 10121
rect 13446 10072 13452 10075
rect 13504 10072 13510 10124
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 14921 10115 14979 10121
rect 14921 10112 14933 10115
rect 13780 10084 14933 10112
rect 13780 10072 13786 10084
rect 14921 10081 14933 10084
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 11480 10016 11652 10044
rect 14936 10044 14964 10075
rect 15010 10072 15016 10124
rect 15068 10072 15074 10124
rect 15194 10072 15200 10124
rect 15252 10072 15258 10124
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 15746 10112 15752 10124
rect 15703 10084 15752 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 15933 10118 15991 10121
rect 16040 10118 16068 10152
rect 16408 10124 16436 10152
rect 16758 10140 16764 10192
rect 16816 10140 16822 10192
rect 16850 10140 16856 10192
rect 16908 10140 16914 10192
rect 16942 10140 16948 10192
rect 17000 10189 17006 10192
rect 17000 10183 17029 10189
rect 17017 10180 17029 10183
rect 17017 10152 17264 10180
rect 17017 10149 17029 10152
rect 17000 10143 17029 10149
rect 17000 10140 17006 10143
rect 15933 10115 16068 10118
rect 15933 10081 15945 10115
rect 15979 10090 16068 10115
rect 16209 10115 16267 10121
rect 15979 10081 15991 10090
rect 15933 10075 15991 10081
rect 16209 10081 16221 10115
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 16224 10044 16252 10075
rect 16390 10072 16396 10124
rect 16448 10072 16454 10124
rect 16666 10072 16672 10124
rect 16724 10072 16730 10124
rect 17126 10072 17132 10124
rect 17184 10072 17190 10124
rect 17236 10112 17264 10152
rect 17310 10140 17316 10192
rect 17368 10189 17374 10192
rect 17368 10183 17431 10189
rect 17368 10149 17385 10183
rect 17419 10149 17431 10183
rect 17368 10143 17431 10149
rect 17368 10140 17374 10143
rect 17586 10140 17592 10192
rect 17644 10140 17650 10192
rect 19306 10112 19334 10220
rect 20346 10208 20352 10220
rect 20404 10248 20410 10260
rect 20714 10248 20720 10260
rect 20404 10220 20720 10248
rect 20404 10208 20410 10220
rect 20714 10208 20720 10220
rect 20772 10208 20778 10260
rect 27430 10248 27436 10260
rect 26160 10220 27436 10248
rect 21082 10180 21088 10192
rect 19720 10152 21088 10180
rect 19720 10121 19748 10152
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 25498 10180 25504 10192
rect 23676 10152 25504 10180
rect 19978 10121 19984 10124
rect 17236 10084 19334 10112
rect 19705 10115 19763 10121
rect 19705 10081 19717 10115
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 19972 10075 19984 10121
rect 19978 10072 19984 10075
rect 20036 10072 20042 10124
rect 22370 10072 22376 10124
rect 22428 10072 22434 10124
rect 23676 10121 23704 10152
rect 25498 10140 25504 10152
rect 25556 10140 25562 10192
rect 26160 10189 26188 10220
rect 27430 10208 27436 10220
rect 27488 10208 27494 10260
rect 27982 10208 27988 10260
rect 28040 10248 28046 10260
rect 29273 10251 29331 10257
rect 28040 10220 28948 10248
rect 28040 10208 28046 10220
rect 28920 10192 28948 10220
rect 29273 10217 29285 10251
rect 29319 10248 29331 10251
rect 30098 10248 30104 10260
rect 29319 10220 30104 10248
rect 29319 10217 29331 10220
rect 29273 10211 29331 10217
rect 30098 10208 30104 10220
rect 30156 10208 30162 10260
rect 26145 10183 26203 10189
rect 26145 10149 26157 10183
rect 26191 10149 26203 10183
rect 26145 10143 26203 10149
rect 26234 10140 26240 10192
rect 26292 10180 26298 10192
rect 26579 10183 26637 10189
rect 26579 10180 26591 10183
rect 26292 10152 26591 10180
rect 26292 10140 26298 10152
rect 26579 10149 26591 10152
rect 26625 10180 26637 10183
rect 27065 10183 27123 10189
rect 26625 10152 27016 10180
rect 26625 10149 26637 10152
rect 26579 10143 26637 10149
rect 23934 10121 23940 10124
rect 23661 10115 23719 10121
rect 23661 10081 23673 10115
rect 23707 10081 23719 10115
rect 23928 10112 23940 10121
rect 23895 10084 23940 10112
rect 23661 10075 23719 10081
rect 23928 10075 23940 10084
rect 23934 10072 23940 10075
rect 23992 10072 23998 10124
rect 25406 10072 25412 10124
rect 25464 10112 25470 10124
rect 25464 10084 26648 10112
rect 25464 10072 25470 10084
rect 14936 10016 16252 10044
rect 16684 10044 16712 10072
rect 18046 10044 18052 10056
rect 16684 10016 18052 10044
rect 11480 10004 11486 10016
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 21821 10047 21879 10053
rect 21821 10044 21833 10047
rect 21468 10016 21833 10044
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 9030 9976 9036 9988
rect 8812 9948 9036 9976
rect 8812 9936 8818 9948
rect 9030 9936 9036 9948
rect 9088 9976 9094 9988
rect 12802 9976 12808 9988
rect 9088 9948 12808 9976
rect 9088 9936 9094 9948
rect 12802 9936 12808 9948
rect 12860 9936 12866 9988
rect 15289 9979 15347 9985
rect 15289 9945 15301 9979
rect 15335 9945 15347 9979
rect 15289 9939 15347 9945
rect 15473 9979 15531 9985
rect 15473 9945 15485 9979
rect 15519 9976 15531 9979
rect 15519 9948 17448 9976
rect 15519 9945 15531 9948
rect 15473 9939 15531 9945
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9908 1915 9911
rect 1946 9908 1952 9920
rect 1903 9880 1952 9908
rect 1903 9877 1915 9880
rect 1857 9871 1915 9877
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 2866 9868 2872 9920
rect 2924 9868 2930 9920
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4709 9911 4767 9917
rect 4709 9908 4721 9911
rect 4120 9880 4721 9908
rect 4120 9868 4126 9880
rect 4709 9877 4721 9880
rect 4755 9877 4767 9911
rect 4709 9871 4767 9877
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5684 9880 5825 9908
rect 5684 9868 5690 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6273 9911 6331 9917
rect 6273 9908 6285 9911
rect 6052 9880 6285 9908
rect 6052 9868 6058 9880
rect 6273 9877 6285 9880
rect 6319 9877 6331 9911
rect 6273 9871 6331 9877
rect 8846 9868 8852 9920
rect 8904 9868 8910 9920
rect 10134 9868 10140 9920
rect 10192 9868 10198 9920
rect 11330 9868 11336 9920
rect 11388 9908 11394 9920
rect 12066 9908 12072 9920
rect 11388 9880 12072 9908
rect 11388 9868 11394 9880
rect 12066 9868 12072 9880
rect 12124 9908 12130 9920
rect 14274 9908 14280 9920
rect 12124 9880 14280 9908
rect 12124 9868 12130 9880
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9908 14611 9911
rect 15102 9908 15108 9920
rect 14599 9880 15108 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15304 9908 15332 9939
rect 16666 9908 16672 9920
rect 15304 9880 16672 9908
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 17420 9917 17448 9948
rect 20806 9936 20812 9988
rect 20864 9976 20870 9988
rect 21269 9979 21327 9985
rect 21269 9976 21281 9979
rect 20864 9948 21281 9976
rect 20864 9936 20870 9948
rect 21269 9945 21281 9948
rect 21315 9945 21327 9979
rect 21269 9939 21327 9945
rect 21468 9920 21496 10016
rect 21821 10013 21833 10016
rect 21867 10013 21879 10047
rect 21821 10007 21879 10013
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10044 22247 10047
rect 23290 10044 23296 10056
rect 22235 10016 23296 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 23290 10004 23296 10016
rect 23348 10044 23354 10056
rect 26421 10047 26479 10053
rect 23348 10016 23428 10044
rect 23348 10004 23354 10016
rect 23400 9920 23428 10016
rect 26421 10013 26433 10047
rect 26467 10013 26479 10047
rect 26620 10044 26648 10084
rect 26694 10072 26700 10124
rect 26752 10072 26758 10124
rect 26786 10072 26792 10124
rect 26844 10072 26850 10124
rect 26881 10115 26939 10121
rect 26881 10081 26893 10115
rect 26927 10081 26939 10115
rect 26988 10112 27016 10152
rect 27065 10149 27077 10183
rect 27111 10180 27123 10183
rect 28626 10180 28632 10192
rect 27111 10152 28120 10180
rect 27111 10149 27123 10152
rect 27065 10143 27123 10149
rect 27295 10115 27353 10121
rect 27295 10112 27307 10115
rect 26988 10084 27307 10112
rect 26881 10075 26939 10081
rect 27295 10081 27307 10084
rect 27341 10081 27353 10115
rect 27295 10075 27353 10081
rect 26896 10044 26924 10075
rect 27430 10072 27436 10124
rect 27488 10072 27494 10124
rect 27522 10072 27528 10124
rect 27580 10072 27586 10124
rect 28092 10121 28120 10152
rect 28276 10152 28632 10180
rect 28276 10121 28304 10152
rect 28626 10140 28632 10152
rect 28684 10140 28690 10192
rect 28902 10140 28908 10192
rect 28960 10140 28966 10192
rect 28997 10183 29055 10189
rect 28997 10149 29009 10183
rect 29043 10180 29055 10183
rect 29914 10180 29920 10192
rect 29043 10152 29920 10180
rect 29043 10149 29055 10152
rect 28997 10143 29055 10149
rect 29914 10140 29920 10152
rect 29972 10140 29978 10192
rect 30006 10140 30012 10192
rect 30064 10180 30070 10192
rect 30478 10183 30536 10189
rect 30478 10180 30490 10183
rect 30064 10152 30490 10180
rect 30064 10140 30070 10152
rect 30478 10149 30490 10152
rect 30524 10149 30536 10183
rect 30478 10143 30536 10149
rect 27617 10115 27675 10121
rect 27617 10081 27629 10115
rect 27663 10081 27675 10115
rect 27617 10075 27675 10081
rect 28077 10115 28135 10121
rect 28077 10081 28089 10115
rect 28123 10081 28135 10115
rect 28077 10075 28135 10081
rect 28261 10115 28319 10121
rect 28261 10081 28273 10115
rect 28307 10081 28319 10115
rect 28261 10075 28319 10081
rect 26620 10016 27108 10044
rect 26421 10007 26479 10013
rect 24596 9948 25268 9976
rect 17405 9911 17463 9917
rect 17405 9877 17417 9911
rect 17451 9877 17463 9911
rect 17405 9871 17463 9877
rect 21085 9911 21143 9917
rect 21085 9877 21097 9911
rect 21131 9908 21143 9911
rect 21450 9908 21456 9920
rect 21131 9880 21456 9908
rect 21131 9877 21143 9880
rect 21085 9871 21143 9877
rect 21450 9868 21456 9880
rect 21508 9868 21514 9920
rect 22554 9868 22560 9920
rect 22612 9868 22618 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 24596 9908 24624 9948
rect 23440 9880 24624 9908
rect 25041 9911 25099 9917
rect 23440 9868 23446 9880
rect 25041 9877 25053 9911
rect 25087 9908 25099 9911
rect 25130 9908 25136 9920
rect 25087 9880 25136 9908
rect 25087 9877 25099 9880
rect 25041 9871 25099 9877
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 25240 9908 25268 9948
rect 25774 9936 25780 9988
rect 25832 9976 25838 9988
rect 26436 9976 26464 10007
rect 26878 9976 26884 9988
rect 25832 9948 26884 9976
rect 25832 9936 25838 9948
rect 26878 9936 26884 9948
rect 26936 9936 26942 9988
rect 27080 9976 27108 10016
rect 27154 10004 27160 10056
rect 27212 10004 27218 10056
rect 27632 9976 27660 10075
rect 28442 10072 28448 10124
rect 28500 10112 28506 10124
rect 28767 10115 28825 10121
rect 28767 10112 28779 10115
rect 28500 10084 28779 10112
rect 28500 10072 28506 10084
rect 28767 10081 28779 10084
rect 28813 10081 28825 10115
rect 28767 10075 28825 10081
rect 29089 10115 29147 10121
rect 29089 10081 29101 10115
rect 29135 10112 29147 10115
rect 29454 10112 29460 10124
rect 29135 10084 29460 10112
rect 29135 10081 29147 10084
rect 29089 10075 29147 10081
rect 29454 10072 29460 10084
rect 29512 10072 29518 10124
rect 30742 10072 30748 10124
rect 30800 10072 30806 10124
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10044 28687 10047
rect 29270 10044 29276 10056
rect 28675 10016 29276 10044
rect 28675 10013 28687 10016
rect 28629 10007 28687 10013
rect 29270 10004 29276 10016
rect 29328 10004 29334 10056
rect 27080 9948 27660 9976
rect 27801 9979 27859 9985
rect 27801 9945 27813 9979
rect 27847 9976 27859 9979
rect 28074 9976 28080 9988
rect 27847 9948 28080 9976
rect 27847 9945 27859 9948
rect 27801 9939 27859 9945
rect 28074 9936 28080 9948
rect 28132 9936 28138 9988
rect 26050 9908 26056 9920
rect 25240 9880 26056 9908
rect 26050 9868 26056 9880
rect 26108 9868 26114 9920
rect 27890 9868 27896 9920
rect 27948 9868 27954 9920
rect 29178 9868 29184 9920
rect 29236 9908 29242 9920
rect 29365 9911 29423 9917
rect 29365 9908 29377 9911
rect 29236 9880 29377 9908
rect 29236 9868 29242 9880
rect 29365 9877 29377 9880
rect 29411 9877 29423 9911
rect 29365 9871 29423 9877
rect 552 9818 31648 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 11436 9818
rect 11488 9766 11500 9818
rect 11552 9766 11564 9818
rect 11616 9766 11628 9818
rect 11680 9766 11692 9818
rect 11744 9766 19210 9818
rect 19262 9766 19274 9818
rect 19326 9766 19338 9818
rect 19390 9766 19402 9818
rect 19454 9766 19466 9818
rect 19518 9766 26984 9818
rect 27036 9766 27048 9818
rect 27100 9766 27112 9818
rect 27164 9766 27176 9818
rect 27228 9766 27240 9818
rect 27292 9766 31648 9818
rect 552 9744 31648 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 3053 9707 3111 9713
rect 3053 9704 3065 9707
rect 2832 9676 3065 9704
rect 2832 9664 2838 9676
rect 3053 9673 3065 9676
rect 3099 9673 3111 9707
rect 3053 9667 3111 9673
rect 4249 9707 4307 9713
rect 4249 9673 4261 9707
rect 4295 9704 4307 9707
rect 4525 9707 4583 9713
rect 4295 9676 4384 9704
rect 4295 9673 4307 9676
rect 4249 9667 4307 9673
rect 3068 9636 3096 9667
rect 3418 9636 3424 9648
rect 3068 9608 3424 9636
rect 3418 9596 3424 9608
rect 3476 9636 3482 9648
rect 3476 9608 4016 9636
rect 3476 9596 3482 9608
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 2924 9540 3801 9568
rect 2924 9528 2930 9540
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 1305 9503 1363 9509
rect 1305 9469 1317 9503
rect 1351 9500 1363 9503
rect 1394 9500 1400 9512
rect 1351 9472 1400 9500
rect 1351 9469 1363 9472
rect 1305 9463 1363 9469
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1946 9509 1952 9512
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1535 9472 1685 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1940 9500 1952 9509
rect 1907 9472 1952 9500
rect 1673 9463 1731 9469
rect 1940 9463 1952 9472
rect 1946 9460 1952 9463
rect 2004 9460 2010 9512
rect 3988 9509 4016 9608
rect 4356 9568 4384 9676
rect 4525 9673 4537 9707
rect 4571 9704 4583 9707
rect 5350 9704 5356 9716
rect 4571 9676 5356 9704
rect 4571 9673 4583 9676
rect 4525 9667 4583 9673
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5445 9707 5503 9713
rect 5445 9673 5457 9707
rect 5491 9704 5503 9707
rect 5718 9704 5724 9716
rect 5491 9676 5724 9704
rect 5491 9673 5503 9676
rect 5445 9667 5503 9673
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 5960 9676 6285 9704
rect 5960 9664 5966 9676
rect 6273 9673 6285 9676
rect 6319 9673 6331 9707
rect 6273 9667 6331 9673
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 8754 9704 8760 9716
rect 7156 9676 8760 9704
rect 7156 9664 7162 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 10410 9704 10416 9716
rect 9692 9676 10416 9704
rect 4433 9639 4491 9645
rect 4433 9605 4445 9639
rect 4479 9636 4491 9639
rect 4706 9636 4712 9648
rect 4479 9608 4712 9636
rect 4479 9605 4491 9608
rect 4433 9599 4491 9605
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 4982 9636 4988 9648
rect 4816 9608 4988 9636
rect 4816 9568 4844 9608
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 5169 9639 5227 9645
rect 5169 9605 5181 9639
rect 5215 9636 5227 9639
rect 5994 9636 6000 9648
rect 5215 9608 6000 9636
rect 5215 9605 5227 9608
rect 5169 9599 5227 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 5626 9568 5632 9580
rect 4356 9540 4844 9568
rect 5000 9540 5632 9568
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9500 4307 9503
rect 4614 9500 4620 9512
rect 4295 9472 4620 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 3237 9435 3295 9441
rect 3237 9432 3249 9435
rect 2648 9404 3249 9432
rect 2648 9392 2654 9404
rect 3237 9401 3249 9404
rect 3283 9401 3295 9435
rect 4724 9432 4752 9463
rect 4890 9460 4896 9512
rect 4948 9460 4954 9512
rect 5000 9509 5028 9540
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6748 9568 6776 9599
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 6880 9608 6960 9636
rect 6880 9596 6886 9608
rect 5776 9540 6776 9568
rect 6932 9568 6960 9608
rect 6932 9540 8524 9568
rect 5776 9528 5782 9540
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 5583 9472 5764 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 5736 9444 5764 9472
rect 5810 9460 5816 9512
rect 5868 9460 5874 9512
rect 5994 9460 6000 9512
rect 6052 9460 6058 9512
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 6362 9500 6368 9512
rect 6227 9472 6368 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 6454 9460 6460 9512
rect 6512 9460 6518 9512
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6932 9500 6960 9540
rect 6871 9472 6960 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 4724 9404 5120 9432
rect 3237 9395 3295 9401
rect 1210 9324 1216 9376
rect 1268 9324 1274 9376
rect 5092 9364 5120 9404
rect 5718 9392 5724 9444
rect 5776 9392 5782 9444
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9432 5963 9435
rect 6564 9432 6592 9463
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 7650 9500 7656 9512
rect 7607 9472 7656 9500
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8294 9500 8300 9512
rect 7975 9472 8300 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 5951 9404 6592 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 5092 9336 5641 9364
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 6564 9364 6592 9404
rect 7282 9392 7288 9444
rect 7340 9392 7346 9444
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7760 9432 7788 9463
rect 7515 9404 7788 9432
rect 7852 9432 7880 9463
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 8496 9500 8524 9540
rect 9692 9500 9720 9676
rect 10410 9664 10416 9676
rect 10468 9704 10474 9716
rect 10468 9676 11100 9704
rect 10468 9664 10474 9676
rect 11072 9636 11100 9676
rect 13446 9664 13452 9716
rect 13504 9704 13510 9716
rect 13633 9707 13691 9713
rect 13633 9704 13645 9707
rect 13504 9676 13645 9704
rect 13504 9664 13510 9676
rect 13633 9673 13645 9676
rect 13679 9673 13691 9707
rect 13633 9667 13691 9673
rect 14645 9707 14703 9713
rect 14645 9673 14657 9707
rect 14691 9704 14703 9707
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14691 9676 14933 9704
rect 14691 9673 14703 9676
rect 14645 9667 14703 9673
rect 14921 9673 14933 9676
rect 14967 9704 14979 9707
rect 14967 9676 17632 9704
rect 14967 9673 14979 9676
rect 14921 9667 14979 9673
rect 17604 9648 17632 9676
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 20073 9707 20131 9713
rect 20073 9704 20085 9707
rect 20036 9676 20085 9704
rect 20036 9664 20042 9676
rect 20073 9673 20085 9676
rect 20119 9673 20131 9707
rect 20073 9667 20131 9673
rect 20530 9664 20536 9716
rect 20588 9704 20594 9716
rect 25774 9704 25780 9716
rect 20588 9676 25780 9704
rect 20588 9664 20594 9676
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 26234 9664 26240 9716
rect 26292 9704 26298 9716
rect 26421 9707 26479 9713
rect 26421 9704 26433 9707
rect 26292 9676 26433 9704
rect 26292 9664 26298 9676
rect 26421 9673 26433 9676
rect 26467 9704 26479 9707
rect 26786 9704 26792 9716
rect 26467 9676 26792 9704
rect 26467 9673 26479 9676
rect 26421 9667 26479 9673
rect 26786 9664 26792 9676
rect 26844 9664 26850 9716
rect 26878 9664 26884 9716
rect 26936 9704 26942 9716
rect 28810 9704 28816 9716
rect 26936 9676 28816 9704
rect 26936 9664 26942 9676
rect 28810 9664 28816 9676
rect 28868 9664 28874 9716
rect 28994 9664 29000 9716
rect 29052 9664 29058 9716
rect 29914 9664 29920 9716
rect 29972 9704 29978 9716
rect 30009 9707 30067 9713
rect 30009 9704 30021 9707
rect 29972 9676 30021 9704
rect 29972 9664 29978 9676
rect 30009 9673 30021 9676
rect 30055 9673 30067 9707
rect 30009 9667 30067 9673
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 11072 9608 11529 9636
rect 11517 9605 11529 9608
rect 11563 9605 11575 9639
rect 11517 9599 11575 9605
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12299 9608 12449 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 14737 9639 14795 9645
rect 14737 9636 14749 9639
rect 12437 9599 12495 9605
rect 13924 9608 14749 9636
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9999 9540 10149 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 8496 9472 9720 9500
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9500 10103 9503
rect 10686 9500 10692 9512
rect 10091 9472 10692 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 10686 9460 10692 9472
rect 10744 9500 10750 9512
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 10744 9472 11805 9500
rect 10744 9460 10750 9472
rect 11793 9469 11805 9472
rect 11839 9469 11851 9503
rect 11793 9463 11851 9469
rect 12066 9460 12072 9512
rect 12124 9460 12130 9512
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9500 12403 9503
rect 12526 9500 12532 9512
rect 12391 9472 12532 9500
rect 12391 9469 12403 9472
rect 12345 9463 12403 9469
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 8656 9435 8714 9441
rect 7852 9404 8340 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 7300 9364 7328 9392
rect 6564 9336 7328 9364
rect 5629 9327 5687 9333
rect 8202 9324 8208 9376
rect 8260 9324 8266 9376
rect 8312 9364 8340 9404
rect 8656 9401 8668 9435
rect 8702 9432 8714 9435
rect 8846 9432 8852 9444
rect 8702 9404 8852 9432
rect 8702 9401 8714 9404
rect 8656 9395 8714 9401
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10382 9435 10440 9441
rect 10382 9432 10394 9435
rect 10192 9404 10394 9432
rect 10192 9392 10198 9404
rect 10382 9401 10394 9404
rect 10428 9401 10440 9435
rect 10382 9395 10440 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 12636 9432 12664 9463
rect 12710 9460 12716 9512
rect 12768 9460 12774 9512
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 13924 9500 13952 9608
rect 14737 9605 14749 9608
rect 14783 9605 14795 9639
rect 14737 9599 14795 9605
rect 16485 9639 16543 9645
rect 16485 9605 16497 9639
rect 16531 9636 16543 9639
rect 17310 9636 17316 9648
rect 16531 9608 17316 9636
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 17586 9596 17592 9648
rect 17644 9636 17650 9648
rect 17644 9608 21119 9636
rect 17644 9596 17650 9608
rect 14550 9568 14556 9580
rect 14016 9540 14556 9568
rect 14016 9509 14044 9540
rect 14550 9528 14556 9540
rect 14608 9568 14614 9580
rect 14608 9540 15792 9568
rect 14608 9528 14614 9540
rect 13863 9472 13952 9500
rect 14001 9503 14059 9509
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 14001 9469 14013 9503
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14108 9432 14136 9463
rect 14274 9460 14280 9512
rect 14332 9460 14338 9512
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 14507 9472 14596 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14568 9444 14596 9472
rect 11112 9404 14136 9432
rect 11112 9392 11118 9404
rect 14550 9392 14556 9444
rect 14608 9392 14614 9444
rect 15105 9435 15163 9441
rect 15105 9401 15117 9435
rect 15151 9432 15163 9435
rect 15194 9432 15200 9444
rect 15151 9404 15200 9432
rect 15151 9401 15163 9404
rect 15105 9395 15163 9401
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 15764 9432 15792 9540
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16301 9571 16359 9577
rect 16301 9568 16313 9571
rect 15988 9540 16313 9568
rect 15988 9528 15994 9540
rect 16301 9537 16313 9540
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 19058 9568 19064 9580
rect 18196 9540 19064 9568
rect 18196 9528 18202 9540
rect 19058 9528 19064 9540
rect 19116 9568 19122 9580
rect 19116 9540 19472 9568
rect 19116 9528 19122 9540
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15896 9472 16037 9500
rect 15896 9460 15902 9472
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 16114 9460 16120 9512
rect 16172 9460 16178 9512
rect 16390 9460 16396 9512
rect 16448 9460 16454 9512
rect 18322 9460 18328 9512
rect 18380 9500 18386 9512
rect 19444 9509 19472 9540
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 18380 9472 19257 9500
rect 18380 9460 18386 9472
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9469 19487 9503
rect 20180 9500 20208 9608
rect 20806 9568 20812 9580
rect 20456 9540 20812 9568
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 20180 9472 20269 9500
rect 19429 9463 19487 9469
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 20346 9460 20352 9512
rect 20404 9460 20410 9512
rect 20456 9509 20484 9540
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 20441 9503 20499 9509
rect 20441 9469 20453 9503
rect 20487 9469 20499 9503
rect 20441 9463 20499 9469
rect 20714 9460 20720 9512
rect 20772 9460 20778 9512
rect 19334 9432 19340 9444
rect 15764 9404 19340 9432
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 20530 9392 20536 9444
rect 20588 9441 20594 9444
rect 20588 9435 20617 9441
rect 20605 9401 20617 9435
rect 21091 9432 21119 9608
rect 21174 9528 21180 9580
rect 21232 9568 21238 9580
rect 22186 9568 22192 9580
rect 21232 9540 22192 9568
rect 21232 9528 21238 9540
rect 22020 9509 22048 9540
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 27801 9571 27859 9577
rect 27801 9537 27813 9571
rect 27847 9568 27859 9571
rect 28445 9571 28503 9577
rect 28445 9568 28457 9571
rect 27847 9540 28457 9568
rect 27847 9537 27859 9540
rect 27801 9531 27859 9537
rect 28445 9537 28457 9540
rect 28491 9537 28503 9571
rect 28445 9531 28503 9537
rect 22554 9509 22560 9512
rect 22005 9503 22063 9509
rect 22005 9469 22017 9503
rect 22051 9469 22063 9503
rect 22005 9463 22063 9469
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9500 22155 9503
rect 22281 9503 22339 9509
rect 22281 9500 22293 9503
rect 22143 9472 22293 9500
rect 22143 9469 22155 9472
rect 22097 9463 22155 9469
rect 22281 9469 22293 9472
rect 22327 9469 22339 9503
rect 22548 9500 22560 9509
rect 22515 9472 22560 9500
rect 22281 9463 22339 9469
rect 22548 9463 22560 9472
rect 22554 9460 22560 9463
rect 22612 9460 22618 9512
rect 23845 9503 23903 9509
rect 23845 9469 23857 9503
rect 23891 9500 23903 9503
rect 24486 9500 24492 9512
rect 23891 9472 24492 9500
rect 23891 9469 23903 9472
rect 23845 9463 23903 9469
rect 24486 9460 24492 9472
rect 24544 9460 24550 9512
rect 25869 9503 25927 9509
rect 25869 9500 25881 9503
rect 25240 9472 25881 9500
rect 23566 9432 23572 9444
rect 21091 9404 23572 9432
rect 20588 9395 20617 9401
rect 20588 9392 20594 9395
rect 23566 9392 23572 9404
rect 23624 9392 23630 9444
rect 24112 9435 24170 9441
rect 24112 9401 24124 9435
rect 24158 9432 24170 9435
rect 24302 9432 24308 9444
rect 24158 9404 24308 9432
rect 24158 9401 24170 9404
rect 24112 9395 24170 9401
rect 24302 9392 24308 9404
rect 24360 9392 24366 9444
rect 25240 9376 25268 9472
rect 25869 9469 25881 9472
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 27545 9503 27603 9509
rect 27545 9469 27557 9503
rect 27591 9500 27603 9503
rect 27890 9500 27896 9512
rect 27591 9472 27896 9500
rect 27591 9469 27603 9472
rect 27545 9463 27603 9469
rect 27890 9460 27896 9472
rect 27948 9460 27954 9512
rect 28077 9503 28135 9509
rect 28077 9469 28089 9503
rect 28123 9500 28135 9503
rect 28166 9500 28172 9512
rect 28123 9472 28172 9500
rect 28123 9469 28135 9472
rect 28077 9463 28135 9469
rect 28166 9460 28172 9472
rect 28224 9460 28230 9512
rect 28261 9503 28319 9509
rect 28261 9469 28273 9503
rect 28307 9469 28319 9503
rect 28261 9463 28319 9469
rect 26050 9392 26056 9444
rect 26108 9432 26114 9444
rect 26108 9404 28120 9432
rect 26108 9392 26114 9404
rect 9122 9364 9128 9376
rect 8312 9336 9128 9364
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11664 9336 11713 9364
rect 11664 9324 11670 9336
rect 11701 9333 11713 9336
rect 11747 9333 11759 9367
rect 11701 9327 11759 9333
rect 11882 9324 11888 9376
rect 11940 9324 11946 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 14895 9367 14953 9373
rect 14895 9364 14907 9367
rect 14792 9336 14907 9364
rect 14792 9324 14798 9336
rect 14895 9333 14907 9336
rect 14941 9333 14953 9367
rect 14895 9327 14953 9333
rect 19521 9367 19579 9373
rect 19521 9333 19533 9367
rect 19567 9364 19579 9367
rect 19610 9364 19616 9376
rect 19567 9336 19616 9364
rect 19567 9333 19579 9336
rect 19521 9327 19579 9333
rect 19610 9324 19616 9336
rect 19668 9364 19674 9376
rect 21634 9364 21640 9376
rect 19668 9336 21640 9364
rect 19668 9324 19674 9336
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 23661 9367 23719 9373
rect 23661 9333 23673 9367
rect 23707 9364 23719 9367
rect 23750 9364 23756 9376
rect 23707 9336 23756 9364
rect 23707 9333 23719 9336
rect 23661 9327 23719 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 25222 9324 25228 9376
rect 25280 9324 25286 9376
rect 25314 9324 25320 9376
rect 25372 9324 25378 9376
rect 27893 9367 27951 9373
rect 27893 9333 27905 9367
rect 27939 9364 27951 9367
rect 27982 9364 27988 9376
rect 27939 9336 27988 9364
rect 27939 9333 27951 9336
rect 27893 9327 27951 9333
rect 27982 9324 27988 9336
rect 28040 9324 28046 9376
rect 28092 9364 28120 9404
rect 28276 9364 28304 9463
rect 28534 9460 28540 9512
rect 28592 9500 28598 9512
rect 28813 9503 28871 9509
rect 28813 9500 28825 9503
rect 28592 9472 28825 9500
rect 28592 9460 28598 9472
rect 28813 9469 28825 9472
rect 28859 9500 28871 9503
rect 29012 9500 29040 9664
rect 29178 9528 29184 9580
rect 29236 9568 29242 9580
rect 29236 9540 29960 9568
rect 29236 9528 29242 9540
rect 29932 9509 29960 9540
rect 29549 9503 29607 9509
rect 29549 9500 29561 9503
rect 28859 9472 29561 9500
rect 28859 9469 28871 9472
rect 28813 9463 28871 9469
rect 29549 9469 29561 9472
rect 29595 9469 29607 9503
rect 29549 9463 29607 9469
rect 29917 9503 29975 9509
rect 29917 9469 29929 9503
rect 29963 9469 29975 9503
rect 29917 9463 29975 9469
rect 28092 9336 28304 9364
rect 28718 9324 28724 9376
rect 28776 9324 28782 9376
rect 29270 9324 29276 9376
rect 29328 9364 29334 9376
rect 29457 9367 29515 9373
rect 29457 9364 29469 9367
rect 29328 9336 29469 9364
rect 29328 9324 29334 9336
rect 29457 9333 29469 9336
rect 29503 9333 29515 9367
rect 29457 9327 29515 9333
rect 552 9274 31648 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 12096 9274
rect 12148 9222 12160 9274
rect 12212 9222 12224 9274
rect 12276 9222 12288 9274
rect 12340 9222 12352 9274
rect 12404 9222 19870 9274
rect 19922 9222 19934 9274
rect 19986 9222 19998 9274
rect 20050 9222 20062 9274
rect 20114 9222 20126 9274
rect 20178 9222 27644 9274
rect 27696 9222 27708 9274
rect 27760 9222 27772 9274
rect 27824 9222 27836 9274
rect 27888 9222 27900 9274
rect 27952 9222 31648 9274
rect 552 9200 31648 9222
rect 5810 9160 5816 9172
rect 3620 9132 5816 9160
rect 1210 8984 1216 9036
rect 1268 9024 1274 9036
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1268 8996 1961 9024
rect 1268 8984 1274 8996
rect 1949 8993 1961 8996
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2216 9027 2274 9033
rect 2216 8993 2228 9027
rect 2262 9024 2274 9027
rect 2498 9024 2504 9036
rect 2262 8996 2504 9024
rect 2262 8993 2274 8996
rect 2216 8987 2274 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 3620 9033 3648 9132
rect 5810 9120 5816 9132
rect 5868 9160 5874 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 5868 9132 6193 9160
rect 5868 9120 5874 9132
rect 6181 9129 6193 9132
rect 6227 9160 6239 9163
rect 6454 9160 6460 9172
rect 6227 9132 6460 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 7340 9132 9045 9160
rect 7340 9120 7346 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9398 9120 9404 9172
rect 9456 9160 9462 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 9456 9132 9505 9160
rect 9456 9120 9462 9132
rect 9493 9129 9505 9132
rect 9539 9129 9551 9163
rect 9493 9123 9551 9129
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 11756 9132 12434 9160
rect 11756 9120 11762 9132
rect 8294 9092 8300 9104
rect 6012 9064 8300 9092
rect 6012 9036 6040 9064
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 8993 3663 9027
rect 3605 8987 3663 8993
rect 5994 8984 6000 9036
rect 6052 8984 6058 9036
rect 7392 9033 7420 9064
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 8754 9052 8760 9104
rect 8812 9092 8818 9104
rect 9125 9095 9183 9101
rect 9125 9092 9137 9095
rect 8812 9064 9137 9092
rect 8812 9052 8818 9064
rect 9125 9061 9137 9064
rect 9171 9061 9183 9095
rect 10318 9092 10324 9104
rect 9125 9055 9183 9061
rect 9232 9064 10324 9092
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 8993 6147 9027
rect 6089 8987 6147 8993
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7920 9027 7978 9033
rect 7920 8993 7932 9027
rect 7966 9024 7978 9027
rect 8202 9024 8208 9036
rect 7966 8996 8208 9024
rect 7966 8993 7978 8996
rect 7920 8987 7978 8993
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3510 8956 3516 8968
rect 3292 8928 3516 8956
rect 3292 8916 3298 8928
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4338 8956 4344 8968
rect 4295 8928 4344 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4982 8916 4988 8968
rect 5040 8916 5046 8968
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8956 5595 8959
rect 6104 8956 6132 8987
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9232 9024 9260 9064
rect 10318 9052 10324 9064
rect 10376 9092 10382 9104
rect 11784 9095 11842 9101
rect 10376 9064 11744 9092
rect 10376 9052 10382 9064
rect 8536 8996 9260 9024
rect 9309 9027 9367 9033
rect 8536 8984 8542 8996
rect 9309 8993 9321 9027
rect 9355 9024 9367 9027
rect 9766 9024 9772 9036
rect 9355 8996 9772 9024
rect 9355 8993 9367 8996
rect 9309 8987 9367 8993
rect 5583 8928 6132 8956
rect 7469 8959 7527 8965
rect 5583 8925 5595 8928
rect 5537 8919 5595 8925
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 7515 8928 7665 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 7653 8925 7665 8928
rect 7699 8925 7711 8959
rect 9324 8956 9352 8987
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 11517 9027 11575 9033
rect 11517 8993 11529 9027
rect 11563 9024 11575 9027
rect 11606 9024 11612 9036
rect 11563 8996 11612 9024
rect 11563 8993 11575 8996
rect 11517 8987 11575 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11716 9024 11744 9064
rect 11784 9061 11796 9095
rect 11830 9092 11842 9095
rect 11882 9092 11888 9104
rect 11830 9064 11888 9092
rect 11830 9061 11842 9064
rect 11784 9055 11842 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 12406 9092 12434 9132
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12584 9132 13001 9160
rect 12584 9120 12590 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 13157 9163 13215 9169
rect 13157 9129 13169 9163
rect 13203 9160 13215 9163
rect 14734 9160 14740 9172
rect 13203 9132 14740 9160
rect 13203 9129 13215 9132
rect 13157 9123 13215 9129
rect 13157 9092 13185 9123
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16172 9132 16957 9160
rect 16172 9120 16178 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 22281 9163 22339 9169
rect 22281 9129 22293 9163
rect 22327 9160 22339 9163
rect 22370 9160 22376 9172
rect 22327 9132 22376 9160
rect 22327 9129 22339 9132
rect 22281 9123 22339 9129
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 22554 9120 22560 9172
rect 22612 9160 22618 9172
rect 22738 9160 22744 9172
rect 22612 9132 22744 9160
rect 22612 9120 22618 9132
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 27430 9160 27436 9172
rect 22888 9132 27436 9160
rect 22888 9120 22894 9132
rect 12406 9064 13185 9092
rect 13357 9095 13415 9101
rect 13357 9061 13369 9095
rect 13403 9092 13415 9095
rect 14550 9092 14556 9104
rect 13403 9064 14556 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 18782 9052 18788 9104
rect 18840 9092 18846 9104
rect 22097 9095 22155 9101
rect 18840 9064 21036 9092
rect 18840 9052 18846 9064
rect 12710 9024 12716 9036
rect 11716 8996 12716 9024
rect 12710 8984 12716 8996
rect 12768 9024 12774 9036
rect 14458 9024 14464 9036
rect 12768 8996 14464 9024
rect 12768 8984 12774 8996
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 15013 9027 15071 9033
rect 15013 8993 15025 9027
rect 15059 9024 15071 9027
rect 15286 9024 15292 9036
rect 15059 8996 15292 9024
rect 15059 8993 15071 8996
rect 15013 8987 15071 8993
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 15565 9027 15623 9033
rect 15565 8993 15577 9027
rect 15611 9024 15623 9027
rect 15654 9024 15660 9036
rect 15611 8996 15660 9024
rect 15611 8993 15623 8996
rect 15565 8987 15623 8993
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 8993 17187 9027
rect 17129 8987 17187 8993
rect 17313 9027 17371 9033
rect 17313 8993 17325 9027
rect 17359 9024 17371 9027
rect 17402 9024 17408 9036
rect 17359 8996 17408 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 7653 8919 7711 8925
rect 9232 8928 9352 8956
rect 15197 8959 15255 8965
rect 3973 8891 4031 8897
rect 3973 8857 3985 8891
rect 4019 8888 4031 8891
rect 4062 8888 4068 8900
rect 4019 8860 4068 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 3329 8823 3387 8829
rect 3329 8789 3341 8823
rect 3375 8820 3387 8823
rect 3510 8820 3516 8832
rect 3375 8792 3516 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 3510 8780 3516 8792
rect 3568 8820 3574 8832
rect 4246 8820 4252 8832
rect 3568 8792 4252 8820
rect 3568 8780 3574 8792
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 5868 8792 5917 8820
rect 5868 8780 5874 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 5905 8783 5963 8789
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 9232 8820 9260 8928
rect 15197 8925 15209 8959
rect 15243 8925 15255 8959
rect 17144 8956 17172 8987
rect 17402 8984 17408 8996
rect 17460 9024 17466 9036
rect 17460 8996 18460 9024
rect 17460 8984 17466 8996
rect 18432 8968 18460 8996
rect 18506 8984 18512 9036
rect 18564 8984 18570 9036
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 9024 19211 9027
rect 20073 9027 20131 9033
rect 19199 8996 20024 9024
rect 19199 8993 19211 8996
rect 19153 8987 19211 8993
rect 18138 8956 18144 8968
rect 17144 8928 18144 8956
rect 15197 8919 15255 8925
rect 12897 8891 12955 8897
rect 12897 8857 12909 8891
rect 12943 8888 12955 8891
rect 12943 8860 13216 8888
rect 12943 8857 12955 8860
rect 12897 8851 12955 8857
rect 13188 8829 13216 8860
rect 14274 8848 14280 8900
rect 14332 8888 14338 8900
rect 15212 8888 15240 8919
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 15381 8891 15439 8897
rect 15381 8888 15393 8891
rect 14332 8860 15393 8888
rect 14332 8848 14338 8860
rect 15381 8857 15393 8860
rect 15427 8857 15439 8891
rect 15381 8851 15439 8857
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 18340 8888 18368 8919
rect 18414 8916 18420 8968
rect 18472 8956 18478 8968
rect 19061 8959 19119 8965
rect 19061 8956 19073 8959
rect 18472 8928 19073 8956
rect 18472 8916 18478 8928
rect 19061 8925 19073 8928
rect 19107 8925 19119 8959
rect 19889 8959 19947 8965
rect 19889 8956 19901 8959
rect 19061 8919 19119 8925
rect 19168 8928 19901 8956
rect 18966 8888 18972 8900
rect 18012 8860 18972 8888
rect 18012 8848 18018 8860
rect 18966 8848 18972 8860
rect 19024 8888 19030 8900
rect 19168 8888 19196 8928
rect 19889 8925 19901 8928
rect 19935 8925 19947 8959
rect 19996 8956 20024 8996
rect 20073 8993 20085 9027
rect 20119 9024 20131 9027
rect 20346 9024 20352 9036
rect 20119 8996 20352 9024
rect 20119 8993 20131 8996
rect 20073 8987 20131 8993
rect 20346 8984 20352 8996
rect 20404 8984 20410 9036
rect 21008 9033 21036 9064
rect 22097 9061 22109 9095
rect 22143 9092 22155 9095
rect 22186 9092 22192 9104
rect 22143 9064 22192 9092
rect 22143 9061 22155 9064
rect 22097 9055 22155 9061
rect 22186 9052 22192 9064
rect 22244 9052 22250 9104
rect 22572 9092 22600 9120
rect 23834 9101 23862 9132
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 23819 9095 23877 9101
rect 22572 9064 22692 9092
rect 20993 9027 21051 9033
rect 20993 8993 21005 9027
rect 21039 9024 21051 9027
rect 21174 9024 21180 9036
rect 21039 8996 21180 9024
rect 21039 8993 21051 8996
rect 20993 8987 21051 8993
rect 21174 8984 21180 8996
rect 21232 8984 21238 9036
rect 21266 8984 21272 9036
rect 21324 8984 21330 9036
rect 22370 8984 22376 9036
rect 22428 9024 22434 9036
rect 22664 9033 22692 9064
rect 23819 9061 23831 9095
rect 23865 9061 23877 9095
rect 23819 9055 23877 9061
rect 23937 9095 23995 9101
rect 23937 9061 23949 9095
rect 23983 9092 23995 9095
rect 25314 9092 25320 9104
rect 23983 9064 25320 9092
rect 23983 9061 23995 9064
rect 23937 9055 23995 9061
rect 25314 9052 25320 9064
rect 25372 9052 25378 9104
rect 26510 9052 26516 9104
rect 26568 9092 26574 9104
rect 27522 9092 27528 9104
rect 26568 9064 27528 9092
rect 26568 9052 26574 9064
rect 27522 9052 27528 9064
rect 27580 9052 27586 9104
rect 27648 9095 27706 9101
rect 27648 9061 27660 9095
rect 27694 9092 27706 9095
rect 27982 9092 27988 9104
rect 27694 9064 27988 9092
rect 27694 9061 27706 9064
rect 27648 9055 27706 9061
rect 27982 9052 27988 9064
rect 28040 9052 28046 9104
rect 29181 9095 29239 9101
rect 29181 9061 29193 9095
rect 29227 9092 29239 9095
rect 29518 9095 29576 9101
rect 29518 9092 29530 9095
rect 29227 9064 29530 9092
rect 29227 9061 29239 9064
rect 29181 9055 29239 9061
rect 29518 9061 29530 9064
rect 29564 9061 29576 9095
rect 29518 9055 29576 9061
rect 22830 9033 22836 9036
rect 22465 9027 22523 9033
rect 22465 9024 22477 9027
rect 22428 8996 22477 9024
rect 22428 8984 22434 8996
rect 22465 8993 22477 8996
rect 22511 8993 22523 9027
rect 22465 8987 22523 8993
rect 22557 9027 22615 9033
rect 22557 8993 22569 9027
rect 22603 8993 22615 9027
rect 22557 8987 22615 8993
rect 22649 9027 22707 9033
rect 22649 8993 22661 9027
rect 22695 8993 22707 9027
rect 22649 8987 22707 8993
rect 22787 9027 22836 9033
rect 22787 8993 22799 9027
rect 22833 8993 22836 9027
rect 22787 8987 22836 8993
rect 22278 8956 22284 8968
rect 19996 8928 22284 8956
rect 19889 8919 19947 8925
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 22572 8956 22600 8987
rect 22830 8984 22836 8987
rect 22888 8984 22894 9036
rect 23566 8984 23572 9036
rect 23624 9024 23630 9036
rect 24026 9024 24032 9036
rect 23624 8996 24032 9024
rect 23624 8984 23630 8996
rect 24026 8984 24032 8996
rect 24084 8984 24090 9036
rect 24118 8984 24124 9036
rect 24176 9024 24182 9036
rect 24581 9027 24639 9033
rect 24176 8996 24532 9024
rect 24176 8984 24182 8996
rect 22572 8928 22692 8956
rect 19702 8888 19708 8900
rect 19024 8860 19196 8888
rect 19306 8860 19708 8888
rect 19024 8848 19030 8860
rect 6420 8792 9260 8820
rect 13173 8823 13231 8829
rect 6420 8780 6426 8792
rect 13173 8789 13185 8823
rect 13219 8820 13231 8823
rect 13538 8820 13544 8832
rect 13219 8792 13544 8820
rect 13219 8789 13231 8792
rect 13173 8783 13231 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 14826 8780 14832 8832
rect 14884 8780 14890 8832
rect 18690 8780 18696 8832
rect 18748 8780 18754 8832
rect 18785 8823 18843 8829
rect 18785 8789 18797 8823
rect 18831 8820 18843 8823
rect 18874 8820 18880 8832
rect 18831 8792 18880 8820
rect 18831 8789 18843 8792
rect 18785 8783 18843 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19153 8823 19211 8829
rect 19153 8789 19165 8823
rect 19199 8820 19211 8823
rect 19306 8820 19334 8860
rect 19702 8848 19708 8860
rect 19760 8888 19766 8900
rect 21818 8888 21824 8900
rect 19760 8860 21824 8888
rect 19760 8848 19766 8860
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 22664 8888 22692 8928
rect 22922 8916 22928 8968
rect 22980 8916 22986 8968
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8956 23719 8959
rect 24210 8956 24216 8968
rect 23707 8928 24216 8956
rect 23707 8925 23719 8928
rect 23661 8919 23719 8925
rect 24210 8916 24216 8928
rect 24268 8916 24274 8968
rect 24302 8916 24308 8968
rect 24360 8916 24366 8968
rect 24504 8956 24532 8996
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 24854 9024 24860 9036
rect 24627 8996 24860 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 27893 9027 27951 9033
rect 27893 8993 27905 9027
rect 27939 9024 27951 9027
rect 28718 9024 28724 9036
rect 27939 8996 28724 9024
rect 27939 8993 27951 8996
rect 27893 8987 27951 8993
rect 28718 8984 28724 8996
rect 28776 8984 28782 9036
rect 28994 8984 29000 9036
rect 29052 8984 29058 9036
rect 29270 8984 29276 9036
rect 29328 8984 29334 9036
rect 24504 8928 26648 8956
rect 23750 8888 23756 8900
rect 22664 8860 23756 8888
rect 23750 8848 23756 8860
rect 23808 8888 23814 8900
rect 24578 8888 24584 8900
rect 23808 8860 24584 8888
rect 23808 8848 23814 8860
rect 24578 8848 24584 8860
rect 24636 8848 24642 8900
rect 26510 8848 26516 8900
rect 26568 8848 26574 8900
rect 19199 8792 19334 8820
rect 20257 8823 20315 8829
rect 19199 8789 19211 8792
rect 19153 8783 19211 8789
rect 20257 8789 20269 8823
rect 20303 8820 20315 8823
rect 20898 8820 20904 8832
rect 20303 8792 20904 8820
rect 20303 8789 20315 8792
rect 20257 8783 20315 8789
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 24486 8780 24492 8832
rect 24544 8780 24550 8832
rect 25774 8780 25780 8832
rect 25832 8820 25838 8832
rect 26326 8820 26332 8832
rect 25832 8792 26332 8820
rect 25832 8780 25838 8792
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 26620 8820 26648 8928
rect 28626 8916 28632 8968
rect 28684 8956 28690 8968
rect 28813 8959 28871 8965
rect 28813 8956 28825 8959
rect 28684 8928 28825 8956
rect 28684 8916 28690 8928
rect 28813 8925 28825 8928
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 29454 8820 29460 8832
rect 26620 8792 29460 8820
rect 29454 8780 29460 8792
rect 29512 8780 29518 8832
rect 30650 8780 30656 8832
rect 30708 8780 30714 8832
rect 552 8730 31648 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 11436 8730
rect 11488 8678 11500 8730
rect 11552 8678 11564 8730
rect 11616 8678 11628 8730
rect 11680 8678 11692 8730
rect 11744 8678 19210 8730
rect 19262 8678 19274 8730
rect 19326 8678 19338 8730
rect 19390 8678 19402 8730
rect 19454 8678 19466 8730
rect 19518 8678 26984 8730
rect 27036 8678 27048 8730
rect 27100 8678 27112 8730
rect 27164 8678 27176 8730
rect 27228 8678 27240 8730
rect 27292 8678 31648 8730
rect 552 8656 31648 8678
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 2593 8619 2651 8625
rect 2593 8616 2605 8619
rect 2556 8588 2605 8616
rect 2556 8576 2562 8588
rect 2593 8585 2605 8588
rect 2639 8585 2651 8619
rect 2593 8579 2651 8585
rect 3234 8576 3240 8628
rect 3292 8576 3298 8628
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 5994 8616 6000 8628
rect 3804 8588 6000 8616
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1452 8452 2912 8480
rect 1452 8440 1458 8452
rect 2590 8372 2596 8424
rect 2648 8372 2654 8424
rect 2884 8421 2912 8452
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8381 2835 8415
rect 2777 8375 2835 8381
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3804 8412 3832 8588
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 8444 8588 8585 8616
rect 8444 8576 8450 8588
rect 8573 8585 8585 8588
rect 8619 8585 8631 8619
rect 8573 8579 8631 8585
rect 13633 8619 13691 8625
rect 13633 8585 13645 8619
rect 13679 8616 13691 8619
rect 17402 8616 17408 8628
rect 13679 8588 17408 8616
rect 13679 8585 13691 8588
rect 13633 8579 13691 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 18966 8576 18972 8628
rect 19024 8616 19030 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19024 8588 20085 8616
rect 19024 8576 19030 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 21324 8588 21588 8616
rect 21324 8576 21330 8588
rect 4338 8508 4344 8560
rect 4396 8508 4402 8560
rect 18690 8508 18696 8560
rect 18748 8508 18754 8560
rect 21560 8548 21588 8588
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 22370 8616 22376 8628
rect 21692 8588 22376 8616
rect 21692 8576 21698 8588
rect 22370 8576 22376 8588
rect 22428 8616 22434 8628
rect 22738 8616 22744 8628
rect 22428 8588 22744 8616
rect 22428 8576 22434 8588
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 22922 8576 22928 8628
rect 22980 8616 22986 8628
rect 25593 8619 25651 8625
rect 25593 8616 25605 8619
rect 22980 8588 25605 8616
rect 22980 8576 22986 8588
rect 25593 8585 25605 8588
rect 25639 8585 25651 8619
rect 25593 8579 25651 8585
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 25958 8616 25964 8628
rect 25740 8588 25964 8616
rect 25740 8576 25746 8588
rect 25958 8576 25964 8588
rect 26016 8576 26022 8628
rect 28534 8616 28540 8628
rect 28092 8588 28540 8616
rect 21560 8520 26556 8548
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4154 8480 4160 8492
rect 4111 8452 4160 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 18708 8480 18736 8508
rect 16347 8452 16896 8480
rect 18708 8452 18828 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 2915 8384 3832 8412
rect 3973 8415 4031 8421
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3973 8381 3985 8415
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 2792 8344 2820 8375
rect 3234 8344 3240 8356
rect 2792 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 3418 8353 3424 8356
rect 3405 8347 3424 8353
rect 3405 8313 3417 8347
rect 3405 8307 3424 8313
rect 3418 8304 3424 8307
rect 3476 8304 3482 8356
rect 3510 8304 3516 8356
rect 3568 8344 3574 8356
rect 3605 8347 3663 8353
rect 3605 8344 3617 8347
rect 3568 8316 3617 8344
rect 3568 8304 3574 8316
rect 3605 8313 3617 8316
rect 3651 8313 3663 8347
rect 3988 8344 4016 8375
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 5546 8415 5604 8421
rect 5546 8412 5558 8415
rect 4856 8384 5558 8412
rect 4856 8372 4862 8384
rect 5546 8381 5558 8384
rect 5592 8381 5604 8415
rect 5546 8375 5604 8381
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 5776 8384 6469 8412
rect 5776 8372 5782 8384
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 8352 8384 8677 8412
rect 8352 8372 8358 8384
rect 8665 8381 8677 8384
rect 8711 8412 8723 8415
rect 9306 8412 9312 8424
rect 8711 8384 9312 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 13538 8372 13544 8424
rect 13596 8372 13602 8424
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 13780 8384 14473 8412
rect 13780 8372 13786 8384
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 14599 8384 14749 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 14737 8381 14749 8384
rect 14783 8381 14795 8415
rect 14737 8375 14795 8381
rect 14826 8372 14832 8424
rect 14884 8412 14890 8424
rect 14993 8415 15051 8421
rect 14993 8412 15005 8415
rect 14884 8384 15005 8412
rect 14884 8372 14890 8384
rect 14993 8381 15005 8384
rect 15039 8381 15051 8415
rect 14993 8375 15051 8381
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8412 16543 8415
rect 16574 8412 16580 8424
rect 16531 8384 16580 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 16758 8372 16764 8424
rect 16816 8372 16822 8424
rect 16868 8412 16896 8452
rect 17954 8412 17960 8424
rect 16868 8384 17960 8412
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 18417 8415 18475 8421
rect 18417 8381 18429 8415
rect 18463 8412 18475 8415
rect 18693 8415 18751 8421
rect 18693 8412 18705 8415
rect 18463 8384 18705 8412
rect 18463 8381 18475 8384
rect 18417 8375 18475 8381
rect 18693 8381 18705 8384
rect 18739 8381 18751 8415
rect 18800 8412 18828 8452
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 24302 8480 24308 8492
rect 22060 8452 24308 8480
rect 22060 8440 22066 8452
rect 20898 8421 20904 8424
rect 18949 8415 19007 8421
rect 18949 8412 18961 8415
rect 18800 8384 18961 8412
rect 18693 8375 18751 8381
rect 18949 8381 18961 8384
rect 18995 8381 19007 8415
rect 18949 8375 19007 8381
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8381 20407 8415
rect 20349 8375 20407 8381
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8412 20499 8415
rect 20625 8415 20683 8421
rect 20625 8412 20637 8415
rect 20487 8384 20637 8412
rect 20487 8381 20499 8384
rect 20441 8375 20499 8381
rect 20625 8381 20637 8384
rect 20671 8381 20683 8415
rect 20892 8412 20904 8421
rect 20859 8384 20904 8412
rect 20625 8375 20683 8381
rect 20892 8375 20904 8384
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 3988 8316 5917 8344
rect 3605 8307 3663 8313
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 5905 8307 5963 8313
rect 16669 8347 16727 8353
rect 16669 8313 16681 8347
rect 16715 8344 16727 8347
rect 17006 8347 17064 8353
rect 17006 8344 17018 8347
rect 16715 8316 17018 8344
rect 16715 8313 16727 8316
rect 16669 8307 16727 8313
rect 17006 8313 17018 8316
rect 17052 8313 17064 8347
rect 18340 8344 18368 8375
rect 18782 8344 18788 8356
rect 17006 8307 17064 8313
rect 17880 8316 18788 8344
rect 2958 8236 2964 8288
rect 3016 8236 3022 8288
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4706 8276 4712 8288
rect 4479 8248 4712 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4706 8236 4712 8248
rect 4764 8276 4770 8288
rect 5718 8276 5724 8288
rect 4764 8248 5724 8276
rect 4764 8236 4770 8248
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11330 8276 11336 8288
rect 11112 8248 11336 8276
rect 11112 8236 11118 8248
rect 11330 8236 11336 8248
rect 11388 8276 11394 8288
rect 11698 8276 11704 8288
rect 11388 8248 11704 8276
rect 11388 8236 11394 8248
rect 11698 8236 11704 8248
rect 11756 8236 11762 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 15838 8276 15844 8288
rect 13044 8248 15844 8276
rect 13044 8236 13050 8248
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 16117 8279 16175 8285
rect 16117 8245 16129 8279
rect 16163 8276 16175 8279
rect 16206 8276 16212 8288
rect 16163 8248 16212 8276
rect 16163 8245 16175 8248
rect 16117 8239 16175 8245
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 17218 8236 17224 8288
rect 17276 8276 17282 8288
rect 17880 8276 17908 8316
rect 18782 8304 18788 8316
rect 18840 8304 18846 8356
rect 19058 8304 19064 8356
rect 19116 8344 19122 8356
rect 20364 8344 20392 8375
rect 20898 8372 20904 8375
rect 20956 8372 20962 8424
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 22281 8415 22339 8421
rect 22281 8412 22293 8415
rect 22152 8384 22293 8412
rect 22152 8372 22158 8384
rect 22281 8381 22293 8384
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 22554 8372 22560 8424
rect 22612 8372 22618 8424
rect 22664 8421 22692 8452
rect 24302 8440 24308 8452
rect 24360 8440 24366 8492
rect 24854 8440 24860 8492
rect 24912 8480 24918 8492
rect 24912 8452 26372 8480
rect 24912 8440 24918 8452
rect 22649 8415 22707 8421
rect 22649 8381 22661 8415
rect 22695 8381 22707 8415
rect 22649 8375 22707 8381
rect 22738 8372 22744 8424
rect 22796 8372 22802 8424
rect 22925 8415 22983 8421
rect 22925 8381 22937 8415
rect 22971 8412 22983 8415
rect 23201 8415 23259 8421
rect 23201 8412 23213 8415
rect 22971 8384 23213 8412
rect 22971 8381 22983 8384
rect 22925 8375 22983 8381
rect 23201 8381 23213 8384
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 23382 8372 23388 8424
rect 23440 8372 23446 8424
rect 23658 8372 23664 8424
rect 23716 8372 23722 8424
rect 25774 8372 25780 8424
rect 25832 8372 25838 8424
rect 25869 8415 25927 8421
rect 25869 8381 25881 8415
rect 25915 8412 25927 8415
rect 26234 8412 26240 8424
rect 25915 8384 26240 8412
rect 25915 8381 25927 8384
rect 25869 8375 25927 8381
rect 26234 8372 26240 8384
rect 26292 8372 26298 8424
rect 20714 8344 20720 8356
rect 19116 8316 19334 8344
rect 20364 8316 20720 8344
rect 19116 8304 19122 8316
rect 17276 8248 17908 8276
rect 17276 8236 17282 8248
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 18141 8279 18199 8285
rect 18141 8276 18153 8279
rect 18012 8248 18153 8276
rect 18012 8236 18018 8248
rect 18141 8245 18153 8248
rect 18187 8245 18199 8279
rect 19306 8276 19334 8316
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 22419 8347 22477 8353
rect 22419 8344 22431 8347
rect 21836 8316 22431 8344
rect 21836 8276 21864 8316
rect 22419 8313 22431 8316
rect 22465 8344 22477 8347
rect 22756 8344 22784 8372
rect 24118 8344 24124 8356
rect 22465 8316 22692 8344
rect 22756 8316 24124 8344
rect 22465 8313 22477 8316
rect 22419 8307 22477 8313
rect 19306 8248 21864 8276
rect 18141 8239 18199 8245
rect 21910 8236 21916 8288
rect 21968 8276 21974 8288
rect 22005 8279 22063 8285
rect 22005 8276 22017 8279
rect 21968 8248 22017 8276
rect 21968 8236 21974 8248
rect 22005 8245 22017 8248
rect 22051 8245 22063 8279
rect 22664 8276 22692 8316
rect 24118 8304 24124 8316
rect 24176 8304 24182 8356
rect 25130 8304 25136 8356
rect 25188 8344 25194 8356
rect 26053 8347 26111 8353
rect 26053 8344 26065 8347
rect 25188 8316 26065 8344
rect 25188 8304 25194 8316
rect 26053 8313 26065 8316
rect 26099 8313 26111 8347
rect 26344 8344 26372 8452
rect 26418 8372 26424 8424
rect 26476 8412 26482 8424
rect 26528 8421 26556 8520
rect 28092 8421 28120 8588
rect 28534 8576 28540 8588
rect 28592 8576 28598 8628
rect 28994 8576 29000 8628
rect 29052 8616 29058 8628
rect 29641 8619 29699 8625
rect 29641 8616 29653 8619
rect 29052 8588 29653 8616
rect 29052 8576 29058 8588
rect 29641 8585 29653 8588
rect 29687 8585 29699 8619
rect 29641 8579 29699 8585
rect 28258 8508 28264 8560
rect 28316 8548 28322 8560
rect 28902 8548 28908 8560
rect 28316 8520 28908 8548
rect 28316 8508 28322 8520
rect 28902 8508 28908 8520
rect 28960 8548 28966 8560
rect 28960 8520 29224 8548
rect 28960 8508 28966 8520
rect 28350 8440 28356 8492
rect 28408 8480 28414 8492
rect 28626 8480 28632 8492
rect 28408 8452 28632 8480
rect 28408 8440 28414 8452
rect 28626 8440 28632 8452
rect 28684 8440 28690 8492
rect 28721 8483 28779 8489
rect 28721 8449 28733 8483
rect 28767 8480 28779 8483
rect 29086 8480 29092 8492
rect 28767 8452 29092 8480
rect 28767 8449 28779 8452
rect 28721 8443 28779 8449
rect 29086 8440 29092 8452
rect 29144 8440 29150 8492
rect 26513 8415 26571 8421
rect 26513 8412 26525 8415
rect 26476 8384 26525 8412
rect 26476 8372 26482 8384
rect 26513 8381 26525 8384
rect 26559 8381 26571 8415
rect 26513 8375 26571 8381
rect 27617 8415 27675 8421
rect 27617 8381 27629 8415
rect 27663 8412 27675 8415
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27663 8384 28089 8412
rect 27663 8381 27675 8384
rect 27617 8375 27675 8381
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 27249 8347 27307 8353
rect 27249 8344 27261 8347
rect 26344 8316 27261 8344
rect 26053 8307 26111 8313
rect 27249 8313 27261 8316
rect 27295 8344 27307 8347
rect 27632 8344 27660 8375
rect 28534 8372 28540 8424
rect 28592 8372 28598 8424
rect 28810 8372 28816 8424
rect 28868 8412 28874 8424
rect 28997 8415 29055 8421
rect 28997 8412 29009 8415
rect 28868 8384 29009 8412
rect 28868 8372 28874 8384
rect 28997 8381 29009 8384
rect 29043 8381 29055 8415
rect 29196 8412 29224 8520
rect 29196 8384 29316 8412
rect 28997 8375 29055 8381
rect 29288 8356 29316 8384
rect 29454 8372 29460 8424
rect 29512 8372 29518 8424
rect 27295 8316 27660 8344
rect 27295 8313 27307 8316
rect 27249 8307 27307 8313
rect 28442 8304 28448 8356
rect 28500 8344 28506 8356
rect 29155 8347 29213 8353
rect 29155 8344 29167 8347
rect 28500 8316 29167 8344
rect 28500 8304 28506 8316
rect 29155 8313 29167 8316
rect 29201 8344 29213 8347
rect 29201 8313 29224 8344
rect 29155 8307 29224 8313
rect 22830 8276 22836 8288
rect 22664 8248 22836 8276
rect 22005 8239 22063 8245
rect 22830 8236 22836 8248
rect 22888 8236 22894 8288
rect 23014 8236 23020 8288
rect 23072 8236 23078 8288
rect 23566 8236 23572 8288
rect 23624 8236 23630 8288
rect 28169 8279 28227 8285
rect 28169 8245 28181 8279
rect 28215 8276 28227 8279
rect 28626 8276 28632 8288
rect 28215 8248 28632 8276
rect 28215 8245 28227 8248
rect 28169 8239 28227 8245
rect 28626 8236 28632 8248
rect 28684 8236 28690 8288
rect 29196 8276 29224 8307
rect 29270 8304 29276 8356
rect 29328 8304 29334 8356
rect 29365 8347 29423 8353
rect 29365 8313 29377 8347
rect 29411 8344 29423 8347
rect 30650 8344 30656 8356
rect 29411 8316 30656 8344
rect 29411 8313 29423 8316
rect 29365 8307 29423 8313
rect 30650 8304 30656 8316
rect 30708 8304 30714 8356
rect 30742 8276 30748 8288
rect 29196 8248 30748 8276
rect 30742 8236 30748 8248
rect 30800 8236 30806 8288
rect 552 8186 31648 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 12096 8186
rect 12148 8134 12160 8186
rect 12212 8134 12224 8186
rect 12276 8134 12288 8186
rect 12340 8134 12352 8186
rect 12404 8134 19870 8186
rect 19922 8134 19934 8186
rect 19986 8134 19998 8186
rect 20050 8134 20062 8186
rect 20114 8134 20126 8186
rect 20178 8134 27644 8186
rect 27696 8134 27708 8186
rect 27760 8134 27772 8186
rect 27824 8134 27836 8186
rect 27888 8134 27900 8186
rect 27952 8134 31648 8186
rect 552 8112 31648 8134
rect 4982 8032 4988 8084
rect 5040 8032 5046 8084
rect 12618 8072 12624 8084
rect 10060 8044 12624 8072
rect 3872 8007 3930 8013
rect 3872 7973 3884 8007
rect 3918 8004 3930 8007
rect 4062 8004 4068 8016
rect 3918 7976 4068 8004
rect 3918 7973 3930 7976
rect 3872 7967 3930 7973
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3605 7939 3663 7945
rect 3605 7936 3617 7939
rect 3016 7908 3617 7936
rect 3016 7896 3022 7908
rect 3605 7905 3617 7908
rect 3651 7905 3663 7939
rect 3605 7899 3663 7905
rect 7742 7896 7748 7948
rect 7800 7896 7806 7948
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 7852 7908 8033 7936
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7852 7868 7880 7908
rect 8021 7905 8033 7908
rect 8067 7936 8079 7939
rect 8202 7936 8208 7948
rect 8067 7908 8208 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 9858 7896 9864 7948
rect 9916 7896 9922 7948
rect 10060 7945 10088 8044
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 14608 8044 14780 8072
rect 14608 8032 14614 8044
rect 10704 7976 12020 8004
rect 10704 7948 10732 7976
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 10597 7939 10655 7945
rect 10597 7936 10609 7939
rect 10192 7908 10609 7936
rect 10192 7896 10198 7908
rect 10597 7905 10609 7908
rect 10643 7936 10655 7939
rect 10686 7936 10692 7948
rect 10643 7908 10692 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11287 7908 11652 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 6880 7840 7880 7868
rect 6880 7828 6886 7840
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 11256 7868 11284 7899
rect 10284 7840 11284 7868
rect 11517 7871 11575 7877
rect 10284 7828 10290 7840
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11624 7868 11652 7908
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 11756 7908 11805 7936
rect 11756 7896 11762 7908
rect 11793 7905 11805 7908
rect 11839 7905 11851 7939
rect 11992 7936 12020 7976
rect 12066 7964 12072 8016
rect 12124 8004 12130 8016
rect 12221 8007 12279 8013
rect 12221 8004 12233 8007
rect 12124 7976 12233 8004
rect 12124 7964 12130 7976
rect 12221 7973 12233 7976
rect 12267 7973 12279 8007
rect 12221 7967 12279 7973
rect 12437 8007 12495 8013
rect 12437 7973 12449 8007
rect 12483 8004 12495 8007
rect 12526 8004 12532 8016
rect 12483 7976 12532 8004
rect 12483 7973 12495 7976
rect 12437 7967 12495 7973
rect 12526 7964 12532 7976
rect 12584 7964 12590 8016
rect 14642 7964 14648 8016
rect 14700 7964 14706 8016
rect 14752 8013 14780 8044
rect 15010 8032 15016 8084
rect 15068 8032 15074 8084
rect 15197 8075 15255 8081
rect 15197 8041 15209 8075
rect 15243 8072 15255 8075
rect 15286 8072 15292 8084
rect 15243 8044 15292 8072
rect 15243 8041 15255 8044
rect 15197 8035 15255 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 16298 8072 16304 8084
rect 15436 8044 16304 8072
rect 15436 8032 15442 8044
rect 16298 8032 16304 8044
rect 16356 8072 16362 8084
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 16356 8044 16405 8072
rect 16356 8032 16362 8044
rect 16393 8041 16405 8044
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16816 8044 16957 8072
rect 16816 8032 16822 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 16945 8035 17003 8041
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 18564 8044 18705 8072
rect 18564 8032 18570 8044
rect 18693 8041 18705 8044
rect 18739 8041 18751 8075
rect 19610 8072 19616 8084
rect 18693 8035 18751 8041
rect 18908 8044 19616 8072
rect 14737 8007 14795 8013
rect 14737 7973 14749 8007
rect 14783 7973 14795 8007
rect 14737 7967 14795 7973
rect 14875 8007 14933 8013
rect 14875 7973 14887 8007
rect 14921 8004 14933 8007
rect 15028 8004 15056 8032
rect 14921 7976 15056 8004
rect 15473 8007 15531 8013
rect 14921 7973 14933 7976
rect 14875 7967 14933 7973
rect 15473 7973 15485 8007
rect 15519 8004 15531 8007
rect 16206 8004 16212 8016
rect 15519 7976 16212 8004
rect 15519 7973 15531 7976
rect 15473 7967 15531 7973
rect 16206 7964 16212 7976
rect 16264 7964 16270 8016
rect 16482 7964 16488 8016
rect 16540 7964 16546 8016
rect 16850 7964 16856 8016
rect 16908 8004 16914 8016
rect 17497 8007 17555 8013
rect 17497 8004 17509 8007
rect 16908 7976 17509 8004
rect 16908 7964 16914 7976
rect 17497 7973 17509 7976
rect 17543 7973 17555 8007
rect 17497 7967 17555 7973
rect 17586 7964 17592 8016
rect 17644 8013 17650 8016
rect 17644 8007 17673 8013
rect 17661 7973 17673 8007
rect 17644 7967 17673 7973
rect 17644 7964 17650 7967
rect 18138 7964 18144 8016
rect 18196 7964 18202 8016
rect 18325 8007 18383 8013
rect 18325 7973 18337 8007
rect 18371 8004 18383 8007
rect 18414 8004 18420 8016
rect 18371 7976 18420 8004
rect 18371 7973 18383 7976
rect 18325 7967 18383 7973
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 11992 7908 12633 7936
rect 11793 7899 11851 7905
rect 12621 7905 12633 7908
rect 12667 7936 12679 7939
rect 13170 7936 13176 7948
rect 12667 7908 13176 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 13170 7896 13176 7908
rect 13228 7936 13234 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13228 7908 13369 7936
rect 13228 7896 13234 7908
rect 13357 7905 13369 7908
rect 13403 7936 13415 7939
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 13403 7908 13645 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13633 7905 13645 7908
rect 13679 7936 13691 7939
rect 13722 7936 13728 7948
rect 13679 7908 13728 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 14093 7939 14151 7945
rect 14093 7905 14105 7939
rect 14139 7936 14151 7939
rect 14369 7939 14427 7945
rect 14369 7936 14381 7939
rect 14139 7908 14381 7936
rect 14139 7905 14151 7908
rect 14093 7899 14151 7905
rect 14369 7905 14381 7908
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 14553 7939 14611 7945
rect 14553 7905 14565 7939
rect 14599 7905 14611 7939
rect 14553 7899 14611 7905
rect 11882 7868 11888 7880
rect 11624 7840 11888 7868
rect 11517 7831 11575 7837
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 9861 7803 9919 7809
rect 9861 7800 9873 7803
rect 8628 7772 9873 7800
rect 8628 7760 8634 7772
rect 9861 7769 9873 7772
rect 9907 7769 9919 7803
rect 11532 7800 11560 7831
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12986 7868 12992 7880
rect 12032 7840 12992 7868
rect 12032 7828 12038 7840
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 14274 7868 14280 7880
rect 13136 7840 14280 7868
rect 13136 7828 13142 7840
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 14568 7868 14596 7899
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 15286 7936 15292 7948
rect 15068 7908 15292 7936
rect 15068 7896 15074 7908
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15381 7939 15439 7945
rect 15381 7905 15393 7939
rect 15427 7905 15439 7939
rect 15381 7899 15439 7905
rect 15396 7868 15424 7899
rect 15562 7896 15568 7948
rect 15620 7896 15626 7948
rect 15654 7896 15660 7948
rect 15712 7945 15718 7948
rect 15712 7939 15741 7945
rect 15729 7905 15741 7939
rect 15712 7899 15741 7905
rect 15712 7896 15718 7899
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 16114 7936 16120 7948
rect 15896 7908 16120 7936
rect 15896 7896 15902 7908
rect 16114 7896 16120 7908
rect 16172 7896 16178 7948
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 17218 7936 17224 7948
rect 17083 7908 17224 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17313 7939 17371 7945
rect 17313 7905 17325 7939
rect 17359 7905 17371 7939
rect 17313 7899 17371 7905
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 14568 7840 15424 7868
rect 15396 7812 15424 7840
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 17129 7871 17187 7877
rect 17129 7868 17141 7871
rect 16632 7840 17141 7868
rect 16632 7828 16638 7840
rect 17129 7837 17141 7840
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 12069 7803 12127 7809
rect 12069 7800 12081 7803
rect 11532 7772 12081 7800
rect 9861 7763 9919 7769
rect 12069 7769 12081 7772
rect 12115 7769 12127 7803
rect 12069 7763 12127 7769
rect 15378 7760 15384 7812
rect 15436 7800 15442 7812
rect 17328 7800 17356 7899
rect 17420 7868 17448 7899
rect 17770 7896 17776 7948
rect 17828 7896 17834 7948
rect 18908 7945 18936 8044
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 20346 8032 20352 8084
rect 20404 8032 20410 8084
rect 22554 8072 22560 8084
rect 20732 8044 22560 8072
rect 18966 7964 18972 8016
rect 19024 7964 19030 8016
rect 20732 8013 20760 8044
rect 22554 8032 22560 8044
rect 22612 8032 22618 8084
rect 24302 8032 24308 8084
rect 24360 8032 24366 8084
rect 28442 8072 28448 8084
rect 28158 8044 28448 8072
rect 19061 8007 19119 8013
rect 19061 7973 19073 8007
rect 19107 8004 19119 8007
rect 20717 8007 20775 8013
rect 20717 8004 20729 8007
rect 19107 7976 20729 8004
rect 19107 7973 19119 7976
rect 19061 7967 19119 7973
rect 20717 7973 20729 7976
rect 20763 7973 20775 8007
rect 20717 7967 20775 7973
rect 20806 7964 20812 8016
rect 20864 8013 20870 8016
rect 20864 8007 20893 8013
rect 20881 7973 20893 8007
rect 21082 8004 21088 8016
rect 20864 7967 20893 7973
rect 21008 7976 21088 8004
rect 20864 7964 20870 7967
rect 17865 7939 17923 7945
rect 17865 7905 17877 7939
rect 17911 7936 17923 7939
rect 18877 7939 18936 7945
rect 17911 7908 18368 7936
rect 17911 7905 17923 7908
rect 17865 7899 17923 7905
rect 18340 7880 18368 7908
rect 18877 7905 18889 7939
rect 18923 7908 18936 7939
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 19150 7896 19156 7948
rect 19208 7945 19214 7948
rect 19208 7939 19237 7945
rect 19225 7905 19237 7939
rect 19208 7899 19237 7905
rect 19208 7896 19214 7899
rect 20438 7896 20444 7948
rect 20496 7936 20502 7948
rect 20533 7939 20591 7945
rect 20533 7936 20545 7939
rect 20496 7908 20545 7936
rect 20496 7896 20502 7908
rect 20533 7905 20545 7908
rect 20579 7905 20591 7939
rect 20533 7899 20591 7905
rect 20622 7896 20628 7948
rect 20680 7896 20686 7948
rect 21008 7945 21036 7976
rect 21082 7964 21088 7976
rect 21140 7964 21146 8016
rect 22278 7964 22284 8016
rect 22336 8004 22342 8016
rect 22833 8007 22891 8013
rect 22833 8004 22845 8007
rect 22336 7976 22845 8004
rect 22336 7964 22342 7976
rect 22833 7973 22845 7976
rect 22879 7973 22891 8007
rect 23566 8004 23572 8016
rect 22833 7967 22891 7973
rect 22940 7976 23572 8004
rect 20993 7939 21051 7945
rect 20993 7905 21005 7939
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 17954 7868 17960 7880
rect 17420 7840 17960 7868
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18046 7828 18052 7880
rect 18104 7828 18110 7880
rect 18322 7828 18328 7880
rect 18380 7828 18386 7880
rect 19337 7871 19395 7877
rect 19337 7837 19349 7871
rect 19383 7868 19395 7871
rect 21008 7868 21036 7899
rect 21450 7896 21456 7948
rect 21508 7896 21514 7948
rect 21634 7896 21640 7948
rect 21692 7936 21698 7948
rect 21729 7939 21787 7945
rect 21729 7936 21741 7939
rect 21692 7908 21741 7936
rect 21692 7896 21698 7908
rect 21729 7905 21741 7908
rect 21775 7905 21787 7939
rect 21729 7899 21787 7905
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 22005 7939 22063 7945
rect 22005 7936 22017 7939
rect 21876 7908 22017 7936
rect 21876 7896 21882 7908
rect 22005 7905 22017 7908
rect 22051 7905 22063 7939
rect 22005 7899 22063 7905
rect 22554 7896 22560 7948
rect 22612 7896 22618 7948
rect 22646 7896 22652 7948
rect 22704 7896 22710 7948
rect 22940 7945 22968 7976
rect 23566 7964 23572 7976
rect 23624 7964 23630 8016
rect 26418 7964 26424 8016
rect 26476 7964 26482 8016
rect 27430 7964 27436 8016
rect 27488 8004 27494 8016
rect 28158 8013 28186 8044
rect 28442 8032 28448 8044
rect 28500 8032 28506 8084
rect 28534 8032 28540 8084
rect 28592 8072 28598 8084
rect 28629 8075 28687 8081
rect 28629 8072 28641 8075
rect 28592 8044 28641 8072
rect 28592 8032 28598 8044
rect 28629 8041 28641 8044
rect 28675 8041 28687 8075
rect 28629 8035 28687 8041
rect 28810 8032 28816 8084
rect 28868 8032 28874 8084
rect 28123 8007 28186 8013
rect 28123 8004 28135 8007
rect 27488 7976 28135 8004
rect 27488 7964 27494 7976
rect 28123 7973 28135 7976
rect 28169 7976 28186 8007
rect 28169 7973 28181 7976
rect 28123 7967 28181 7973
rect 28258 7964 28264 8016
rect 28316 7964 28322 8016
rect 28353 8007 28411 8013
rect 28353 7973 28365 8007
rect 28399 8004 28411 8007
rect 28828 8004 28856 8032
rect 28966 8007 29024 8013
rect 28966 8004 28978 8007
rect 28399 7976 28580 8004
rect 28828 7976 28978 8004
rect 28399 7973 28411 7976
rect 28353 7967 28411 7973
rect 28552 7948 28580 7976
rect 28966 7973 28978 7976
rect 29012 7973 29024 8007
rect 28966 7967 29024 7973
rect 29270 7964 29276 8016
rect 29328 8004 29334 8016
rect 30742 8013 30748 8016
rect 30561 8007 30619 8013
rect 30561 8004 30573 8007
rect 29328 7976 30573 8004
rect 29328 7964 29334 7976
rect 30561 7973 30573 7976
rect 30607 7973 30619 8007
rect 30561 7967 30619 7973
rect 30699 8007 30748 8013
rect 30699 7973 30711 8007
rect 30745 7973 30748 8007
rect 30699 7967 30748 7973
rect 30742 7964 30748 7967
rect 30800 7964 30806 8016
rect 22925 7939 22983 7945
rect 22925 7905 22937 7939
rect 22971 7905 22983 7939
rect 22925 7899 22983 7905
rect 23014 7896 23020 7948
rect 23072 7936 23078 7948
rect 23181 7939 23239 7945
rect 23181 7936 23193 7939
rect 23072 7908 23193 7936
rect 23072 7896 23078 7908
rect 23181 7905 23193 7908
rect 23227 7905 23239 7939
rect 23181 7899 23239 7905
rect 26237 7939 26295 7945
rect 26237 7905 26249 7939
rect 26283 7936 26295 7939
rect 27157 7939 27215 7945
rect 27157 7936 27169 7939
rect 26283 7908 27169 7936
rect 26283 7905 26295 7908
rect 26237 7899 26295 7905
rect 27157 7905 27169 7908
rect 27203 7936 27215 7939
rect 27890 7936 27896 7948
rect 27203 7908 27896 7936
rect 27203 7905 27215 7908
rect 27157 7899 27215 7905
rect 27890 7896 27896 7908
rect 27948 7896 27954 7948
rect 28445 7939 28503 7945
rect 28445 7905 28457 7939
rect 28491 7905 28503 7939
rect 28445 7899 28503 7905
rect 19383 7840 21036 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 21545 7871 21603 7877
rect 21545 7868 21557 7871
rect 21140 7840 21557 7868
rect 21140 7828 21146 7840
rect 21545 7837 21557 7840
rect 21591 7837 21603 7871
rect 21545 7831 21603 7837
rect 27985 7871 28043 7877
rect 27985 7837 27997 7871
rect 28031 7868 28043 7871
rect 28074 7868 28080 7880
rect 28031 7840 28080 7868
rect 28031 7837 28043 7840
rect 27985 7831 28043 7837
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 28460 7868 28488 7899
rect 28534 7896 28540 7948
rect 28592 7896 28598 7948
rect 28626 7896 28632 7948
rect 28684 7936 28690 7948
rect 28721 7939 28779 7945
rect 28721 7936 28733 7939
rect 28684 7908 28733 7936
rect 28684 7896 28690 7908
rect 28721 7905 28733 7908
rect 28767 7905 28779 7939
rect 29454 7936 29460 7948
rect 28721 7899 28779 7905
rect 28828 7908 29460 7936
rect 28828 7868 28856 7908
rect 29454 7896 29460 7908
rect 29512 7936 29518 7948
rect 30377 7939 30435 7945
rect 30377 7936 30389 7939
rect 29512 7908 30389 7936
rect 29512 7896 29518 7908
rect 30377 7905 30389 7908
rect 30423 7905 30435 7939
rect 30377 7899 30435 7905
rect 30469 7939 30527 7945
rect 30469 7905 30481 7939
rect 30515 7905 30527 7939
rect 30469 7899 30527 7905
rect 30484 7868 30512 7899
rect 30834 7896 30840 7948
rect 30892 7896 30898 7948
rect 28460 7840 28856 7868
rect 30392 7840 30512 7868
rect 18064 7800 18092 7828
rect 20438 7800 20444 7812
rect 15436 7772 20444 7800
rect 15436 7760 15442 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 22094 7760 22100 7812
rect 22152 7760 22158 7812
rect 30193 7803 30251 7809
rect 30193 7800 30205 7803
rect 29656 7772 30205 7800
rect 7558 7692 7564 7744
rect 7616 7692 7622 7744
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8662 7732 8668 7744
rect 8159 7704 8668 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 10686 7692 10692 7744
rect 10744 7692 10750 7744
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10928 7704 11069 7732
rect 10928 7692 10934 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11425 7735 11483 7741
rect 11425 7701 11437 7735
rect 11471 7732 11483 7735
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11471 7704 11621 7732
rect 11471 7701 11483 7704
rect 11425 7695 11483 7701
rect 11609 7701 11621 7704
rect 11655 7701 11667 7735
rect 11609 7695 11667 7701
rect 12250 7692 12256 7744
rect 12308 7692 12314 7744
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 13722 7692 13728 7744
rect 13780 7692 13786 7744
rect 13909 7735 13967 7741
rect 13909 7701 13921 7735
rect 13955 7732 13967 7735
rect 13998 7732 14004 7744
rect 13955 7704 14004 7732
rect 13955 7701 13967 7704
rect 13909 7695 13967 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 18141 7735 18199 7741
rect 18141 7732 18153 7735
rect 18104 7704 18153 7732
rect 18104 7692 18110 7704
rect 18141 7701 18153 7704
rect 18187 7701 18199 7735
rect 18141 7695 18199 7701
rect 20622 7692 20628 7744
rect 20680 7732 20686 7744
rect 21634 7732 21640 7744
rect 20680 7704 21640 7732
rect 20680 7692 20686 7704
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 21913 7735 21971 7741
rect 21913 7701 21925 7735
rect 21959 7732 21971 7735
rect 22278 7732 22284 7744
rect 21959 7704 22284 7732
rect 21959 7701 21971 7704
rect 21913 7695 21971 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 22557 7735 22615 7741
rect 22557 7732 22569 7735
rect 22520 7704 22569 7732
rect 22520 7692 22526 7704
rect 22557 7701 22569 7704
rect 22603 7732 22615 7735
rect 23290 7732 23296 7744
rect 22603 7704 23296 7732
rect 22603 7701 22615 7704
rect 22557 7695 22615 7701
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 28626 7692 28632 7744
rect 28684 7732 28690 7744
rect 29656 7732 29684 7772
rect 30193 7769 30205 7772
rect 30239 7769 30251 7803
rect 30193 7763 30251 7769
rect 28684 7704 29684 7732
rect 28684 7692 28690 7704
rect 30098 7692 30104 7744
rect 30156 7732 30162 7744
rect 30392 7732 30420 7840
rect 30156 7704 30420 7732
rect 30156 7692 30162 7704
rect 552 7642 31648 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 11436 7642
rect 11488 7590 11500 7642
rect 11552 7590 11564 7642
rect 11616 7590 11628 7642
rect 11680 7590 11692 7642
rect 11744 7590 19210 7642
rect 19262 7590 19274 7642
rect 19326 7590 19338 7642
rect 19390 7590 19402 7642
rect 19454 7590 19466 7642
rect 19518 7590 26984 7642
rect 27036 7590 27048 7642
rect 27100 7590 27112 7642
rect 27164 7590 27176 7642
rect 27228 7590 27240 7642
rect 27292 7590 31648 7642
rect 552 7568 31648 7590
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 7800 7500 8401 7528
rect 7800 7488 7806 7500
rect 8389 7497 8401 7500
rect 8435 7497 8447 7531
rect 8389 7491 8447 7497
rect 10413 7531 10471 7537
rect 10413 7497 10425 7531
rect 10459 7528 10471 7531
rect 11514 7528 11520 7540
rect 10459 7500 11520 7528
rect 10459 7497 10471 7500
rect 10413 7491 10471 7497
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 12161 7531 12219 7537
rect 12161 7497 12173 7531
rect 12207 7528 12219 7531
rect 12526 7528 12532 7540
rect 12207 7500 12532 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 14458 7528 14464 7540
rect 13280 7500 14464 7528
rect 8205 7463 8263 7469
rect 8205 7429 8217 7463
rect 8251 7429 8263 7463
rect 8205 7423 8263 7429
rect 11977 7463 12035 7469
rect 11977 7429 11989 7463
rect 12023 7460 12035 7463
rect 12250 7460 12256 7472
rect 12023 7432 12256 7460
rect 12023 7429 12035 7432
rect 11977 7423 12035 7429
rect 8220 7392 8248 7423
rect 12250 7420 12256 7432
rect 12308 7460 12314 7472
rect 13280 7460 13308 7500
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 15105 7531 15163 7537
rect 15105 7528 15117 7531
rect 14792 7500 15117 7528
rect 14792 7488 14798 7500
rect 15105 7497 15117 7500
rect 15151 7528 15163 7531
rect 17586 7528 17592 7540
rect 15151 7500 17592 7528
rect 15151 7497 15163 7500
rect 15105 7491 15163 7497
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 17681 7531 17739 7537
rect 17681 7497 17693 7531
rect 17727 7528 17739 7531
rect 17954 7528 17960 7540
rect 17727 7500 17960 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 17954 7488 17960 7500
rect 18012 7528 18018 7540
rect 18782 7528 18788 7540
rect 18012 7500 18788 7528
rect 18012 7488 18018 7500
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 18874 7488 18880 7540
rect 18932 7488 18938 7540
rect 22554 7488 22560 7540
rect 22612 7528 22618 7540
rect 25866 7528 25872 7540
rect 22612 7500 25872 7528
rect 22612 7488 22618 7500
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 28810 7488 28816 7540
rect 28868 7488 28874 7540
rect 30098 7528 30104 7540
rect 29012 7500 30104 7528
rect 12308 7432 13308 7460
rect 12308 7420 12314 7432
rect 16390 7420 16396 7472
rect 16448 7460 16454 7472
rect 18693 7463 18751 7469
rect 18693 7460 18705 7463
rect 16448 7432 18705 7460
rect 16448 7420 16454 7432
rect 18693 7429 18705 7432
rect 18739 7429 18751 7463
rect 22370 7460 22376 7472
rect 18693 7423 18751 7429
rect 19076 7432 22376 7460
rect 8846 7392 8852 7404
rect 8220 7364 8852 7392
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6687 7296 6837 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7092 7327 7150 7333
rect 7092 7293 7104 7327
rect 7138 7324 7150 7327
rect 7558 7324 7564 7336
rect 7138 7296 7564 7324
rect 7138 7293 7150 7296
rect 7092 7287 7150 7293
rect 6564 7256 6592 7287
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 8570 7284 8576 7336
rect 8628 7284 8634 7336
rect 8680 7333 8708 7364
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9030 7352 9036 7404
rect 9088 7352 9094 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 9907 7364 10609 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 13078 7392 13084 7404
rect 11940 7364 13084 7392
rect 11940 7352 11946 7364
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13170 7352 13176 7404
rect 13228 7352 13234 7404
rect 13722 7352 13728 7404
rect 13780 7352 13786 7404
rect 17494 7352 17500 7404
rect 17552 7352 17558 7404
rect 19076 7401 19104 7432
rect 22370 7420 22376 7432
rect 22428 7420 22434 7472
rect 26326 7420 26332 7472
rect 26384 7460 26390 7472
rect 26513 7463 26571 7469
rect 26513 7460 26525 7463
rect 26384 7432 26525 7460
rect 26384 7420 26390 7432
rect 26513 7429 26525 7432
rect 26559 7429 26571 7463
rect 29012 7460 29040 7500
rect 30098 7488 30104 7500
rect 30156 7488 30162 7540
rect 26513 7423 26571 7429
rect 27172 7432 29040 7460
rect 19061 7395 19119 7401
rect 17696 7364 19012 7392
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 9766 7324 9772 7336
rect 9355 7296 9772 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7324 10011 7327
rect 10134 7324 10140 7336
rect 9999 7296 10140 7324
rect 9999 7293 10011 7296
rect 9953 7287 10011 7293
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10226 7284 10232 7336
rect 10284 7284 10290 7336
rect 10870 7333 10876 7336
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7293 10563 7327
rect 10864 7324 10876 7333
rect 10831 7296 10876 7324
rect 10505 7287 10563 7293
rect 10864 7287 10876 7296
rect 6564 7228 6868 7256
rect 6840 7200 6868 7228
rect 8754 7216 8760 7268
rect 8812 7216 8818 7268
rect 8895 7259 8953 7265
rect 8895 7225 8907 7259
rect 8941 7225 8953 7259
rect 10520 7256 10548 7287
rect 10870 7284 10876 7287
rect 10928 7284 10934 7336
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 13998 7333 14004 7336
rect 13992 7324 14004 7333
rect 13959 7296 14004 7324
rect 13992 7287 14004 7296
rect 13998 7284 14004 7287
rect 14056 7284 14062 7336
rect 15378 7284 15384 7336
rect 15436 7284 15442 7336
rect 15562 7284 15568 7336
rect 15620 7284 15626 7336
rect 15654 7284 15660 7336
rect 15712 7333 15718 7336
rect 15712 7327 15761 7333
rect 15712 7293 15715 7327
rect 15749 7293 15761 7327
rect 15712 7287 15761 7293
rect 15712 7284 15718 7287
rect 15838 7284 15844 7336
rect 15896 7324 15902 7336
rect 16022 7324 16028 7336
rect 15896 7296 16028 7324
rect 15896 7284 15902 7296
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 16206 7284 16212 7336
rect 16264 7324 16270 7336
rect 17696 7333 17724 7364
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 16264 7296 17417 7324
rect 16264 7284 16270 7296
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 17681 7327 17739 7333
rect 17681 7293 17693 7327
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 11146 7256 11152 7268
rect 10520 7228 11152 7256
rect 8895 7219 8953 7225
rect 6822 7148 6828 7200
rect 6880 7148 6886 7200
rect 8910 7188 8938 7219
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 12253 7259 12311 7265
rect 12253 7225 12265 7259
rect 12299 7225 12311 7259
rect 12253 7219 12311 7225
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8910 7160 9137 7188
rect 9125 7157 9137 7160
rect 9171 7188 9183 7191
rect 9214 7188 9220 7200
rect 9171 7160 9220 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 11054 7188 11060 7200
rect 10091 7160 11060 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 12268 7188 12296 7219
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 15197 7259 15255 7265
rect 15197 7256 15209 7259
rect 13872 7228 15209 7256
rect 13872 7216 13878 7228
rect 15197 7225 15209 7228
rect 15243 7225 15255 7259
rect 15197 7219 15255 7225
rect 15286 7216 15292 7268
rect 15344 7256 15350 7268
rect 15473 7259 15531 7265
rect 15473 7256 15485 7259
rect 15344 7228 15485 7256
rect 15344 7216 15350 7228
rect 15473 7225 15485 7228
rect 15519 7225 15531 7259
rect 15473 7219 15531 7225
rect 14550 7188 14556 7200
rect 12268 7160 14556 7188
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 15488 7188 15516 7219
rect 17696 7188 17724 7287
rect 18690 7284 18696 7336
rect 18748 7324 18754 7336
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18748 7296 18889 7324
rect 18748 7284 18754 7296
rect 18877 7293 18889 7296
rect 18923 7293 18935 7327
rect 18984 7324 19012 7364
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 22462 7392 22468 7404
rect 20763 7364 22468 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 19334 7324 19340 7336
rect 18984 7296 19340 7324
rect 18877 7287 18935 7293
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 20346 7284 20352 7336
rect 20404 7284 20410 7336
rect 19153 7259 19211 7265
rect 19153 7256 19165 7259
rect 17880 7228 19165 7256
rect 17880 7197 17908 7228
rect 19153 7225 19165 7228
rect 19199 7225 19211 7259
rect 20456 7256 20484 7355
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 24026 7352 24032 7404
rect 24084 7392 24090 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 24084 7364 24317 7392
rect 24084 7352 24090 7364
rect 24305 7361 24317 7364
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24765 7395 24823 7401
rect 24765 7361 24777 7395
rect 24811 7392 24823 7395
rect 25222 7392 25228 7404
rect 24811 7364 25228 7392
rect 24811 7361 24823 7364
rect 24765 7355 24823 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 20806 7284 20812 7336
rect 20864 7284 20870 7336
rect 24670 7284 24676 7336
rect 24728 7284 24734 7336
rect 25130 7284 25136 7336
rect 25188 7284 25194 7336
rect 27172 7333 27200 7432
rect 28261 7395 28319 7401
rect 28261 7361 28273 7395
rect 28307 7392 28319 7395
rect 28997 7395 29055 7401
rect 28997 7392 29009 7395
rect 28307 7364 29009 7392
rect 28307 7361 28319 7364
rect 28261 7355 28319 7361
rect 28997 7361 29009 7364
rect 29043 7361 29055 7395
rect 28997 7355 29055 7361
rect 25961 7327 26019 7333
rect 25961 7293 25973 7327
rect 26007 7293 26019 7327
rect 25961 7287 26019 7293
rect 26145 7327 26203 7333
rect 26145 7293 26157 7327
rect 26191 7324 26203 7327
rect 27157 7327 27215 7333
rect 27157 7324 27169 7327
rect 26191 7296 27169 7324
rect 26191 7293 26203 7296
rect 26145 7287 26203 7293
rect 27157 7293 27169 7296
rect 27203 7293 27215 7327
rect 27157 7287 27215 7293
rect 20990 7256 20996 7268
rect 20456 7228 20996 7256
rect 19153 7219 19211 7225
rect 20990 7216 20996 7228
rect 21048 7216 21054 7268
rect 22830 7256 22836 7268
rect 21560 7228 22836 7256
rect 21560 7200 21588 7228
rect 22830 7216 22836 7228
rect 22888 7216 22894 7268
rect 25976 7256 26004 7287
rect 27890 7284 27896 7336
rect 27948 7324 27954 7336
rect 28074 7324 28080 7336
rect 27948 7296 28080 7324
rect 27948 7284 27954 7296
rect 28074 7284 28080 7296
rect 28132 7324 28138 7336
rect 28169 7327 28227 7333
rect 28169 7324 28181 7327
rect 28132 7296 28181 7324
rect 28132 7284 28138 7296
rect 28169 7293 28181 7296
rect 28215 7293 28227 7327
rect 28169 7287 28227 7293
rect 28350 7284 28356 7336
rect 28408 7324 28414 7336
rect 28445 7327 28503 7333
rect 28445 7324 28457 7327
rect 28408 7296 28457 7324
rect 28408 7284 28414 7296
rect 28445 7293 28457 7296
rect 28491 7293 28503 7327
rect 28445 7287 28503 7293
rect 28626 7284 28632 7336
rect 28684 7284 28690 7336
rect 29086 7284 29092 7336
rect 29144 7324 29150 7336
rect 29253 7327 29311 7333
rect 29253 7324 29265 7327
rect 29144 7296 29265 7324
rect 29144 7284 29150 7296
rect 29253 7293 29265 7296
rect 29299 7293 29311 7327
rect 29253 7287 29311 7293
rect 26237 7259 26295 7265
rect 26237 7256 26249 7259
rect 25976 7228 26249 7256
rect 26237 7225 26249 7228
rect 26283 7256 26295 7259
rect 26602 7256 26608 7268
rect 26283 7228 26608 7256
rect 26283 7225 26295 7228
rect 26237 7219 26295 7225
rect 26602 7216 26608 7228
rect 26660 7256 26666 7268
rect 26973 7259 27031 7265
rect 26973 7256 26985 7259
rect 26660 7228 26985 7256
rect 26660 7216 26666 7228
rect 26973 7225 26985 7228
rect 27019 7225 27031 7259
rect 26973 7219 27031 7225
rect 15488 7160 17724 7188
rect 17865 7191 17923 7197
rect 17865 7157 17877 7191
rect 17911 7157 17923 7191
rect 17865 7151 17923 7157
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 21542 7188 21548 7200
rect 18012 7160 21548 7188
rect 18012 7148 18018 7160
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 22094 7148 22100 7200
rect 22152 7188 22158 7200
rect 23842 7188 23848 7200
rect 22152 7160 23848 7188
rect 22152 7148 22158 7160
rect 23842 7148 23848 7160
rect 23900 7148 23906 7200
rect 24394 7148 24400 7200
rect 24452 7188 24458 7200
rect 25041 7191 25099 7197
rect 25041 7188 25053 7191
rect 24452 7160 25053 7188
rect 24452 7148 24458 7160
rect 25041 7157 25053 7160
rect 25087 7157 25099 7191
rect 25041 7151 25099 7157
rect 25222 7148 25228 7200
rect 25280 7188 25286 7200
rect 25961 7191 26019 7197
rect 25961 7188 25973 7191
rect 25280 7160 25973 7188
rect 25280 7148 25286 7160
rect 25961 7157 25973 7160
rect 26007 7157 26019 7191
rect 25961 7151 26019 7157
rect 26694 7148 26700 7200
rect 26752 7148 26758 7200
rect 26786 7148 26792 7200
rect 26844 7148 26850 7200
rect 28534 7148 28540 7200
rect 28592 7188 28598 7200
rect 29914 7188 29920 7200
rect 28592 7160 29920 7188
rect 28592 7148 28598 7160
rect 29914 7148 29920 7160
rect 29972 7188 29978 7200
rect 30377 7191 30435 7197
rect 30377 7188 30389 7191
rect 29972 7160 30389 7188
rect 29972 7148 29978 7160
rect 30377 7157 30389 7160
rect 30423 7157 30435 7191
rect 30377 7151 30435 7157
rect 552 7098 31648 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 12096 7098
rect 12148 7046 12160 7098
rect 12212 7046 12224 7098
rect 12276 7046 12288 7098
rect 12340 7046 12352 7098
rect 12404 7046 19870 7098
rect 19922 7046 19934 7098
rect 19986 7046 19998 7098
rect 20050 7046 20062 7098
rect 20114 7046 20126 7098
rect 20178 7046 27644 7098
rect 27696 7046 27708 7098
rect 27760 7046 27772 7098
rect 27824 7046 27836 7098
rect 27888 7046 27900 7098
rect 27952 7046 31648 7098
rect 552 7024 31648 7046
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 12526 6984 12532 6996
rect 8812 6956 12532 6984
rect 8812 6944 8818 6956
rect 4246 6916 4252 6928
rect 3896 6888 4252 6916
rect 3142 6808 3148 6860
rect 3200 6848 3206 6860
rect 3896 6857 3924 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 6822 6876 6828 6928
rect 6880 6916 6886 6928
rect 7009 6919 7067 6925
rect 7009 6916 7021 6919
rect 6880 6888 7021 6916
rect 6880 6876 6886 6888
rect 7009 6885 7021 6888
rect 7055 6885 7067 6919
rect 7009 6879 7067 6885
rect 8312 6888 8524 6916
rect 3605 6851 3663 6857
rect 3605 6848 3617 6851
rect 3200 6820 3617 6848
rect 3200 6808 3206 6820
rect 3605 6817 3617 6820
rect 3651 6817 3663 6851
rect 3605 6811 3663 6817
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6817 3939 6851
rect 3881 6811 3939 6817
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6848 4215 6851
rect 5166 6848 5172 6860
rect 4203 6820 5172 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3804 6780 3832 6811
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 7098 6848 7104 6860
rect 6319 6820 7104 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 8312 6848 8340 6888
rect 7300 6820 8340 6848
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 3016 6752 4353 6780
rect 3016 6740 3022 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4890 6740 4896 6792
rect 4948 6740 4954 6792
rect 7300 6721 7328 6820
rect 8386 6808 8392 6860
rect 8444 6857 8450 6860
rect 8444 6811 8456 6857
rect 8496 6848 8524 6888
rect 8570 6876 8576 6928
rect 8628 6916 8634 6928
rect 9140 6925 9168 6956
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 16114 6984 16120 6996
rect 15988 6956 16120 6984
rect 15988 6944 15994 6956
rect 16114 6944 16120 6956
rect 16172 6984 16178 6996
rect 17773 6987 17831 6993
rect 17773 6984 17785 6987
rect 16172 6956 17785 6984
rect 16172 6944 16178 6956
rect 17773 6953 17785 6956
rect 17819 6953 17831 6987
rect 17773 6947 17831 6953
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 20901 6987 20959 6993
rect 20901 6984 20913 6987
rect 18196 6956 20913 6984
rect 18196 6944 18202 6956
rect 20901 6953 20913 6956
rect 20947 6953 20959 6987
rect 20901 6947 20959 6953
rect 22462 6944 22468 6996
rect 22520 6944 22526 6996
rect 22646 6944 22652 6996
rect 22704 6984 22710 6996
rect 23014 6984 23020 6996
rect 22704 6956 23020 6984
rect 22704 6944 22710 6956
rect 23014 6944 23020 6956
rect 23072 6984 23078 6996
rect 23072 6956 23336 6984
rect 23072 6944 23078 6956
rect 9125 6919 9183 6925
rect 8628 6888 8984 6916
rect 8628 6876 8634 6888
rect 8496 6820 8616 6848
rect 8444 6808 8450 6811
rect 8588 6780 8616 6820
rect 8662 6808 8668 6860
rect 8720 6808 8726 6860
rect 8956 6857 8984 6888
rect 9125 6885 9137 6919
rect 9171 6885 9183 6919
rect 11330 6916 11336 6928
rect 9125 6879 9183 6885
rect 10612 6888 11336 6916
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 9030 6808 9036 6860
rect 9088 6808 9094 6860
rect 9214 6808 9220 6860
rect 9272 6857 9278 6860
rect 9272 6851 9301 6857
rect 9289 6817 9301 6851
rect 9272 6811 9301 6817
rect 9272 6808 9278 6811
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10612 6857 10640 6888
rect 11330 6876 11336 6888
rect 11388 6916 11394 6928
rect 12342 6916 12348 6928
rect 11388 6888 12348 6916
rect 11388 6876 11394 6888
rect 12342 6876 12348 6888
rect 12400 6916 12406 6928
rect 13814 6916 13820 6928
rect 12400 6888 12664 6916
rect 12400 6876 12406 6888
rect 10413 6851 10471 6857
rect 10413 6848 10425 6851
rect 9732 6820 10425 6848
rect 9732 6808 9738 6820
rect 10413 6817 10425 6820
rect 10459 6817 10471 6851
rect 10413 6811 10471 6817
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10744 6820 10977 6848
rect 10744 6808 10750 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11221 6851 11279 6857
rect 11221 6848 11233 6851
rect 11112 6820 11233 6848
rect 11112 6808 11118 6820
rect 11221 6817 11233 6820
rect 11267 6817 11279 6851
rect 11221 6811 11279 6817
rect 11514 6808 11520 6860
rect 11572 6848 11578 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 11572 6820 12541 6848
rect 11572 6808 11578 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12636 6848 12664 6888
rect 13372 6888 13820 6916
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12636 6820 12725 6848
rect 12529 6811 12587 6817
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 12802 6808 12808 6860
rect 12860 6808 12866 6860
rect 13078 6808 13084 6860
rect 13136 6808 13142 6860
rect 13173 6851 13231 6857
rect 13173 6817 13185 6851
rect 13219 6848 13231 6851
rect 13372 6848 13400 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 18230 6876 18236 6928
rect 18288 6916 18294 6928
rect 18288 6888 18904 6916
rect 18288 6876 18294 6888
rect 13219 6820 13400 6848
rect 13219 6817 13231 6820
rect 13173 6811 13231 6817
rect 13446 6808 13452 6860
rect 13504 6808 13510 6860
rect 13705 6851 13763 6857
rect 13705 6848 13717 6851
rect 13556 6820 13717 6848
rect 9048 6780 9076 6808
rect 8588 6752 9076 6780
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13556 6780 13584 6820
rect 13705 6817 13717 6820
rect 13751 6817 13763 6851
rect 13705 6811 13763 6817
rect 15562 6808 15568 6860
rect 15620 6808 15626 6860
rect 18049 6851 18107 6857
rect 18049 6817 18061 6851
rect 18095 6848 18107 6851
rect 18690 6848 18696 6860
rect 18095 6820 18696 6848
rect 18095 6817 18107 6820
rect 18049 6811 18107 6817
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 13403 6752 13584 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 7285 6715 7343 6721
rect 7285 6681 7297 6715
rect 7331 6681 7343 6715
rect 7285 6675 7343 6681
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 9416 6712 9444 6743
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 15473 6783 15531 6789
rect 15473 6780 15485 6783
rect 14516 6752 15485 6780
rect 14516 6740 14522 6752
rect 15473 6749 15485 6752
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 17184 6752 17509 6780
rect 17184 6740 17190 6752
rect 17497 6749 17509 6752
rect 17543 6780 17555 6783
rect 17954 6780 17960 6792
rect 17543 6752 17960 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6780 18199 6783
rect 18187 6752 18552 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 9582 6712 9588 6724
rect 8996 6684 9588 6712
rect 8996 6672 9002 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 14829 6715 14887 6721
rect 14829 6681 14841 6715
rect 14875 6712 14887 6715
rect 15286 6712 15292 6724
rect 14875 6684 15292 6712
rect 14875 6681 14887 6684
rect 14829 6675 14887 6681
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 18524 6721 18552 6752
rect 18782 6740 18788 6792
rect 18840 6740 18846 6792
rect 18876 6780 18904 6888
rect 18966 6876 18972 6928
rect 19024 6916 19030 6928
rect 19024 6888 19472 6916
rect 19024 6876 19030 6888
rect 19061 6851 19119 6857
rect 19061 6817 19073 6851
rect 19107 6817 19119 6851
rect 19061 6811 19119 6817
rect 19076 6780 19104 6811
rect 19242 6808 19248 6860
rect 19300 6808 19306 6860
rect 19334 6808 19340 6860
rect 19392 6808 19398 6860
rect 19444 6848 19472 6888
rect 20714 6876 20720 6928
rect 20772 6916 20778 6928
rect 22005 6919 22063 6925
rect 22005 6916 22017 6919
rect 20772 6888 22017 6916
rect 20772 6876 20778 6888
rect 22005 6885 22017 6888
rect 22051 6885 22063 6919
rect 22480 6916 22508 6944
rect 23308 6916 23336 6956
rect 25866 6944 25872 6996
rect 25924 6984 25930 6996
rect 26510 6984 26516 6996
rect 25924 6956 26516 6984
rect 25924 6944 25930 6956
rect 26510 6944 26516 6956
rect 26568 6944 26574 6996
rect 23569 6919 23627 6925
rect 23569 6916 23581 6919
rect 22480 6888 23244 6916
rect 23308 6888 23581 6916
rect 22005 6879 22063 6885
rect 19610 6848 19616 6860
rect 19444 6820 19616 6848
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 21085 6851 21143 6857
rect 21085 6817 21097 6851
rect 21131 6848 21143 6851
rect 21174 6848 21180 6860
rect 21131 6820 21180 6848
rect 21131 6817 21143 6820
rect 21085 6811 21143 6817
rect 21174 6808 21180 6820
rect 21232 6808 21238 6860
rect 21266 6808 21272 6860
rect 21324 6808 21330 6860
rect 21358 6808 21364 6860
rect 21416 6848 21422 6860
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 21416 6820 22477 6848
rect 21416 6808 21422 6820
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 22738 6808 22744 6860
rect 22796 6808 22802 6860
rect 23216 6857 23244 6888
rect 23569 6885 23581 6888
rect 23615 6885 23627 6919
rect 23569 6879 23627 6885
rect 24302 6876 24308 6928
rect 24360 6876 24366 6928
rect 26326 6876 26332 6928
rect 26384 6916 26390 6928
rect 26881 6919 26939 6925
rect 26881 6916 26893 6919
rect 26384 6888 26893 6916
rect 26384 6876 26390 6888
rect 26881 6885 26893 6888
rect 26927 6885 26939 6919
rect 26881 6879 26939 6885
rect 23201 6851 23259 6857
rect 23201 6817 23213 6851
rect 23247 6817 23259 6851
rect 23201 6811 23259 6817
rect 23290 6808 23296 6860
rect 23348 6808 23354 6860
rect 23474 6808 23480 6860
rect 23532 6808 23538 6860
rect 23934 6808 23940 6860
rect 23992 6808 23998 6860
rect 24026 6808 24032 6860
rect 24084 6808 24090 6860
rect 24578 6857 24584 6860
rect 24122 6851 24180 6857
rect 24122 6817 24134 6851
rect 24168 6817 24180 6851
rect 24122 6811 24180 6817
rect 24397 6851 24455 6857
rect 24397 6817 24409 6851
rect 24443 6817 24455 6851
rect 24397 6811 24455 6817
rect 24535 6851 24584 6857
rect 24535 6817 24547 6851
rect 24581 6817 24584 6851
rect 24535 6811 24584 6817
rect 18876 6752 19104 6780
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19208 6752 19441 6780
rect 19208 6740 19214 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 22554 6780 22560 6792
rect 19429 6743 19487 6749
rect 19536 6752 22560 6780
rect 18509 6715 18567 6721
rect 18509 6681 18521 6715
rect 18555 6681 18567 6715
rect 18509 6675 18567 6681
rect 18690 6672 18696 6724
rect 18748 6712 18754 6724
rect 19536 6712 19564 6752
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6780 22707 6783
rect 22695 6752 23428 6780
rect 22695 6749 22707 6752
rect 22649 6743 22707 6749
rect 18748 6684 19564 6712
rect 19705 6715 19763 6721
rect 18748 6672 18754 6684
rect 19705 6681 19717 6715
rect 19751 6681 19763 6715
rect 19705 6675 19763 6681
rect 19889 6715 19947 6721
rect 19889 6681 19901 6715
rect 19935 6712 19947 6715
rect 19935 6684 21036 6712
rect 19935 6681 19947 6684
rect 19889 6675 19947 6681
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3568 6616 3617 6644
rect 3568 6604 3574 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 3605 6607 3663 6613
rect 4062 6604 4068 6656
rect 4120 6604 4126 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8076 6616 8769 6644
rect 8076 6604 8082 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 10781 6647 10839 6653
rect 10781 6613 10793 6647
rect 10827 6644 10839 6647
rect 11330 6644 11336 6656
rect 10827 6616 11336 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 12216 6616 12357 6644
rect 12216 6604 12222 6616
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 12345 6607 12403 6613
rect 15930 6604 15936 6656
rect 15988 6604 15994 6656
rect 18966 6604 18972 6656
rect 19024 6604 19030 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19720 6644 19748 6675
rect 19392 6616 19748 6644
rect 21008 6644 21036 6684
rect 21726 6672 21732 6724
rect 21784 6712 21790 6724
rect 22925 6715 22983 6721
rect 21784 6684 22508 6712
rect 21784 6672 21790 6684
rect 22278 6644 22284 6656
rect 21008 6616 22284 6644
rect 19392 6604 19398 6616
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 22480 6653 22508 6684
rect 22925 6681 22937 6715
rect 22971 6712 22983 6715
rect 23290 6712 23296 6724
rect 22971 6684 23296 6712
rect 22971 6681 22983 6684
rect 22925 6675 22983 6681
rect 23290 6672 23296 6684
rect 23348 6672 23354 6724
rect 23400 6712 23428 6752
rect 23750 6740 23756 6792
rect 23808 6780 23814 6792
rect 24136 6780 24164 6811
rect 23808 6752 24164 6780
rect 23808 6740 23814 6752
rect 23658 6712 23664 6724
rect 23400 6684 23664 6712
rect 23658 6672 23664 6684
rect 23716 6712 23722 6724
rect 24412 6712 24440 6811
rect 24578 6808 24584 6811
rect 24636 6808 24642 6860
rect 24949 6851 25007 6857
rect 24949 6848 24961 6851
rect 24688 6820 24961 6848
rect 24486 6712 24492 6724
rect 23716 6684 23796 6712
rect 24412 6684 24492 6712
rect 23716 6672 23722 6684
rect 22465 6647 22523 6653
rect 22465 6613 22477 6647
rect 22511 6613 22523 6647
rect 22465 6607 22523 6613
rect 22554 6604 22560 6656
rect 22612 6644 22618 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22612 6616 23029 6644
rect 22612 6604 22618 6616
rect 23017 6613 23029 6616
rect 23063 6613 23075 6647
rect 23017 6607 23075 6613
rect 23474 6604 23480 6656
rect 23532 6604 23538 6656
rect 23768 6653 23796 6684
rect 24486 6672 24492 6684
rect 24544 6672 24550 6724
rect 24688 6721 24716 6820
rect 24949 6817 24961 6820
rect 24995 6817 25007 6851
rect 24949 6811 25007 6817
rect 25038 6808 25044 6860
rect 25096 6808 25102 6860
rect 25222 6808 25228 6860
rect 25280 6808 25286 6860
rect 25317 6851 25375 6857
rect 25317 6817 25329 6851
rect 25363 6848 25375 6851
rect 26786 6848 26792 6860
rect 25363 6820 26792 6848
rect 25363 6817 25375 6820
rect 25317 6811 25375 6817
rect 26786 6808 26792 6820
rect 26844 6808 26850 6860
rect 28994 6808 29000 6860
rect 29052 6848 29058 6860
rect 29089 6851 29147 6857
rect 29089 6848 29101 6851
rect 29052 6820 29101 6848
rect 29052 6808 29058 6820
rect 29089 6817 29101 6820
rect 29135 6817 29147 6851
rect 29549 6851 29607 6857
rect 29549 6848 29561 6851
rect 29089 6811 29147 6817
rect 29472 6820 29561 6848
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6780 25835 6783
rect 26234 6780 26240 6792
rect 25823 6752 26004 6780
rect 25823 6749 25835 6752
rect 25777 6743 25835 6749
rect 24673 6715 24731 6721
rect 24673 6681 24685 6715
rect 24719 6681 24731 6715
rect 24673 6675 24731 6681
rect 23753 6647 23811 6653
rect 23753 6613 23765 6647
rect 23799 6613 23811 6647
rect 23753 6607 23811 6613
rect 23842 6604 23848 6656
rect 23900 6604 23906 6656
rect 25498 6604 25504 6656
rect 25556 6604 25562 6656
rect 25976 6644 26004 6752
rect 26068 6752 26240 6780
rect 26068 6721 26096 6752
rect 26234 6740 26240 6752
rect 26292 6780 26298 6792
rect 26973 6783 27031 6789
rect 26973 6780 26985 6783
rect 26292 6752 26985 6780
rect 26292 6740 26298 6752
rect 26973 6749 26985 6752
rect 27019 6749 27031 6783
rect 26973 6743 27031 6749
rect 29178 6740 29184 6792
rect 29236 6740 29242 6792
rect 29472 6789 29500 6820
rect 29549 6817 29561 6820
rect 29595 6817 29607 6851
rect 29549 6811 29607 6817
rect 29638 6808 29644 6860
rect 29696 6808 29702 6860
rect 29822 6808 29828 6860
rect 29880 6808 29886 6860
rect 30098 6857 30104 6860
rect 29917 6851 29975 6857
rect 29917 6817 29929 6851
rect 29963 6817 29975 6851
rect 29917 6811 29975 6817
rect 30055 6851 30104 6857
rect 30055 6817 30067 6851
rect 30101 6817 30104 6851
rect 30055 6811 30104 6817
rect 29457 6783 29515 6789
rect 29457 6749 29469 6783
rect 29503 6749 29515 6783
rect 29932 6780 29960 6811
rect 30098 6808 30104 6811
rect 30156 6808 30162 6860
rect 30374 6808 30380 6860
rect 30432 6848 30438 6860
rect 30469 6851 30527 6857
rect 30469 6848 30481 6851
rect 30432 6820 30481 6848
rect 30432 6808 30438 6820
rect 30469 6817 30481 6820
rect 30515 6817 30527 6851
rect 30469 6811 30527 6817
rect 30650 6808 30656 6860
rect 30708 6808 30714 6860
rect 30285 6783 30343 6789
rect 30285 6780 30297 6783
rect 29932 6752 30297 6780
rect 29457 6743 29515 6749
rect 30285 6749 30297 6752
rect 30331 6749 30343 6783
rect 30285 6743 30343 6749
rect 26053 6715 26111 6721
rect 26053 6681 26065 6715
rect 26099 6681 26111 6715
rect 26053 6675 26111 6681
rect 26160 6684 26556 6712
rect 26160 6644 26188 6684
rect 25976 6616 26188 6644
rect 26237 6647 26295 6653
rect 26237 6613 26249 6647
rect 26283 6644 26295 6647
rect 26326 6644 26332 6656
rect 26283 6616 26332 6644
rect 26283 6613 26295 6616
rect 26237 6607 26295 6613
rect 26326 6604 26332 6616
rect 26384 6604 26390 6656
rect 26418 6604 26424 6656
rect 26476 6604 26482 6656
rect 26528 6644 26556 6684
rect 26602 6672 26608 6724
rect 26660 6672 26666 6724
rect 27341 6715 27399 6721
rect 27341 6681 27353 6715
rect 27387 6712 27399 6715
rect 27387 6684 28120 6712
rect 27387 6681 27399 6684
rect 27341 6675 27399 6681
rect 27356 6644 27384 6675
rect 26528 6616 27384 6644
rect 27430 6604 27436 6656
rect 27488 6604 27494 6656
rect 28092 6644 28120 6684
rect 30190 6672 30196 6724
rect 30248 6672 30254 6724
rect 30374 6644 30380 6656
rect 28092 6616 30380 6644
rect 30374 6604 30380 6616
rect 30432 6604 30438 6656
rect 552 6554 31648 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 11436 6554
rect 11488 6502 11500 6554
rect 11552 6502 11564 6554
rect 11616 6502 11628 6554
rect 11680 6502 11692 6554
rect 11744 6502 19210 6554
rect 19262 6502 19274 6554
rect 19326 6502 19338 6554
rect 19390 6502 19402 6554
rect 19454 6502 19466 6554
rect 19518 6502 26984 6554
rect 27036 6502 27048 6554
rect 27100 6502 27112 6554
rect 27164 6502 27176 6554
rect 27228 6502 27240 6554
rect 27292 6502 31648 6554
rect 552 6480 31648 6502
rect 8205 6443 8263 6449
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8386 6440 8392 6452
rect 8251 6412 8392 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 9640 6412 11100 6440
rect 9640 6400 9646 6412
rect 3510 6332 3516 6384
rect 3568 6332 3574 6384
rect 11072 6372 11100 6412
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11204 6412 11529 6440
rect 11204 6400 11210 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6440 11759 6443
rect 12158 6440 12164 6452
rect 11747 6412 12164 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 12268 6412 13860 6440
rect 12268 6372 12296 6412
rect 11072 6344 12296 6372
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 12400 6344 13492 6372
rect 12400 6332 12406 6344
rect 3528 6304 3556 6332
rect 9861 6307 9919 6313
rect 3528 6276 3648 6304
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 3375 6208 3525 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3620 6236 3648 6276
rect 7300 6276 8156 6304
rect 3769 6239 3827 6245
rect 3769 6236 3781 6239
rect 3620 6208 3781 6236
rect 3513 6199 3571 6205
rect 3769 6205 3781 6208
rect 3815 6205 3827 6239
rect 3769 6199 3827 6205
rect 2038 6128 2044 6180
rect 2096 6168 2102 6180
rect 3252 6168 3280 6199
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7300 6245 7328 6276
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6880 6208 7297 6236
rect 6880 6196 6886 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7926 6196 7932 6248
rect 7984 6196 7990 6248
rect 8018 6196 8024 6248
rect 8076 6196 8082 6248
rect 8128 6236 8156 6276
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9907 6276 10057 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 12434 6304 12440 6316
rect 10045 6267 10103 6273
rect 10152 6276 12440 6304
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 8128 6208 9965 6236
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 6365 6171 6423 6177
rect 2096 6140 5212 6168
rect 2096 6128 2102 6140
rect 5184 6112 5212 6140
rect 6365 6137 6377 6171
rect 6411 6137 6423 6171
rect 6365 6131 6423 6137
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 4246 6100 4252 6112
rect 2924 6072 4252 6100
rect 2924 6060 2930 6072
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4890 6060 4896 6112
rect 4948 6060 4954 6112
rect 5166 6060 5172 6112
rect 5224 6100 5230 6112
rect 6380 6100 6408 6131
rect 7098 6128 7104 6180
rect 7156 6168 7162 6180
rect 7156 6140 8616 6168
rect 7156 6128 7162 6140
rect 8110 6100 8116 6112
rect 5224 6072 8116 6100
rect 5224 6060 5230 6072
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 8444 6072 8493 6100
rect 8444 6060 8450 6072
rect 8481 6069 8493 6072
rect 8527 6069 8539 6103
rect 8588 6100 8616 6140
rect 8662 6128 8668 6180
rect 8720 6168 8726 6180
rect 9594 6171 9652 6177
rect 9594 6168 9606 6171
rect 8720 6140 9606 6168
rect 8720 6128 8726 6140
rect 9594 6137 9606 6140
rect 9640 6137 9652 6171
rect 9594 6131 9652 6137
rect 10152 6100 10180 6276
rect 12434 6264 12440 6276
rect 12492 6304 12498 6316
rect 12492 6276 13400 6304
rect 12492 6264 12498 6276
rect 12158 6196 12164 6248
rect 12216 6196 12222 6248
rect 12526 6236 12532 6248
rect 12406 6208 12532 6236
rect 11685 6171 11743 6177
rect 11685 6137 11697 6171
rect 11731 6168 11743 6171
rect 11790 6168 11796 6180
rect 11731 6140 11796 6168
rect 11731 6137 11743 6140
rect 11685 6131 11743 6137
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 11885 6171 11943 6177
rect 11885 6137 11897 6171
rect 11931 6168 11943 6171
rect 12406 6168 12434 6208
rect 12526 6196 12532 6208
rect 12584 6236 12590 6248
rect 12802 6236 12808 6248
rect 12584 6208 12808 6236
rect 12584 6196 12590 6208
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 13372 6245 13400 6276
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6205 13415 6239
rect 13357 6199 13415 6205
rect 13464 6236 13492 6344
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 13832 6304 13860 6412
rect 18782 6400 18788 6452
rect 18840 6440 18846 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 18840 6412 19441 6440
rect 18840 6400 18846 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 20533 6443 20591 6449
rect 19576 6412 20300 6440
rect 19576 6400 19582 6412
rect 18417 6375 18475 6381
rect 18417 6341 18429 6375
rect 18463 6372 18475 6375
rect 18463 6344 19932 6372
rect 18463 6341 18475 6344
rect 18417 6335 18475 6341
rect 15010 6304 15016 6316
rect 13587 6276 15016 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 16482 6264 16488 6316
rect 16540 6264 16546 6316
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 17402 6304 17408 6316
rect 17267 6276 17408 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 17543 6276 18368 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13464 6208 13737 6236
rect 11931 6140 12434 6168
rect 12621 6171 12679 6177
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12621 6137 12633 6171
rect 12667 6168 12679 6171
rect 13170 6168 13176 6180
rect 12667 6140 13176 6168
rect 12667 6137 12679 6140
rect 12621 6131 12679 6137
rect 13170 6128 13176 6140
rect 13228 6128 13234 6180
rect 13262 6128 13268 6180
rect 13320 6168 13326 6180
rect 13464 6168 13492 6208
rect 13725 6205 13737 6208
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 15620 6208 16129 6236
rect 15620 6196 15626 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 17129 6239 17187 6245
rect 17129 6205 17141 6239
rect 17175 6236 17187 6239
rect 17865 6239 17923 6245
rect 17865 6236 17877 6239
rect 17175 6208 17877 6236
rect 17175 6205 17187 6208
rect 17129 6199 17187 6205
rect 17865 6205 17877 6208
rect 17911 6205 17923 6239
rect 17865 6199 17923 6205
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18340 6236 18368 6276
rect 18874 6264 18880 6316
rect 18932 6304 18938 6316
rect 19518 6304 19524 6316
rect 18932 6276 19524 6304
rect 18932 6264 18938 6276
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 18682 6239 18740 6245
rect 18682 6236 18694 6239
rect 18340 6208 18694 6236
rect 18233 6199 18291 6205
rect 18682 6205 18694 6208
rect 18728 6205 18740 6239
rect 18682 6199 18740 6205
rect 18786 6239 18844 6245
rect 18786 6205 18798 6239
rect 18832 6205 18844 6239
rect 19150 6236 19156 6248
rect 19208 6245 19214 6248
rect 19116 6208 19156 6236
rect 18786 6199 18844 6205
rect 17144 6168 17172 6199
rect 17218 6168 17224 6180
rect 13320 6140 13492 6168
rect 13832 6140 17080 6168
rect 17144 6140 17224 6168
rect 13320 6128 13326 6140
rect 8588 6072 10180 6100
rect 12253 6103 12311 6109
rect 8481 6063 8539 6069
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 13832 6100 13860 6140
rect 12299 6072 13860 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 13906 6060 13912 6112
rect 13964 6060 13970 6112
rect 17052 6100 17080 6140
rect 17218 6128 17224 6140
rect 17276 6128 17282 6180
rect 17310 6128 17316 6180
rect 17368 6168 17374 6180
rect 17494 6168 17500 6180
rect 17368 6140 17500 6168
rect 17368 6128 17374 6140
rect 17494 6128 17500 6140
rect 17552 6168 17558 6180
rect 18049 6171 18107 6177
rect 18049 6168 18061 6171
rect 17552 6140 18061 6168
rect 17552 6128 17558 6140
rect 18049 6137 18061 6140
rect 18095 6137 18107 6171
rect 18049 6131 18107 6137
rect 18138 6128 18144 6180
rect 18196 6128 18202 6180
rect 18248 6100 18276 6199
rect 18690 6100 18696 6112
rect 17052 6072 18696 6100
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 18801 6100 18829 6199
rect 19150 6196 19156 6208
rect 19208 6199 19216 6245
rect 19610 6236 19616 6248
rect 19260 6208 19616 6236
rect 19208 6196 19214 6199
rect 19260 6180 19288 6208
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 19702 6196 19708 6248
rect 19760 6196 19766 6248
rect 19904 6245 19932 6344
rect 19889 6239 19947 6245
rect 19889 6205 19901 6239
rect 19935 6205 19947 6239
rect 19889 6199 19947 6205
rect 19978 6196 19984 6248
rect 20036 6196 20042 6248
rect 20272 6245 20300 6412
rect 20533 6409 20545 6443
rect 20579 6440 20591 6443
rect 22002 6440 22008 6452
rect 20579 6412 22008 6440
rect 20579 6409 20591 6412
rect 20533 6403 20591 6409
rect 22002 6400 22008 6412
rect 22060 6400 22066 6452
rect 22097 6443 22155 6449
rect 22097 6409 22109 6443
rect 22143 6440 22155 6443
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 22143 6412 22385 6440
rect 22143 6409 22155 6412
rect 22097 6403 22155 6409
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 22925 6443 22983 6449
rect 22925 6440 22937 6443
rect 22612 6412 22937 6440
rect 22612 6400 22618 6412
rect 22925 6409 22937 6412
rect 22971 6409 22983 6443
rect 22925 6403 22983 6409
rect 23566 6400 23572 6452
rect 23624 6440 23630 6452
rect 26145 6443 26203 6449
rect 26145 6440 26157 6443
rect 23624 6412 26157 6440
rect 23624 6400 23630 6412
rect 26145 6409 26157 6412
rect 26191 6409 26203 6443
rect 26145 6403 26203 6409
rect 26605 6443 26663 6449
rect 26605 6409 26617 6443
rect 26651 6440 26663 6443
rect 26694 6440 26700 6452
rect 26651 6412 26700 6440
rect 26651 6409 26663 6412
rect 26605 6403 26663 6409
rect 26694 6400 26700 6412
rect 26752 6440 26758 6452
rect 26881 6443 26939 6449
rect 26881 6440 26893 6443
rect 26752 6412 26893 6440
rect 26752 6400 26758 6412
rect 26881 6409 26893 6412
rect 26927 6409 26939 6443
rect 26881 6403 26939 6409
rect 29638 6400 29644 6452
rect 29696 6400 29702 6452
rect 29822 6400 29828 6452
rect 29880 6400 29886 6452
rect 30098 6400 30104 6452
rect 30156 6400 30162 6452
rect 22278 6372 22284 6384
rect 22066 6344 22284 6372
rect 22066 6304 22094 6344
rect 22278 6332 22284 6344
rect 22336 6332 22342 6384
rect 23014 6332 23020 6384
rect 23072 6332 23078 6384
rect 23106 6332 23112 6384
rect 23164 6372 23170 6384
rect 23750 6372 23756 6384
rect 23164 6344 23756 6372
rect 23164 6332 23170 6344
rect 23750 6332 23756 6344
rect 23808 6372 23814 6384
rect 23937 6375 23995 6381
rect 23937 6372 23949 6375
rect 23808 6344 23949 6372
rect 23808 6332 23814 6344
rect 23937 6341 23949 6344
rect 23983 6341 23995 6375
rect 23937 6335 23995 6341
rect 26252 6344 27568 6372
rect 20640 6276 22094 6304
rect 22741 6307 22799 6313
rect 20257 6239 20315 6245
rect 20257 6205 20269 6239
rect 20303 6205 20315 6239
rect 20257 6199 20315 6205
rect 20346 6196 20352 6248
rect 20404 6196 20410 6248
rect 20640 6245 20668 6276
rect 22741 6273 22753 6307
rect 22787 6304 22799 6307
rect 22787 6276 25268 6304
rect 22787 6273 22799 6276
rect 22741 6267 22799 6273
rect 20625 6239 20683 6245
rect 20625 6205 20637 6239
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 22002 6196 22008 6248
rect 22060 6196 22066 6248
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6236 22155 6239
rect 22186 6236 22192 6248
rect 22143 6208 22192 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 22186 6196 22192 6208
rect 22244 6196 22250 6248
rect 22462 6196 22468 6248
rect 22520 6236 22526 6248
rect 22557 6239 22615 6245
rect 22557 6236 22569 6239
rect 22520 6208 22569 6236
rect 22520 6196 22526 6208
rect 22557 6205 22569 6208
rect 22603 6205 22615 6239
rect 22557 6199 22615 6205
rect 24029 6239 24087 6245
rect 24029 6205 24041 6239
rect 24075 6205 24087 6239
rect 24029 6199 24087 6205
rect 18966 6128 18972 6180
rect 19024 6128 19030 6180
rect 19058 6128 19064 6180
rect 19116 6128 19122 6180
rect 19242 6128 19248 6180
rect 19300 6128 19306 6180
rect 21726 6168 21732 6180
rect 19352 6140 21732 6168
rect 19150 6100 19156 6112
rect 18801 6072 19156 6100
rect 19150 6060 19156 6072
rect 19208 6060 19214 6112
rect 19352 6109 19380 6140
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 21818 6128 21824 6180
rect 21876 6128 21882 6180
rect 22370 6128 22376 6180
rect 22428 6168 22434 6180
rect 22833 6171 22891 6177
rect 22833 6168 22845 6171
rect 22428 6140 22845 6168
rect 22428 6128 22434 6140
rect 22833 6137 22845 6140
rect 22879 6137 22891 6171
rect 22833 6131 22891 6137
rect 23385 6171 23443 6177
rect 23385 6137 23397 6171
rect 23431 6168 23443 6171
rect 24044 6168 24072 6199
rect 25130 6168 25136 6180
rect 23431 6140 25136 6168
rect 23431 6137 23443 6140
rect 23385 6131 23443 6137
rect 25130 6128 25136 6140
rect 25188 6128 25194 6180
rect 25240 6168 25268 6276
rect 26142 6264 26148 6316
rect 26200 6304 26206 6316
rect 26252 6304 26280 6344
rect 26200 6276 26280 6304
rect 26513 6307 26571 6313
rect 26200 6264 26206 6276
rect 26513 6273 26525 6307
rect 26559 6304 26571 6307
rect 26559 6276 27108 6304
rect 26559 6273 26571 6276
rect 26513 6267 26571 6273
rect 26326 6196 26332 6248
rect 26384 6236 26390 6248
rect 27080 6245 27108 6276
rect 26881 6239 26939 6245
rect 26881 6236 26893 6239
rect 26384 6208 26893 6236
rect 26384 6196 26390 6208
rect 26881 6205 26893 6208
rect 26927 6205 26939 6239
rect 26881 6199 26939 6205
rect 27065 6239 27123 6245
rect 27065 6205 27077 6239
rect 27111 6236 27123 6239
rect 27430 6236 27436 6248
rect 27111 6208 27436 6236
rect 27111 6205 27123 6208
rect 27065 6199 27123 6205
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 26418 6168 26424 6180
rect 25240 6140 26424 6168
rect 26418 6128 26424 6140
rect 26476 6168 26482 6180
rect 26605 6171 26663 6177
rect 26605 6168 26617 6171
rect 26476 6140 26617 6168
rect 26476 6128 26482 6140
rect 26605 6137 26617 6140
rect 26651 6137 26663 6171
rect 27540 6168 27568 6344
rect 29288 6276 29960 6304
rect 29288 6245 29316 6276
rect 29932 6248 29960 6276
rect 29273 6239 29331 6245
rect 29273 6205 29285 6239
rect 29319 6205 29331 6239
rect 29273 6199 29331 6205
rect 29457 6239 29515 6245
rect 29457 6205 29469 6239
rect 29503 6236 29515 6239
rect 29733 6239 29791 6245
rect 29733 6236 29745 6239
rect 29503 6208 29745 6236
rect 29503 6205 29515 6208
rect 29457 6199 29515 6205
rect 29733 6205 29745 6208
rect 29779 6205 29791 6239
rect 29733 6199 29791 6205
rect 29472 6168 29500 6199
rect 29914 6196 29920 6248
rect 29972 6196 29978 6248
rect 30009 6239 30067 6245
rect 30009 6205 30021 6239
rect 30055 6205 30067 6239
rect 30009 6199 30067 6205
rect 30193 6239 30251 6245
rect 30193 6205 30205 6239
rect 30239 6236 30251 6239
rect 30650 6236 30656 6248
rect 30239 6208 30656 6236
rect 30239 6205 30251 6208
rect 30193 6199 30251 6205
rect 27540 6140 29500 6168
rect 30024 6168 30052 6199
rect 30650 6196 30656 6208
rect 30708 6196 30714 6248
rect 30374 6168 30380 6180
rect 30024 6140 30380 6168
rect 26605 6131 26663 6137
rect 30374 6128 30380 6140
rect 30432 6128 30438 6180
rect 19337 6103 19395 6109
rect 19337 6069 19349 6103
rect 19383 6069 19395 6103
rect 19337 6063 19395 6069
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 19668 6072 20085 6100
rect 19668 6060 19674 6072
rect 20073 6069 20085 6072
rect 20119 6069 20131 6103
rect 20073 6063 20131 6069
rect 22281 6103 22339 6109
rect 22281 6069 22293 6103
rect 22327 6100 22339 6103
rect 23106 6100 23112 6112
rect 22327 6072 23112 6100
rect 22327 6069 22339 6072
rect 22281 6063 22339 6069
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 23198 6060 23204 6112
rect 23256 6100 23262 6112
rect 23842 6100 23848 6112
rect 23256 6072 23848 6100
rect 23256 6060 23262 6072
rect 23842 6060 23848 6072
rect 23900 6060 23906 6112
rect 26694 6060 26700 6112
rect 26752 6060 26758 6112
rect 552 6010 31648 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 12096 6010
rect 12148 5958 12160 6010
rect 12212 5958 12224 6010
rect 12276 5958 12288 6010
rect 12340 5958 12352 6010
rect 12404 5958 19870 6010
rect 19922 5958 19934 6010
rect 19986 5958 19998 6010
rect 20050 5958 20062 6010
rect 20114 5958 20126 6010
rect 20178 5958 27644 6010
rect 27696 5958 27708 6010
rect 27760 5958 27772 6010
rect 27824 5958 27836 6010
rect 27888 5958 27900 6010
rect 27952 5958 31648 6010
rect 552 5936 31648 5958
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 3142 5896 3148 5908
rect 2731 5868 3148 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 4890 5896 4896 5908
rect 3344 5868 4896 5896
rect 2866 5720 2872 5772
rect 2924 5720 2930 5772
rect 2958 5720 2964 5772
rect 3016 5720 3022 5772
rect 3344 5769 3372 5868
rect 4890 5856 4896 5868
rect 4948 5896 4954 5908
rect 8205 5899 8263 5905
rect 4948 5868 6960 5896
rect 4948 5856 4954 5868
rect 4062 5828 4068 5840
rect 3712 5800 4068 5828
rect 3712 5769 3740 5800
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 4154 5788 4160 5840
rect 4212 5788 4218 5840
rect 4246 5788 4252 5840
rect 4304 5828 4310 5840
rect 6932 5837 6960 5868
rect 8205 5865 8217 5899
rect 8251 5896 8263 5899
rect 8662 5896 8668 5908
rect 8251 5868 8668 5896
rect 8251 5865 8263 5868
rect 8205 5859 8263 5865
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9582 5896 9588 5908
rect 8812 5868 9588 5896
rect 8812 5856 8818 5868
rect 6701 5831 6759 5837
rect 6701 5828 6713 5831
rect 4304 5800 6713 5828
rect 4304 5788 4310 5800
rect 6701 5797 6713 5800
rect 6747 5797 6759 5831
rect 6701 5791 6759 5797
rect 6917 5831 6975 5837
rect 6917 5797 6929 5831
rect 6963 5797 6975 5831
rect 6917 5791 6975 5797
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 8864 5837 8892 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 15838 5896 15844 5908
rect 12406 5868 15844 5896
rect 8849 5831 8907 5837
rect 8444 5800 8800 5828
rect 8444 5788 8450 5800
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5729 3387 5763
rect 3329 5723 3387 5729
rect 3697 5763 3755 5769
rect 3697 5729 3709 5763
rect 3743 5729 3755 5763
rect 3953 5763 4011 5769
rect 3953 5760 3965 5763
rect 3697 5723 3755 5729
rect 3804 5732 3965 5760
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2372 5664 2697 5692
rect 2372 5652 2378 5664
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3160 5624 3188 5655
rect 3234 5652 3240 5704
rect 3292 5652 3298 5704
rect 3418 5652 3424 5704
rect 3476 5652 3482 5704
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 3804 5692 3832 5732
rect 3953 5729 3965 5732
rect 3999 5729 4011 5763
rect 4172 5760 4200 5788
rect 8772 5772 8800 5800
rect 8849 5797 8861 5831
rect 8895 5797 8907 5831
rect 12406 5828 12434 5868
rect 8849 5791 8907 5797
rect 9140 5800 12434 5828
rect 5353 5763 5411 5769
rect 5353 5760 5365 5763
rect 4172 5732 5365 5760
rect 3953 5723 4011 5729
rect 5353 5729 5365 5732
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 7926 5720 7932 5772
rect 7984 5720 7990 5772
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8067 5732 8493 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8481 5729 8493 5732
rect 8527 5729 8539 5763
rect 8481 5723 8539 5729
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 8665 5763 8723 5769
rect 8665 5760 8677 5763
rect 8628 5732 8677 5760
rect 8628 5720 8634 5732
rect 8665 5729 8677 5732
rect 8711 5729 8723 5763
rect 8665 5723 8723 5729
rect 3568 5664 3832 5692
rect 5629 5695 5687 5701
rect 3568 5652 3574 5664
rect 5629 5661 5641 5695
rect 5675 5692 5687 5695
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5675 5664 5825 5692
rect 5675 5661 5687 5664
rect 5629 5655 5687 5661
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 6328 5664 6377 5692
rect 6328 5652 6334 5664
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 3160 5596 3740 5624
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 3384 5528 3617 5556
rect 3384 5516 3390 5528
rect 3605 5525 3617 5528
rect 3651 5525 3663 5559
rect 3712 5556 3740 5596
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 5169 5627 5227 5633
rect 5169 5624 5181 5627
rect 4764 5596 5181 5624
rect 4764 5584 4770 5596
rect 5169 5593 5181 5596
rect 5215 5593 5227 5627
rect 5902 5624 5908 5636
rect 5169 5587 5227 5593
rect 5460 5596 5908 5624
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 3712 5528 5089 5556
rect 3605 5519 3663 5525
rect 5077 5525 5089 5528
rect 5123 5556 5135 5559
rect 5460 5556 5488 5596
rect 5902 5584 5908 5596
rect 5960 5624 5966 5636
rect 8680 5624 8708 5723
rect 8754 5720 8760 5772
rect 8812 5720 8818 5772
rect 9140 5769 9168 5800
rect 12986 5788 12992 5840
rect 13044 5828 13050 5840
rect 13630 5828 13636 5840
rect 13044 5800 13636 5828
rect 13044 5788 13050 5800
rect 13630 5788 13636 5800
rect 13688 5788 13694 5840
rect 8967 5763 9025 5769
rect 8967 5729 8979 5763
rect 9013 5760 9025 5763
rect 9125 5763 9183 5769
rect 9013 5729 9030 5760
rect 8967 5723 9030 5729
rect 9125 5729 9137 5763
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 9002 5692 9030 5723
rect 9398 5720 9404 5772
rect 9456 5720 9462 5772
rect 9490 5720 9496 5772
rect 9548 5720 9554 5772
rect 9582 5720 9588 5772
rect 9640 5720 9646 5772
rect 9703 5763 9761 5769
rect 9703 5760 9715 5763
rect 9692 5729 9715 5760
rect 9749 5729 9761 5763
rect 9692 5723 9761 5729
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5760 9919 5763
rect 10042 5760 10048 5772
rect 9907 5732 10048 5760
rect 9907 5729 9919 5732
rect 9861 5723 9919 5729
rect 9214 5692 9220 5704
rect 9002 5664 9220 5692
rect 9214 5652 9220 5664
rect 9272 5692 9278 5704
rect 9692 5692 9720 5723
rect 10042 5720 10048 5732
rect 10100 5760 10106 5772
rect 11149 5763 11207 5769
rect 11149 5760 11161 5763
rect 10100 5732 11161 5760
rect 10100 5720 10106 5732
rect 11149 5729 11161 5732
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 11238 5720 11244 5772
rect 11296 5760 11302 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11296 5732 11345 5760
rect 11296 5720 11302 5732
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 9272 5664 9720 5692
rect 12912 5692 12940 5723
rect 13262 5720 13268 5772
rect 13320 5720 13326 5772
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 13372 5732 13737 5760
rect 13170 5692 13176 5704
rect 12912 5664 13176 5692
rect 9272 5652 9278 5664
rect 13170 5652 13176 5664
rect 13228 5692 13234 5704
rect 13372 5692 13400 5732
rect 13725 5729 13737 5732
rect 13771 5729 13783 5763
rect 13725 5723 13783 5729
rect 13228 5664 13400 5692
rect 13449 5695 13507 5701
rect 13228 5652 13234 5664
rect 13449 5661 13461 5695
rect 13495 5692 13507 5695
rect 13832 5692 13860 5868
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 19702 5896 19708 5908
rect 18892 5868 19708 5896
rect 18892 5769 18920 5868
rect 19702 5856 19708 5868
rect 19760 5856 19766 5908
rect 19794 5856 19800 5908
rect 19852 5896 19858 5908
rect 20346 5896 20352 5908
rect 19852 5868 20352 5896
rect 19852 5856 19858 5868
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 21358 5856 21364 5908
rect 21416 5856 21422 5908
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 21836 5868 21925 5896
rect 19610 5828 19616 5840
rect 19444 5800 19616 5828
rect 19444 5769 19472 5800
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 21836 5837 21864 5868
rect 21913 5865 21925 5868
rect 21959 5865 21971 5899
rect 22922 5896 22928 5908
rect 21913 5859 21971 5865
rect 22112 5868 22928 5896
rect 21821 5831 21879 5837
rect 21821 5797 21833 5831
rect 21867 5797 21879 5831
rect 21821 5791 21879 5797
rect 22112 5772 22140 5868
rect 22922 5856 22928 5868
rect 22980 5856 22986 5908
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 23532 5868 23857 5896
rect 23532 5856 23538 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 23845 5859 23903 5865
rect 22278 5828 22284 5840
rect 22204 5800 22284 5828
rect 18877 5763 18935 5769
rect 18877 5729 18889 5763
rect 18923 5729 18935 5763
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18877 5723 18935 5729
rect 18984 5732 19257 5760
rect 18984 5704 19012 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19429 5763 19487 5769
rect 19429 5729 19441 5763
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 19521 5763 19579 5769
rect 19521 5729 19533 5763
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 19705 5763 19763 5769
rect 19705 5729 19717 5763
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 21545 5763 21603 5769
rect 21545 5729 21557 5763
rect 21591 5760 21603 5763
rect 22002 5760 22008 5772
rect 21591 5732 22008 5760
rect 21591 5729 21603 5732
rect 21545 5723 21603 5729
rect 13495 5664 13860 5692
rect 13495 5661 13507 5664
rect 13449 5655 13507 5661
rect 18966 5652 18972 5704
rect 19024 5652 19030 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5661 19119 5695
rect 19061 5655 19119 5661
rect 9398 5624 9404 5636
rect 5960 5596 6776 5624
rect 8680 5596 9404 5624
rect 5960 5584 5966 5596
rect 5123 5528 5488 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 6748 5565 6776 5596
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 13633 5627 13691 5633
rect 13633 5624 13645 5627
rect 12952 5596 13645 5624
rect 12952 5584 12958 5596
rect 13633 5593 13645 5596
rect 13679 5593 13691 5627
rect 13633 5587 13691 5593
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 19076 5624 19104 5655
rect 19150 5652 19156 5704
rect 19208 5692 19214 5704
rect 19536 5692 19564 5723
rect 19720 5692 19748 5723
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 22094 5720 22100 5772
rect 22152 5720 22158 5772
rect 19208 5664 19564 5692
rect 19628 5664 19748 5692
rect 21729 5695 21787 5701
rect 19208 5652 19214 5664
rect 19242 5624 19248 5636
rect 16540 5596 19012 5624
rect 19076 5596 19248 5624
rect 16540 5584 16546 5596
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 5592 5528 6561 5556
rect 5592 5516 5598 5528
rect 6549 5525 6561 5528
rect 6595 5525 6607 5559
rect 6549 5519 6607 5525
rect 6733 5559 6791 5565
rect 6733 5525 6745 5559
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9217 5559 9275 5565
rect 9217 5556 9229 5559
rect 9180 5528 9229 5556
rect 9180 5516 9186 5528
rect 9217 5525 9229 5528
rect 9263 5525 9275 5559
rect 9217 5519 9275 5525
rect 11517 5559 11575 5565
rect 11517 5525 11529 5559
rect 11563 5556 11575 5559
rect 12158 5556 12164 5568
rect 11563 5528 12164 5556
rect 11563 5525 11575 5528
rect 11517 5519 11575 5525
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 13078 5516 13084 5568
rect 13136 5516 13142 5568
rect 18690 5516 18696 5568
rect 18748 5516 18754 5568
rect 18984 5556 19012 5596
rect 19242 5584 19248 5596
rect 19300 5584 19306 5636
rect 19334 5584 19340 5636
rect 19392 5624 19398 5636
rect 19628 5624 19656 5664
rect 21729 5661 21741 5695
rect 21775 5692 21787 5695
rect 21818 5692 21824 5704
rect 21775 5664 21824 5692
rect 21775 5661 21787 5664
rect 21729 5655 21787 5661
rect 21818 5652 21824 5664
rect 21876 5692 21882 5704
rect 22204 5692 22232 5800
rect 22278 5788 22284 5800
rect 22336 5788 22342 5840
rect 22370 5788 22376 5840
rect 22428 5788 22434 5840
rect 23014 5788 23020 5840
rect 23072 5828 23078 5840
rect 23658 5828 23664 5840
rect 23072 5800 23428 5828
rect 23072 5788 23078 5800
rect 22465 5763 22523 5769
rect 22465 5729 22477 5763
rect 22511 5729 22523 5763
rect 22465 5723 22523 5729
rect 21876 5664 22232 5692
rect 22281 5695 22339 5701
rect 21876 5652 21882 5664
rect 22281 5661 22293 5695
rect 22327 5692 22339 5695
rect 22370 5692 22376 5704
rect 22327 5664 22376 5692
rect 22327 5661 22339 5664
rect 22281 5655 22339 5661
rect 22370 5652 22376 5664
rect 22428 5652 22434 5704
rect 22480 5692 22508 5723
rect 22646 5720 22652 5772
rect 22704 5720 22710 5772
rect 23198 5760 23204 5772
rect 22756 5732 23204 5760
rect 22756 5692 22784 5732
rect 23198 5720 23204 5732
rect 23256 5720 23262 5772
rect 23293 5763 23351 5769
rect 23293 5729 23305 5763
rect 23339 5729 23351 5763
rect 23293 5723 23351 5729
rect 22480 5664 22784 5692
rect 22922 5652 22928 5704
rect 22980 5652 22986 5704
rect 19392 5596 19656 5624
rect 19705 5627 19763 5633
rect 19392 5584 19398 5596
rect 19705 5593 19717 5627
rect 19751 5624 19763 5627
rect 23308 5624 23336 5723
rect 23400 5692 23428 5800
rect 23492 5800 23664 5828
rect 23492 5769 23520 5800
rect 23658 5788 23664 5800
rect 23716 5788 23722 5840
rect 23934 5788 23940 5840
rect 23992 5828 23998 5840
rect 24305 5831 24363 5837
rect 23992 5800 24164 5828
rect 23992 5788 23998 5800
rect 23477 5763 23535 5769
rect 23477 5729 23489 5763
rect 23523 5729 23535 5763
rect 23477 5723 23535 5729
rect 23566 5720 23572 5772
rect 23624 5720 23630 5772
rect 24026 5720 24032 5772
rect 24084 5720 24090 5772
rect 24136 5760 24164 5800
rect 24305 5797 24317 5831
rect 24351 5828 24363 5831
rect 24946 5828 24952 5840
rect 24351 5800 24952 5828
rect 24351 5797 24363 5800
rect 24305 5791 24363 5797
rect 24946 5788 24952 5800
rect 25004 5788 25010 5840
rect 26602 5788 26608 5840
rect 26660 5828 26666 5840
rect 26660 5800 28304 5828
rect 26660 5788 26666 5800
rect 24394 5760 24400 5772
rect 24136 5732 24400 5760
rect 24394 5720 24400 5732
rect 24452 5720 24458 5772
rect 24581 5763 24639 5769
rect 24581 5729 24593 5763
rect 24627 5760 24639 5763
rect 24670 5760 24676 5772
rect 24627 5732 24676 5760
rect 24627 5729 24639 5732
rect 24581 5723 24639 5729
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 25406 5720 25412 5772
rect 25464 5720 25470 5772
rect 25501 5763 25559 5769
rect 25501 5729 25513 5763
rect 25547 5760 25559 5763
rect 26050 5760 26056 5772
rect 25547 5732 26056 5760
rect 25547 5729 25559 5732
rect 25501 5723 25559 5729
rect 26050 5720 26056 5732
rect 26108 5720 26114 5772
rect 28077 5763 28135 5769
rect 28077 5729 28089 5763
rect 28123 5760 28135 5763
rect 28166 5760 28172 5772
rect 28123 5732 28172 5760
rect 28123 5729 28135 5732
rect 28077 5723 28135 5729
rect 28166 5720 28172 5732
rect 28224 5720 28230 5772
rect 28276 5769 28304 5800
rect 28626 5788 28632 5840
rect 28684 5828 28690 5840
rect 28905 5831 28963 5837
rect 28905 5828 28917 5831
rect 28684 5800 28917 5828
rect 28684 5788 28690 5800
rect 28905 5797 28917 5800
rect 28951 5797 28963 5831
rect 28905 5791 28963 5797
rect 28994 5788 29000 5840
rect 29052 5828 29058 5840
rect 29365 5831 29423 5837
rect 29365 5828 29377 5831
rect 29052 5800 29377 5828
rect 29052 5788 29058 5800
rect 29365 5797 29377 5800
rect 29411 5797 29423 5831
rect 29365 5791 29423 5797
rect 28261 5763 28319 5769
rect 28261 5729 28273 5763
rect 28307 5760 28319 5763
rect 28442 5760 28448 5772
rect 28307 5732 28448 5760
rect 28307 5729 28319 5732
rect 28261 5723 28319 5729
rect 28442 5720 28448 5732
rect 28500 5720 28506 5772
rect 28718 5720 28724 5772
rect 28776 5760 28782 5772
rect 29181 5763 29239 5769
rect 29181 5760 29193 5763
rect 28776 5732 29193 5760
rect 28776 5720 28782 5732
rect 29181 5729 29193 5732
rect 29227 5729 29239 5763
rect 29181 5723 29239 5729
rect 23400 5664 24072 5692
rect 19751 5596 23336 5624
rect 19751 5593 19763 5596
rect 19705 5587 19763 5593
rect 21358 5556 21364 5568
rect 18984 5528 21364 5556
rect 21358 5516 21364 5528
rect 21416 5516 21422 5568
rect 21560 5565 21588 5596
rect 23474 5584 23480 5636
rect 23532 5624 23538 5636
rect 23934 5624 23940 5636
rect 23532 5596 23940 5624
rect 23532 5584 23538 5596
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 21545 5559 21603 5565
rect 21545 5525 21557 5559
rect 21591 5525 21603 5559
rect 21545 5519 21603 5525
rect 21726 5516 21732 5568
rect 21784 5556 21790 5568
rect 22097 5559 22155 5565
rect 22097 5556 22109 5559
rect 21784 5528 22109 5556
rect 21784 5516 21790 5528
rect 22097 5525 22109 5528
rect 22143 5556 22155 5559
rect 22186 5556 22192 5568
rect 22143 5528 22192 5556
rect 22143 5525 22155 5528
rect 22097 5519 22155 5525
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 22738 5516 22744 5568
rect 22796 5516 22802 5568
rect 22833 5559 22891 5565
rect 22833 5525 22845 5559
rect 22879 5556 22891 5559
rect 22922 5556 22928 5568
rect 22879 5528 22928 5556
rect 22879 5525 22891 5528
rect 22833 5519 22891 5525
rect 22922 5516 22928 5528
rect 22980 5516 22986 5568
rect 23198 5516 23204 5568
rect 23256 5516 23262 5568
rect 23290 5516 23296 5568
rect 23348 5516 23354 5568
rect 23750 5516 23756 5568
rect 23808 5516 23814 5568
rect 24044 5565 24072 5664
rect 24210 5652 24216 5704
rect 24268 5652 24274 5704
rect 28534 5584 28540 5636
rect 28592 5584 28598 5636
rect 24029 5559 24087 5565
rect 24029 5525 24041 5559
rect 24075 5525 24087 5559
rect 24029 5519 24087 5525
rect 24302 5516 24308 5568
rect 24360 5556 24366 5568
rect 24397 5559 24455 5565
rect 24397 5556 24409 5559
rect 24360 5528 24409 5556
rect 24360 5516 24366 5528
rect 24397 5525 24409 5528
rect 24443 5525 24455 5559
rect 24397 5519 24455 5525
rect 28445 5559 28503 5565
rect 28445 5525 28457 5559
rect 28491 5556 28503 5559
rect 28905 5559 28963 5565
rect 28905 5556 28917 5559
rect 28491 5528 28917 5556
rect 28491 5525 28503 5528
rect 28445 5519 28503 5525
rect 28905 5525 28917 5528
rect 28951 5525 28963 5559
rect 28905 5519 28963 5525
rect 29086 5516 29092 5568
rect 29144 5516 29150 5568
rect 29546 5516 29552 5568
rect 29604 5516 29610 5568
rect 552 5466 31648 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 11436 5466
rect 11488 5414 11500 5466
rect 11552 5414 11564 5466
rect 11616 5414 11628 5466
rect 11680 5414 11692 5466
rect 11744 5414 19210 5466
rect 19262 5414 19274 5466
rect 19326 5414 19338 5466
rect 19390 5414 19402 5466
rect 19454 5414 19466 5466
rect 19518 5414 26984 5466
rect 27036 5414 27048 5466
rect 27100 5414 27112 5466
rect 27164 5414 27176 5466
rect 27228 5414 27240 5466
rect 27292 5414 31648 5466
rect 552 5392 31648 5414
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3602 5352 3608 5364
rect 3476 5324 3608 5352
rect 3476 5312 3482 5324
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 5626 5352 5632 5364
rect 5552 5324 5632 5352
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 5552 5225 5580 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 11388 5324 11621 5352
rect 11388 5312 11394 5324
rect 11609 5321 11621 5324
rect 11655 5321 11667 5355
rect 11609 5315 11667 5321
rect 12158 5312 12164 5364
rect 12216 5312 12222 5364
rect 12526 5312 12532 5364
rect 12584 5361 12590 5364
rect 12584 5352 12596 5361
rect 12584 5324 12629 5352
rect 12584 5315 12596 5324
rect 12584 5312 12590 5315
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 13136 5324 13277 5352
rect 13136 5312 13142 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 13906 5312 13912 5364
rect 13964 5312 13970 5364
rect 14277 5355 14335 5361
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 14458 5352 14464 5364
rect 14323 5324 14464 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 21453 5355 21511 5361
rect 21453 5321 21465 5355
rect 21499 5352 21511 5355
rect 21726 5352 21732 5364
rect 21499 5324 21732 5352
rect 21499 5321 21511 5324
rect 21453 5315 21511 5321
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 22557 5355 22615 5361
rect 22557 5352 22569 5355
rect 22336 5324 22569 5352
rect 22336 5312 22342 5324
rect 22557 5321 22569 5324
rect 22603 5321 22615 5355
rect 22557 5315 22615 5321
rect 23385 5355 23443 5361
rect 23385 5321 23397 5355
rect 23431 5352 23443 5355
rect 23750 5352 23756 5364
rect 23431 5324 23756 5352
rect 23431 5321 23443 5324
rect 23385 5315 23443 5321
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 24581 5355 24639 5361
rect 24581 5352 24593 5355
rect 24268 5324 24593 5352
rect 24268 5312 24274 5324
rect 24581 5321 24593 5324
rect 24627 5321 24639 5355
rect 24581 5315 24639 5321
rect 24762 5312 24768 5364
rect 24820 5352 24826 5364
rect 24857 5355 24915 5361
rect 24857 5352 24869 5355
rect 24820 5324 24869 5352
rect 24820 5312 24826 5324
rect 24857 5321 24869 5324
rect 24903 5321 24915 5355
rect 24857 5315 24915 5321
rect 28166 5312 28172 5364
rect 28224 5352 28230 5364
rect 28629 5355 28687 5361
rect 28224 5324 28304 5352
rect 28224 5312 28230 5324
rect 7926 5244 7932 5296
rect 7984 5284 7990 5296
rect 12345 5287 12403 5293
rect 12345 5284 12357 5287
rect 7984 5256 9352 5284
rect 7984 5244 7990 5256
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 6270 5216 6276 5228
rect 5868 5188 6276 5216
rect 5868 5176 5874 5188
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 9324 5225 9352 5256
rect 11716 5256 12357 5284
rect 11716 5225 11744 5256
rect 12345 5253 12357 5256
rect 12391 5253 12403 5287
rect 14093 5287 14151 5293
rect 14093 5284 14105 5287
rect 12345 5247 12403 5253
rect 13372 5256 14105 5284
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 9309 5219 9367 5225
rect 6779 5188 8432 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 1673 5151 1731 5157
rect 1673 5148 1685 5151
rect 1535 5120 1685 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 1673 5117 1685 5120
rect 1719 5117 1731 5151
rect 1673 5111 1731 5117
rect 1412 5012 1440 5111
rect 3418 5108 3424 5160
rect 3476 5108 3482 5160
rect 3688 5151 3746 5157
rect 3688 5117 3700 5151
rect 3734 5148 3746 5151
rect 4706 5148 4712 5160
rect 3734 5120 4712 5148
rect 3734 5117 3746 5120
rect 3688 5111 3746 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 1946 5089 1952 5092
rect 1940 5043 1952 5089
rect 1946 5040 1952 5043
rect 2004 5040 2010 5092
rect 3234 5080 3240 5092
rect 3068 5052 3240 5080
rect 2038 5012 2044 5024
rect 1412 4984 2044 5012
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 3068 5021 3096 5052
rect 3234 5040 3240 5052
rect 3292 5080 3298 5092
rect 3786 5080 3792 5092
rect 3292 5052 3792 5080
rect 3292 5040 3298 5052
rect 3786 5040 3792 5052
rect 3844 5080 3850 5092
rect 5092 5080 5120 5111
rect 5902 5108 5908 5160
rect 5960 5157 5966 5160
rect 5960 5151 5988 5157
rect 5976 5117 5988 5151
rect 5960 5111 5988 5117
rect 5960 5108 5966 5111
rect 6086 5108 6092 5160
rect 6144 5108 6150 5160
rect 8110 5108 8116 5160
rect 8168 5108 8174 5160
rect 8404 5157 8432 5188
rect 9309 5185 9321 5219
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 12986 5216 12992 5228
rect 11701 5179 11759 5185
rect 11992 5188 12992 5216
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 8846 5108 8852 5160
rect 8904 5108 8910 5160
rect 9122 5108 9128 5160
rect 9180 5108 9186 5160
rect 11146 5108 11152 5160
rect 11204 5108 11210 5160
rect 11992 5157 12020 5188
rect 12986 5176 12992 5188
rect 13044 5216 13050 5228
rect 13372 5225 13400 5256
rect 14093 5253 14105 5256
rect 14139 5253 14151 5287
rect 18322 5284 18328 5296
rect 14093 5247 14151 5253
rect 15948 5256 18328 5284
rect 13357 5219 13415 5225
rect 13044 5188 13124 5216
rect 13044 5176 13050 5188
rect 11425 5151 11483 5157
rect 11425 5117 11437 5151
rect 11471 5117 11483 5151
rect 11425 5111 11483 5117
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12434 5148 12440 5160
rect 12299 5120 12440 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 3844 5052 5120 5080
rect 8481 5083 8539 5089
rect 3844 5040 3850 5052
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 9490 5080 9496 5092
rect 8527 5052 9496 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 11440 5080 11468 5111
rect 11992 5080 12020 5111
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 13096 5157 13124 5188
rect 13357 5185 13369 5219
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15252 5188 15853 5216
rect 15252 5176 15258 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 13081 5151 13139 5157
rect 13081 5117 13093 5151
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 13630 5108 13636 5160
rect 13688 5148 13694 5160
rect 13725 5151 13783 5157
rect 13725 5148 13737 5151
rect 13688 5120 13737 5148
rect 13688 5108 13694 5120
rect 13725 5117 13737 5120
rect 13771 5117 13783 5151
rect 13725 5111 13783 5117
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14366 5148 14372 5160
rect 14047 5120 14372 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 15948 5157 15976 5256
rect 18322 5244 18328 5256
rect 18380 5284 18386 5296
rect 21269 5287 21327 5293
rect 21269 5284 21281 5287
rect 18380 5256 21281 5284
rect 18380 5244 18386 5256
rect 21269 5253 21281 5256
rect 21315 5284 21327 5287
rect 21542 5284 21548 5296
rect 21315 5256 21548 5284
rect 21315 5253 21327 5256
rect 21269 5247 21327 5253
rect 21542 5244 21548 5256
rect 21600 5244 21606 5296
rect 21821 5287 21879 5293
rect 21821 5253 21833 5287
rect 21867 5253 21879 5287
rect 21821 5247 21879 5253
rect 20993 5219 21051 5225
rect 20993 5185 21005 5219
rect 21039 5216 21051 5219
rect 21450 5216 21456 5228
rect 21039 5188 21456 5216
rect 21039 5185 21051 5188
rect 20993 5179 21051 5185
rect 21450 5176 21456 5188
rect 21508 5216 21514 5228
rect 21836 5216 21864 5247
rect 22002 5244 22008 5296
rect 22060 5244 22066 5296
rect 23106 5244 23112 5296
rect 23164 5284 23170 5296
rect 23477 5287 23535 5293
rect 23477 5284 23489 5287
rect 23164 5256 23489 5284
rect 23164 5244 23170 5256
rect 23477 5253 23489 5256
rect 23523 5253 23535 5287
rect 23477 5247 23535 5253
rect 23658 5244 23664 5296
rect 23716 5244 23722 5296
rect 24121 5287 24179 5293
rect 24121 5253 24133 5287
rect 24167 5284 24179 5287
rect 24670 5284 24676 5296
rect 24167 5256 24676 5284
rect 24167 5253 24179 5256
rect 24121 5247 24179 5253
rect 24670 5244 24676 5256
rect 24728 5284 24734 5296
rect 25133 5287 25191 5293
rect 25133 5284 25145 5287
rect 24728 5256 25145 5284
rect 24728 5244 24734 5256
rect 25133 5253 25145 5256
rect 25179 5253 25191 5287
rect 25133 5247 25191 5253
rect 25317 5287 25375 5293
rect 25317 5253 25329 5287
rect 25363 5284 25375 5287
rect 25363 5256 25820 5284
rect 25363 5253 25375 5256
rect 25317 5247 25375 5253
rect 21508 5188 21864 5216
rect 21508 5176 21514 5188
rect 23198 5176 23204 5228
rect 23256 5216 23262 5228
rect 23293 5219 23351 5225
rect 23293 5216 23305 5219
rect 23256 5188 23305 5216
rect 23256 5176 23262 5188
rect 23293 5185 23305 5188
rect 23339 5185 23351 5219
rect 24210 5216 24216 5228
rect 23293 5179 23351 5185
rect 23768 5188 24216 5216
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18656 5120 18705 5148
rect 18656 5108 18662 5120
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18785 5151 18843 5157
rect 18785 5117 18797 5151
rect 18831 5148 18843 5151
rect 22094 5148 22100 5160
rect 18831 5120 22100 5148
rect 18831 5117 18843 5120
rect 18785 5111 18843 5117
rect 22094 5108 22100 5120
rect 22152 5108 22158 5160
rect 22738 5108 22744 5160
rect 22796 5108 22802 5160
rect 22833 5151 22891 5157
rect 22833 5117 22845 5151
rect 22879 5117 22891 5151
rect 22833 5111 22891 5117
rect 11440 5052 12020 5080
rect 12713 5083 12771 5089
rect 12713 5049 12725 5083
rect 12759 5080 12771 5083
rect 12802 5080 12808 5092
rect 12759 5052 12808 5080
rect 12759 5049 12771 5052
rect 12713 5043 12771 5049
rect 12802 5040 12808 5052
rect 12860 5080 12866 5092
rect 14461 5083 14519 5089
rect 14461 5080 14473 5083
rect 12860 5052 14473 5080
rect 12860 5040 12866 5052
rect 14461 5049 14473 5052
rect 14507 5080 14519 5083
rect 14734 5080 14740 5092
rect 14507 5052 14740 5080
rect 14507 5049 14519 5052
rect 14461 5043 14519 5049
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 21542 5040 21548 5092
rect 21600 5040 21606 5092
rect 21634 5040 21640 5092
rect 21692 5080 21698 5092
rect 22370 5080 22376 5092
rect 21692 5052 22376 5080
rect 21692 5040 21698 5052
rect 22370 5040 22376 5052
rect 22428 5080 22434 5092
rect 22848 5080 22876 5111
rect 22922 5108 22928 5160
rect 22980 5148 22986 5160
rect 23768 5148 23796 5188
rect 24210 5176 24216 5188
rect 24268 5176 24274 5228
rect 24302 5176 24308 5228
rect 24360 5176 24366 5228
rect 24949 5219 25007 5225
rect 24949 5185 24961 5219
rect 24995 5216 25007 5219
rect 25685 5219 25743 5225
rect 25685 5216 25697 5219
rect 24995 5188 25697 5216
rect 24995 5185 25007 5188
rect 24949 5179 25007 5185
rect 25240 5160 25268 5188
rect 25685 5185 25697 5188
rect 25731 5185 25743 5219
rect 25792 5216 25820 5256
rect 25866 5244 25872 5296
rect 25924 5244 25930 5296
rect 28276 5293 28304 5324
rect 28629 5321 28641 5355
rect 28675 5352 28687 5355
rect 29546 5352 29552 5364
rect 28675 5324 29552 5352
rect 28675 5321 28687 5324
rect 28629 5315 28687 5321
rect 29546 5312 29552 5324
rect 29604 5312 29610 5364
rect 28261 5287 28319 5293
rect 28261 5253 28273 5287
rect 28307 5253 28319 5287
rect 28261 5247 28319 5253
rect 28813 5287 28871 5293
rect 28813 5253 28825 5287
rect 28859 5253 28871 5287
rect 28813 5247 28871 5253
rect 26142 5216 26148 5228
rect 25792 5188 26148 5216
rect 25685 5179 25743 5185
rect 26142 5176 26148 5188
rect 26200 5176 26206 5228
rect 22980 5120 23796 5148
rect 22980 5108 22986 5120
rect 23842 5108 23848 5160
rect 23900 5108 23906 5160
rect 23934 5108 23940 5160
rect 23992 5148 23998 5160
rect 24029 5151 24087 5157
rect 24029 5148 24041 5151
rect 23992 5120 24041 5148
rect 23992 5108 23998 5120
rect 24029 5117 24041 5120
rect 24075 5148 24087 5151
rect 24118 5148 24124 5160
rect 24075 5120 24124 5148
rect 24075 5117 24087 5120
rect 24029 5111 24087 5117
rect 24118 5108 24124 5120
rect 24176 5108 24182 5160
rect 25038 5108 25044 5160
rect 25096 5108 25102 5160
rect 25222 5108 25228 5160
rect 25280 5108 25286 5160
rect 27154 5148 27160 5160
rect 25516 5120 27160 5148
rect 22428 5052 22876 5080
rect 23109 5083 23167 5089
rect 22428 5040 22434 5052
rect 23109 5049 23121 5083
rect 23155 5049 23167 5083
rect 23109 5043 23167 5049
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 4981 3111 5015
rect 3053 4975 3111 4981
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3970 5012 3976 5024
rect 3384 4984 3976 5012
rect 3384 4972 3390 4984
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4801 5015 4859 5021
rect 4801 4981 4813 5015
rect 4847 5012 4859 5015
rect 5810 5012 5816 5024
rect 4847 4984 5816 5012
rect 4847 4981 4859 4984
rect 4801 4975 4859 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7892 4984 8033 5012
rect 7892 4972 7898 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 8021 4975 8079 4981
rect 8573 5015 8631 5021
rect 8573 4981 8585 5015
rect 8619 5012 8631 5015
rect 8662 5012 8668 5024
rect 8619 4984 8668 5012
rect 8619 4981 8631 4984
rect 8573 4975 8631 4981
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 8938 4972 8944 5024
rect 8996 4972 9002 5024
rect 10962 4972 10968 5024
rect 11020 5012 11026 5024
rect 11057 5015 11115 5021
rect 11057 5012 11069 5015
rect 11020 4984 11069 5012
rect 11020 4972 11026 4984
rect 11057 4981 11069 4984
rect 11103 4981 11115 5015
rect 11057 4975 11115 4981
rect 11238 4972 11244 5024
rect 11296 4972 11302 5024
rect 11790 4972 11796 5024
rect 11848 4972 11854 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12503 5015 12561 5021
rect 12503 5012 12515 5015
rect 11940 4984 12515 5012
rect 11940 4972 11946 4984
rect 12503 4981 12515 4984
rect 12549 4981 12561 5015
rect 12503 4975 12561 4981
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 5012 12955 5015
rect 12986 5012 12992 5024
rect 12943 4984 12992 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 13541 5015 13599 5021
rect 13541 4981 13553 5015
rect 13587 5012 13599 5015
rect 13814 5012 13820 5024
rect 13587 4984 13820 5012
rect 13587 4981 13599 4984
rect 13541 4975 13599 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14274 5021 14280 5024
rect 14261 5015 14280 5021
rect 14261 4981 14273 5015
rect 14261 4975 14280 4981
rect 14274 4972 14280 4975
rect 14332 4972 14338 5024
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 17310 5012 17316 5024
rect 16347 4984 17316 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 23124 5012 23152 5043
rect 23198 5040 23204 5092
rect 23256 5040 23262 5092
rect 23382 5040 23388 5092
rect 23440 5080 23446 5092
rect 23661 5083 23719 5089
rect 23661 5080 23673 5083
rect 23440 5052 23673 5080
rect 23440 5040 23446 5052
rect 23661 5049 23673 5052
rect 23707 5049 23719 5083
rect 24136 5080 24164 5108
rect 25516 5080 25544 5120
rect 27154 5108 27160 5120
rect 27212 5148 27218 5160
rect 27801 5151 27859 5157
rect 27801 5148 27813 5151
rect 27212 5120 27813 5148
rect 27212 5108 27218 5120
rect 27801 5117 27813 5120
rect 27847 5117 27859 5151
rect 27801 5111 27859 5117
rect 24136 5052 25544 5080
rect 25593 5083 25651 5089
rect 23661 5043 23719 5049
rect 25593 5049 25605 5083
rect 25639 5080 25651 5083
rect 25866 5080 25872 5092
rect 25639 5052 25872 5080
rect 25639 5049 25651 5052
rect 25593 5043 25651 5049
rect 25866 5040 25872 5052
rect 25924 5040 25930 5092
rect 23474 5012 23480 5024
rect 23124 4984 23480 5012
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 23566 4972 23572 5024
rect 23624 5012 23630 5024
rect 24673 5015 24731 5021
rect 24673 5012 24685 5015
rect 23624 4984 24685 5012
rect 23624 4972 23630 4984
rect 24673 4981 24685 4984
rect 24719 4981 24731 5015
rect 27816 5012 27844 5111
rect 27982 5108 27988 5160
rect 28040 5148 28046 5160
rect 28258 5148 28264 5160
rect 28040 5120 28264 5148
rect 28040 5108 28046 5120
rect 28258 5108 28264 5120
rect 28316 5148 28322 5160
rect 28718 5148 28724 5160
rect 28316 5120 28724 5148
rect 28316 5108 28322 5120
rect 28718 5108 28724 5120
rect 28776 5108 28782 5160
rect 28828 5148 28856 5247
rect 28994 5244 29000 5296
rect 29052 5284 29058 5296
rect 29089 5287 29147 5293
rect 29089 5284 29101 5287
rect 29052 5256 29101 5284
rect 29052 5244 29058 5256
rect 29089 5253 29101 5256
rect 29135 5253 29147 5287
rect 29089 5247 29147 5253
rect 30202 5151 30260 5157
rect 30202 5148 30214 5151
rect 28828 5120 30214 5148
rect 30202 5117 30214 5120
rect 30248 5117 30260 5151
rect 30202 5111 30260 5117
rect 30469 5151 30527 5157
rect 30469 5117 30481 5151
rect 30515 5148 30527 5151
rect 30653 5151 30711 5157
rect 30653 5148 30665 5151
rect 30515 5120 30665 5148
rect 30515 5117 30527 5120
rect 30469 5111 30527 5117
rect 30653 5117 30665 5120
rect 30699 5117 30711 5151
rect 30653 5111 30711 5117
rect 30745 5151 30803 5157
rect 30745 5117 30757 5151
rect 30791 5148 30803 5151
rect 30837 5151 30895 5157
rect 30837 5148 30849 5151
rect 30791 5120 30849 5148
rect 30791 5117 30803 5120
rect 30745 5111 30803 5117
rect 30837 5117 30849 5120
rect 30883 5117 30895 5151
rect 30837 5111 30895 5117
rect 28074 5040 28080 5092
rect 28132 5080 28138 5092
rect 28132 5052 30144 5080
rect 28132 5040 28138 5052
rect 28166 5012 28172 5024
rect 27816 4984 28172 5012
rect 24673 4975 24731 4981
rect 28166 4972 28172 4984
rect 28224 4972 28230 5024
rect 28626 4972 28632 5024
rect 28684 4972 28690 5024
rect 30116 5012 30144 5052
rect 30760 5012 30788 5111
rect 30116 4984 30788 5012
rect 30926 4972 30932 5024
rect 30984 4972 30990 5024
rect 552 4922 31648 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 12096 4922
rect 12148 4870 12160 4922
rect 12212 4870 12224 4922
rect 12276 4870 12288 4922
rect 12340 4870 12352 4922
rect 12404 4870 19870 4922
rect 19922 4870 19934 4922
rect 19986 4870 19998 4922
rect 20050 4870 20062 4922
rect 20114 4870 20126 4922
rect 20178 4870 27644 4922
rect 27696 4870 27708 4922
rect 27760 4870 27772 4922
rect 27824 4870 27836 4922
rect 27888 4870 27900 4922
rect 27952 4870 31648 4922
rect 552 4848 31648 4870
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 1946 4808 1952 4820
rect 1903 4780 1952 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 3418 4808 3424 4820
rect 2179 4780 3424 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 3568 4780 3893 4808
rect 3568 4768 3574 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 4028 4780 4077 4808
rect 4028 4768 4034 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 4065 4771 4123 4777
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9490 4808 9496 4820
rect 9263 4780 9496 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 12434 4768 12440 4820
rect 12492 4768 12498 4820
rect 12728 4780 13492 4808
rect 2317 4743 2375 4749
rect 2317 4740 2329 4743
rect 1964 4712 2329 4740
rect 1762 4632 1768 4684
rect 1820 4632 1826 4684
rect 1964 4681 1992 4712
rect 2317 4709 2329 4712
rect 2363 4709 2375 4743
rect 3145 4743 3203 4749
rect 3145 4740 3157 4743
rect 2317 4703 2375 4709
rect 2608 4712 3157 4740
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4641 2007 4675
rect 1949 4635 2007 4641
rect 2038 4632 2044 4684
rect 2096 4632 2102 4684
rect 2608 4681 2636 4712
rect 3145 4709 3157 4712
rect 3191 4709 3203 4743
rect 3145 4703 3203 4709
rect 4246 4700 4252 4752
rect 4304 4740 4310 4752
rect 4677 4743 4735 4749
rect 4677 4740 4689 4743
rect 4304 4712 4689 4740
rect 4304 4700 4310 4712
rect 4677 4709 4689 4712
rect 4723 4709 4735 4743
rect 4677 4703 4735 4709
rect 4890 4700 4896 4752
rect 4948 4700 4954 4752
rect 8104 4743 8162 4749
rect 8104 4709 8116 4743
rect 8150 4740 8162 4743
rect 8938 4740 8944 4752
rect 8150 4712 8944 4740
rect 8150 4709 8162 4712
rect 8104 4703 8162 4709
rect 8938 4700 8944 4712
rect 8996 4700 9002 4752
rect 11238 4749 11244 4752
rect 11232 4740 11244 4749
rect 11199 4712 11244 4740
rect 11232 4703 11244 4712
rect 11238 4700 11244 4703
rect 11296 4700 11302 4752
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 12589 4743 12647 4749
rect 12589 4740 12601 4743
rect 11940 4712 12601 4740
rect 11940 4700 11946 4712
rect 12589 4709 12601 4712
rect 12635 4740 12647 4743
rect 12728 4740 12756 4780
rect 12635 4712 12756 4740
rect 12635 4709 12647 4712
rect 12589 4703 12647 4709
rect 12802 4700 12808 4752
rect 12860 4700 12866 4752
rect 13464 4740 13492 4780
rect 14366 4768 14372 4820
rect 14424 4768 14430 4820
rect 16114 4768 16120 4820
rect 16172 4808 16178 4820
rect 16482 4808 16488 4820
rect 16172 4780 16488 4808
rect 16172 4768 16178 4780
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 18230 4768 18236 4820
rect 18288 4768 18294 4820
rect 18509 4811 18567 4817
rect 18509 4777 18521 4811
rect 18555 4808 18567 4811
rect 18690 4808 18696 4820
rect 18555 4780 18696 4808
rect 18555 4777 18567 4780
rect 18509 4771 18567 4777
rect 18690 4768 18696 4780
rect 18748 4768 18754 4820
rect 19610 4808 19616 4820
rect 18984 4780 19616 4808
rect 14274 4740 14280 4752
rect 13464 4712 14280 4740
rect 14274 4700 14280 4712
rect 14332 4740 14338 4752
rect 14521 4743 14579 4749
rect 14521 4740 14533 4743
rect 14332 4712 14533 4740
rect 14332 4700 14338 4712
rect 14521 4709 14533 4712
rect 14567 4709 14579 4743
rect 14521 4703 14579 4709
rect 14734 4700 14740 4752
rect 14792 4700 14798 4752
rect 17402 4740 17408 4752
rect 14844 4712 17408 4740
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4641 2651 4675
rect 2593 4635 2651 4641
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4641 2927 4675
rect 2869 4635 2927 4641
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4672 3111 4675
rect 3786 4672 3792 4684
rect 3099 4644 3792 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 2314 4564 2320 4616
rect 2372 4564 2378 4616
rect 2501 4539 2559 4545
rect 2501 4505 2513 4539
rect 2547 4536 2559 4539
rect 2884 4536 2912 4635
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 5166 4632 5172 4684
rect 5224 4632 5230 4684
rect 7834 4632 7840 4684
rect 7892 4632 7898 4684
rect 10962 4632 10968 4684
rect 11020 4632 11026 4684
rect 12894 4632 12900 4684
rect 12952 4632 12958 4684
rect 12986 4632 12992 4684
rect 13044 4672 13050 4684
rect 13153 4675 13211 4681
rect 13153 4672 13165 4675
rect 13044 4644 13165 4672
rect 13044 4632 13050 4644
rect 13153 4641 13165 4644
rect 13199 4641 13211 4675
rect 13153 4635 13211 4641
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 13688 4644 14320 4672
rect 13688 4632 13694 4644
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 5534 4604 5540 4616
rect 4479 4576 5540 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 14292 4604 14320 4644
rect 14366 4632 14372 4684
rect 14424 4672 14430 4684
rect 14844 4672 14872 4712
rect 17402 4700 17408 4712
rect 17460 4740 17466 4752
rect 18984 4749 19012 4780
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 22557 4811 22615 4817
rect 22557 4777 22569 4811
rect 22603 4808 22615 4811
rect 22922 4808 22928 4820
rect 22603 4780 22928 4808
rect 22603 4777 22615 4780
rect 22557 4771 22615 4777
rect 22922 4768 22928 4780
rect 22980 4768 22986 4820
rect 23014 4768 23020 4820
rect 23072 4808 23078 4820
rect 23201 4811 23259 4817
rect 23201 4808 23213 4811
rect 23072 4780 23213 4808
rect 23072 4768 23078 4780
rect 23201 4777 23213 4780
rect 23247 4777 23259 4811
rect 23201 4771 23259 4777
rect 23382 4768 23388 4820
rect 23440 4768 23446 4820
rect 27154 4817 27160 4820
rect 24305 4811 24363 4817
rect 24305 4808 24317 4811
rect 23860 4780 24317 4808
rect 18969 4743 19027 4749
rect 17460 4712 17724 4740
rect 17460 4700 17466 4712
rect 14424 4644 14872 4672
rect 14921 4675 14979 4681
rect 14424 4632 14430 4644
rect 14921 4641 14933 4675
rect 14967 4641 14979 4675
rect 14921 4635 14979 4641
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 15470 4672 15476 4684
rect 15151 4644 15476 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 14936 4604 14964 4635
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 16114 4632 16120 4684
rect 16172 4632 16178 4684
rect 16206 4632 16212 4684
rect 16264 4632 16270 4684
rect 16393 4675 16451 4681
rect 16393 4641 16405 4675
rect 16439 4672 16451 4675
rect 16485 4675 16543 4681
rect 16485 4672 16497 4675
rect 16439 4644 16497 4672
rect 16439 4641 16451 4644
rect 16393 4635 16451 4641
rect 16485 4641 16497 4644
rect 16531 4641 16543 4675
rect 16485 4635 16543 4641
rect 14292 4576 14964 4604
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 16408 4604 16436 4635
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 16669 4675 16727 4681
rect 16669 4672 16681 4675
rect 16632 4644 16681 4672
rect 16632 4632 16638 4644
rect 16669 4641 16681 4644
rect 16715 4641 16727 4675
rect 16669 4635 16727 4641
rect 17310 4632 17316 4684
rect 17368 4632 17374 4684
rect 17494 4632 17500 4684
rect 17552 4632 17558 4684
rect 17696 4681 17724 4712
rect 18969 4709 18981 4743
rect 19015 4709 19027 4743
rect 18969 4703 19027 4709
rect 19521 4743 19579 4749
rect 19521 4709 19533 4743
rect 19567 4740 19579 4743
rect 23750 4740 23756 4752
rect 19567 4712 23756 4740
rect 19567 4709 19579 4712
rect 19521 4703 19579 4709
rect 23750 4700 23756 4712
rect 23808 4700 23814 4752
rect 23860 4749 23888 4780
rect 24305 4777 24317 4780
rect 24351 4777 24363 4811
rect 24305 4771 24363 4777
rect 26421 4811 26479 4817
rect 26421 4777 26433 4811
rect 26467 4777 26479 4811
rect 26421 4771 26479 4777
rect 27141 4811 27160 4817
rect 27141 4777 27153 4811
rect 27141 4771 27160 4777
rect 23845 4743 23903 4749
rect 23845 4709 23857 4743
rect 23891 4709 23903 4743
rect 23845 4703 23903 4709
rect 24026 4700 24032 4752
rect 24084 4700 24090 4752
rect 24486 4740 24492 4752
rect 24136 4712 24492 4740
rect 17681 4675 17739 4681
rect 17681 4641 17693 4675
rect 17727 4641 17739 4675
rect 17681 4635 17739 4641
rect 17865 4675 17923 4681
rect 17865 4641 17877 4675
rect 17911 4672 17923 4675
rect 17954 4672 17960 4684
rect 17911 4644 17960 4672
rect 17911 4641 17923 4644
rect 17865 4635 17923 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 18138 4632 18144 4684
rect 18196 4672 18202 4684
rect 19153 4675 19211 4681
rect 19153 4672 19165 4675
rect 18196 4644 19165 4672
rect 18196 4632 18202 4644
rect 19153 4641 19165 4644
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 19246 4675 19304 4681
rect 19246 4641 19258 4675
rect 19292 4641 19304 4675
rect 19246 4635 19304 4641
rect 15068 4576 16436 4604
rect 15068 4564 15074 4576
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 17276 4576 17601 4604
rect 17276 4564 17282 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 18095 4576 18429 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 18506 4564 18512 4616
rect 18564 4604 18570 4616
rect 19260 4604 19288 4635
rect 19426 4632 19432 4684
rect 19484 4632 19490 4684
rect 19659 4675 19717 4681
rect 19659 4641 19671 4675
rect 19705 4672 19717 4675
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 19705 4644 19993 4672
rect 19705 4641 19717 4644
rect 19659 4635 19717 4641
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 19981 4635 20039 4641
rect 20073 4675 20131 4681
rect 20073 4641 20085 4675
rect 20119 4672 20131 4675
rect 20622 4672 20628 4684
rect 20119 4644 20628 4672
rect 20119 4641 20131 4644
rect 20073 4635 20131 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 22646 4632 22652 4684
rect 22704 4632 22710 4684
rect 22830 4632 22836 4684
rect 22888 4632 22894 4684
rect 22925 4675 22983 4681
rect 22925 4641 22937 4675
rect 22971 4641 22983 4675
rect 22925 4635 22983 4641
rect 23017 4675 23075 4681
rect 23017 4641 23029 4675
rect 23063 4672 23075 4675
rect 23290 4672 23296 4684
rect 23063 4644 23296 4672
rect 23063 4641 23075 4644
rect 23017 4635 23075 4641
rect 18564 4576 19288 4604
rect 19352 4576 19840 4604
rect 18564 4564 18570 4576
rect 3602 4536 3608 4548
rect 2547 4508 3608 4536
rect 2547 4505 2559 4508
rect 2501 4499 2559 4505
rect 3602 4496 3608 4508
rect 3660 4536 3666 4548
rect 12345 4539 12403 4545
rect 3660 4508 4568 4536
rect 3660 4496 3666 4508
rect 4540 4480 4568 4508
rect 12345 4505 12357 4539
rect 12391 4536 12403 4539
rect 12526 4536 12532 4548
rect 12391 4508 12532 4536
rect 12391 4505 12403 4508
rect 12345 4499 12403 4505
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 14277 4539 14335 4545
rect 14277 4505 14289 4539
rect 14323 4536 14335 4539
rect 14458 4536 14464 4548
rect 14323 4508 14464 4536
rect 14323 4505 14335 4508
rect 14277 4499 14335 4505
rect 14458 4496 14464 4508
rect 14516 4536 14522 4548
rect 18969 4539 19027 4545
rect 14516 4508 17908 4536
rect 14516 4496 14522 4508
rect 17880 4480 17908 4508
rect 18969 4505 18981 4539
rect 19015 4536 19027 4539
rect 19352 4536 19380 4576
rect 19812 4545 19840 4576
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 22940 4604 22968 4635
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 23569 4675 23627 4681
rect 23569 4641 23581 4675
rect 23615 4641 23627 4675
rect 23569 4635 23627 4641
rect 23474 4604 23480 4616
rect 22940 4576 23480 4604
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 23591 4604 23619 4635
rect 23658 4632 23664 4684
rect 23716 4672 23722 4684
rect 24136 4681 24164 4712
rect 24486 4700 24492 4712
rect 24544 4700 24550 4752
rect 25038 4700 25044 4752
rect 25096 4740 25102 4752
rect 25501 4743 25559 4749
rect 25501 4740 25513 4743
rect 25096 4712 25513 4740
rect 25096 4700 25102 4712
rect 25501 4709 25513 4712
rect 25547 4740 25559 4743
rect 26436 4740 26464 4771
rect 27154 4768 27160 4771
rect 27212 4768 27218 4820
rect 28077 4811 28135 4817
rect 28077 4808 28089 4811
rect 28000 4780 28089 4808
rect 28000 4749 28028 4780
rect 28077 4777 28089 4780
rect 28123 4808 28135 4811
rect 28534 4808 28540 4820
rect 28123 4780 28540 4808
rect 28123 4777 28135 4780
rect 28077 4771 28135 4777
rect 28534 4768 28540 4780
rect 28592 4768 28598 4820
rect 28813 4811 28871 4817
rect 28813 4777 28825 4811
rect 28859 4777 28871 4811
rect 28813 4771 28871 4777
rect 28258 4749 28264 4752
rect 25547 4712 26464 4740
rect 27341 4743 27399 4749
rect 25547 4709 25559 4712
rect 25501 4703 25559 4709
rect 27341 4709 27353 4743
rect 27387 4709 27399 4743
rect 27341 4703 27399 4709
rect 27985 4743 28043 4749
rect 27985 4709 27997 4743
rect 28031 4709 28043 4743
rect 27985 4703 28043 4709
rect 28245 4743 28264 4749
rect 28245 4709 28257 4743
rect 28245 4703 28264 4709
rect 23937 4675 23995 4681
rect 23937 4672 23949 4675
rect 23716 4644 23949 4672
rect 23716 4632 23722 4644
rect 23937 4641 23949 4644
rect 23983 4641 23995 4675
rect 23937 4635 23995 4641
rect 24121 4675 24179 4681
rect 24121 4641 24133 4675
rect 24167 4641 24179 4675
rect 24121 4635 24179 4641
rect 24210 4632 24216 4684
rect 24268 4672 24274 4684
rect 24673 4675 24731 4681
rect 24673 4672 24685 4675
rect 24268 4644 24685 4672
rect 24268 4632 24274 4644
rect 24673 4641 24685 4644
rect 24719 4641 24731 4675
rect 24673 4635 24731 4641
rect 25222 4632 25228 4684
rect 25280 4632 25286 4684
rect 25958 4632 25964 4684
rect 26016 4672 26022 4684
rect 26881 4675 26939 4681
rect 26881 4672 26893 4675
rect 26016 4644 26893 4672
rect 26016 4632 26022 4644
rect 26881 4641 26893 4644
rect 26927 4641 26939 4675
rect 26881 4635 26939 4641
rect 27356 4672 27384 4703
rect 28258 4700 28264 4703
rect 28316 4700 28322 4752
rect 28442 4700 28448 4752
rect 28500 4740 28506 4752
rect 28828 4740 28856 4771
rect 28500 4712 28856 4740
rect 28500 4700 28506 4712
rect 29086 4700 29092 4752
rect 29144 4740 29150 4752
rect 29926 4743 29984 4749
rect 29926 4740 29938 4743
rect 29144 4712 29938 4740
rect 29144 4700 29150 4712
rect 29926 4709 29938 4712
rect 29972 4709 29984 4743
rect 29926 4703 29984 4709
rect 27801 4675 27859 4681
rect 27801 4672 27813 4675
rect 27356 4644 27813 4672
rect 23753 4607 23811 4613
rect 23591 4576 23704 4604
rect 19015 4508 19380 4536
rect 19797 4539 19855 4545
rect 19015 4505 19027 4508
rect 18969 4499 19027 4505
rect 19797 4505 19809 4539
rect 19843 4505 19855 4539
rect 19797 4499 19855 4505
rect 22370 4496 22376 4548
rect 22428 4496 22434 4548
rect 23676 4536 23704 4576
rect 23753 4573 23765 4607
rect 23799 4604 23811 4607
rect 24302 4604 24308 4616
rect 23799 4576 24308 4604
rect 23799 4573 23811 4576
rect 23753 4567 23811 4573
rect 24302 4564 24308 4576
rect 24360 4564 24366 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 24627 4576 25329 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 25317 4573 25329 4576
rect 25363 4604 25375 4607
rect 25593 4607 25651 4613
rect 25593 4604 25605 4607
rect 25363 4576 25605 4604
rect 25363 4573 25375 4576
rect 25317 4567 25375 4573
rect 25593 4573 25605 4576
rect 25639 4573 25651 4607
rect 25593 4567 25651 4573
rect 24026 4536 24032 4548
rect 22480 4508 23612 4536
rect 23676 4508 24032 4536
rect 2682 4428 2688 4480
rect 2740 4428 2746 4480
rect 4062 4428 4068 4480
rect 4120 4428 4126 4480
rect 4522 4428 4528 4480
rect 4580 4428 4586 4480
rect 4706 4428 4712 4480
rect 4764 4428 4770 4480
rect 5074 4428 5080 4480
rect 5132 4428 5138 4480
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 14366 4468 14372 4480
rect 12676 4440 14372 4468
rect 12676 4428 12682 4440
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 14550 4428 14556 4480
rect 14608 4428 14614 4480
rect 14918 4428 14924 4480
rect 14976 4468 14982 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14976 4440 15025 4468
rect 14976 4428 14982 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 16356 4440 16405 4468
rect 16356 4428 16362 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 16393 4431 16451 4437
rect 16669 4471 16727 4477
rect 16669 4437 16681 4471
rect 16715 4468 16727 4471
rect 16942 4468 16948 4480
rect 16715 4440 16948 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 19426 4468 19432 4480
rect 17920 4440 19432 4468
rect 17920 4428 17926 4440
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 22002 4428 22008 4480
rect 22060 4468 22066 4480
rect 22480 4468 22508 4508
rect 23584 4477 23612 4508
rect 24026 4496 24032 4508
rect 24084 4496 24090 4548
rect 24946 4496 24952 4548
rect 25004 4536 25010 4548
rect 25041 4539 25099 4545
rect 25041 4536 25053 4539
rect 25004 4508 25053 4536
rect 25004 4496 25010 4508
rect 25041 4505 25053 4508
rect 25087 4505 25099 4539
rect 25041 4499 25099 4505
rect 25777 4539 25835 4545
rect 25777 4505 25789 4539
rect 25823 4536 25835 4539
rect 25976 4536 26004 4632
rect 26050 4564 26056 4616
rect 26108 4604 26114 4616
rect 26108 4576 26648 4604
rect 26108 4564 26114 4576
rect 26620 4545 26648 4576
rect 25823 4508 26004 4536
rect 26605 4539 26663 4545
rect 25823 4505 25835 4508
rect 25777 4499 25835 4505
rect 26605 4505 26617 4539
rect 26651 4536 26663 4539
rect 27356 4536 27384 4644
rect 27801 4641 27813 4644
rect 27847 4672 27859 4675
rect 28902 4672 28908 4684
rect 27847 4644 28908 4672
rect 27847 4641 27859 4644
rect 27801 4635 27859 4641
rect 28902 4632 28908 4644
rect 28960 4632 28966 4684
rect 30193 4675 30251 4681
rect 30193 4641 30205 4675
rect 30239 4672 30251 4675
rect 30926 4672 30932 4684
rect 30239 4644 30932 4672
rect 30239 4641 30251 4644
rect 30193 4635 30251 4641
rect 30926 4632 30932 4644
rect 30984 4632 30990 4684
rect 28442 4536 28448 4548
rect 26651 4508 27384 4536
rect 27448 4508 28448 4536
rect 26651 4505 26663 4508
rect 26605 4499 26663 4505
rect 22060 4440 22508 4468
rect 23569 4471 23627 4477
rect 22060 4428 22066 4440
rect 23569 4437 23581 4471
rect 23615 4437 23627 4471
rect 23569 4431 23627 4437
rect 24670 4428 24676 4480
rect 24728 4428 24734 4480
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 25225 4471 25283 4477
rect 25225 4468 25237 4471
rect 24820 4440 25237 4468
rect 24820 4428 24826 4440
rect 25225 4437 25237 4440
rect 25271 4437 25283 4471
rect 25225 4431 25283 4437
rect 26878 4428 26884 4480
rect 26936 4468 26942 4480
rect 26973 4471 27031 4477
rect 26973 4468 26985 4471
rect 26936 4440 26985 4468
rect 26936 4428 26942 4440
rect 26973 4437 26985 4440
rect 27019 4437 27031 4471
rect 26973 4431 27031 4437
rect 27157 4471 27215 4477
rect 27157 4437 27169 4471
rect 27203 4468 27215 4471
rect 27448 4468 27476 4508
rect 28442 4496 28448 4508
rect 28500 4496 28506 4548
rect 27203 4440 27476 4468
rect 27203 4437 27215 4440
rect 27157 4431 27215 4437
rect 27614 4428 27620 4480
rect 27672 4428 27678 4480
rect 28166 4428 28172 4480
rect 28224 4468 28230 4480
rect 28261 4471 28319 4477
rect 28261 4468 28273 4471
rect 28224 4440 28273 4468
rect 28224 4428 28230 4440
rect 28261 4437 28273 4440
rect 28307 4468 28319 4471
rect 28994 4468 29000 4480
rect 28307 4440 29000 4468
rect 28307 4437 28319 4440
rect 28261 4431 28319 4437
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 552 4378 31648 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 11436 4378
rect 11488 4326 11500 4378
rect 11552 4326 11564 4378
rect 11616 4326 11628 4378
rect 11680 4326 11692 4378
rect 11744 4326 19210 4378
rect 19262 4326 19274 4378
rect 19326 4326 19338 4378
rect 19390 4326 19402 4378
rect 19454 4326 19466 4378
rect 19518 4326 26984 4378
rect 27036 4326 27048 4378
rect 27100 4326 27112 4378
rect 27164 4326 27176 4378
rect 27228 4326 27240 4378
rect 27292 4326 31648 4378
rect 552 4304 31648 4326
rect 2424 4236 3004 4264
rect 2038 4020 2044 4072
rect 2096 4020 2102 4072
rect 2424 4069 2452 4236
rect 2682 4156 2688 4208
rect 2740 4156 2746 4208
rect 2976 4205 3004 4236
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 4157 4267 4215 4273
rect 4157 4264 4169 4267
rect 4120 4236 4169 4264
rect 4120 4224 4126 4236
rect 4157 4233 4169 4236
rect 4203 4233 4215 4267
rect 4157 4227 4215 4233
rect 7576 4236 8432 4264
rect 2961 4199 3019 4205
rect 2961 4165 2973 4199
rect 3007 4196 3019 4199
rect 3418 4196 3424 4208
rect 3007 4168 3424 4196
rect 3007 4165 3019 4168
rect 2961 4159 3019 4165
rect 3418 4156 3424 4168
rect 3476 4196 3482 4208
rect 4246 4196 4252 4208
rect 3476 4168 4252 4196
rect 3476 4156 3482 4168
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 4522 4156 4528 4208
rect 4580 4156 4586 4208
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 4764 4168 5764 4196
rect 4764 4156 4770 4168
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2777 4131 2835 4137
rect 2777 4128 2789 4131
rect 2556 4100 2789 4128
rect 2556 4088 2562 4100
rect 2777 4097 2789 4100
rect 2823 4128 2835 4131
rect 4062 4128 4068 4140
rect 2823 4100 4068 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5534 4128 5540 4140
rect 5215 4100 5540 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 5736 4128 5764 4168
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5736 4100 5917 4128
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 7576 4128 7604 4236
rect 7837 4199 7895 4205
rect 7837 4165 7849 4199
rect 7883 4196 7895 4199
rect 8404 4196 8432 4236
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8904 4236 9045 4264
rect 8904 4224 8910 4236
rect 9033 4233 9045 4236
rect 9079 4233 9091 4267
rect 9033 4227 9091 4233
rect 14550 4224 14556 4276
rect 14608 4264 14614 4276
rect 14921 4267 14979 4273
rect 14921 4264 14933 4267
rect 14608 4236 14933 4264
rect 14608 4224 14614 4236
rect 14921 4233 14933 4236
rect 14967 4233 14979 4267
rect 14921 4227 14979 4233
rect 16206 4224 16212 4276
rect 16264 4264 16270 4276
rect 16264 4236 16712 4264
rect 16264 4224 16270 4236
rect 9122 4196 9128 4208
rect 7883 4168 8340 4196
rect 8404 4168 9128 4196
rect 7883 4165 7895 4168
rect 7837 4159 7895 4165
rect 6236 4100 7604 4128
rect 6236 4088 6242 4100
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2363 4032 2421 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2866 4060 2872 4072
rect 2409 4023 2467 4029
rect 2516 4032 2872 4060
rect 2148 3992 2176 4023
rect 2516 3992 2544 4032
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4060 3111 4063
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 3099 4032 3249 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 3237 4029 3249 4032
rect 3283 4029 3295 4063
rect 3237 4023 3295 4029
rect 2148 3964 2544 3992
rect 2685 3995 2743 4001
rect 2685 3961 2697 3995
rect 2731 3992 2743 3995
rect 2777 3995 2835 4001
rect 2777 3992 2789 3995
rect 2731 3964 2789 3992
rect 2731 3961 2743 3964
rect 2685 3955 2743 3961
rect 2777 3961 2789 3964
rect 2823 3961 2835 3995
rect 2777 3955 2835 3961
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 1820 3896 1961 3924
rect 1820 3884 1826 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 1949 3887 2007 3893
rect 2222 3884 2228 3936
rect 2280 3884 2286 3936
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 3068 3924 3096 4023
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 3384 4032 3893 4060
rect 3384 4020 3390 4032
rect 3881 4029 3893 4032
rect 3927 4060 3939 4063
rect 4890 4060 4896 4072
rect 3927 4032 4896 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 4982 4020 4988 4072
rect 5040 4020 5046 4072
rect 5994 4020 6000 4072
rect 6052 4069 6058 4072
rect 6052 4063 6080 4069
rect 6068 4029 6080 4063
rect 6052 4023 6080 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 8051 4063 8109 4069
rect 8051 4060 8063 4063
rect 6871 4032 8063 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 8051 4029 8063 4032
rect 8097 4029 8109 4063
rect 8051 4023 8109 4029
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4029 8263 4063
rect 8312 4060 8340 4168
rect 9122 4156 9128 4168
rect 9180 4156 9186 4208
rect 16684 4205 16712 4236
rect 18138 4224 18144 4276
rect 18196 4224 18202 4276
rect 18325 4267 18383 4273
rect 18325 4233 18337 4267
rect 18371 4264 18383 4267
rect 19337 4267 19395 4273
rect 18371 4236 18736 4264
rect 18371 4233 18383 4236
rect 18325 4227 18383 4233
rect 16669 4199 16727 4205
rect 16669 4165 16681 4199
rect 16715 4196 16727 4199
rect 18598 4196 18604 4208
rect 16715 4168 18604 4196
rect 16715 4165 16727 4168
rect 16669 4159 16727 4165
rect 9490 4128 9496 4140
rect 9048 4100 9496 4128
rect 8603 4063 8661 4069
rect 8603 4060 8615 4063
rect 8312 4032 8615 4060
rect 8205 4023 8263 4029
rect 8603 4029 8615 4032
rect 8649 4029 8661 4063
rect 8603 4023 8661 4029
rect 6052 4020 6058 4023
rect 8220 3992 8248 4023
rect 9048 3992 9076 4100
rect 9490 4088 9496 4100
rect 9548 4128 9554 4140
rect 17328 4137 17356 4168
rect 18598 4156 18604 4168
rect 18656 4156 18662 4208
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9548 4100 9781 4128
rect 9548 4088 9554 4100
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4128 10379 4131
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10367 4100 10517 4128
rect 10367 4097 10379 4100
rect 10321 4091 10379 4097
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17460 4100 17509 4128
rect 17460 4088 17466 4100
rect 17497 4097 17509 4100
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 17957 4131 18015 4137
rect 17957 4097 17969 4131
rect 18003 4128 18015 4131
rect 18506 4128 18512 4140
rect 18003 4100 18512 4128
rect 18003 4097 18015 4100
rect 17957 4091 18015 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18708 4128 18736 4236
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19610 4264 19616 4276
rect 19383 4236 19616 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19610 4224 19616 4236
rect 19668 4224 19674 4276
rect 23474 4224 23480 4276
rect 23532 4264 23538 4276
rect 23937 4267 23995 4273
rect 23937 4264 23949 4267
rect 23532 4236 23949 4264
rect 23532 4224 23538 4236
rect 23937 4233 23949 4236
rect 23983 4264 23995 4267
rect 24486 4264 24492 4276
rect 23983 4236 24492 4264
rect 23983 4233 23995 4236
rect 23937 4227 23995 4233
rect 24486 4224 24492 4236
rect 24544 4224 24550 4276
rect 27614 4224 27620 4276
rect 27672 4264 27678 4276
rect 28629 4267 28687 4273
rect 28629 4264 28641 4267
rect 27672 4236 28641 4264
rect 27672 4224 27678 4236
rect 28629 4233 28641 4236
rect 28675 4233 28687 4267
rect 28629 4227 28687 4233
rect 22186 4156 22192 4208
rect 22244 4196 22250 4208
rect 23201 4199 23259 4205
rect 23201 4196 23213 4199
rect 22244 4168 23213 4196
rect 22244 4156 22250 4168
rect 23201 4165 23213 4168
rect 23247 4165 23259 4199
rect 23201 4159 23259 4165
rect 18708 4100 18828 4128
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 9171 4032 9260 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 8220 3964 9076 3992
rect 2547 3896 3096 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 3970 3884 3976 3936
rect 4028 3884 4034 3936
rect 4154 3884 4160 3936
rect 4212 3884 4218 3936
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 5994 3924 6000 3936
rect 4948 3896 6000 3924
rect 4948 3884 4954 3896
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 8478 3884 8484 3936
rect 8536 3884 8542 3936
rect 8662 3884 8668 3936
rect 8720 3884 8726 3936
rect 9232 3933 9260 4032
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9640 4032 9689 4060
rect 9640 4020 9646 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4060 10471 4063
rect 11146 4060 11152 4072
rect 10459 4032 11152 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 11146 4020 11152 4032
rect 11204 4060 11210 4072
rect 13170 4060 13176 4072
rect 11204 4032 13176 4060
rect 11204 4020 11210 4032
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13814 4069 13820 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13311 4032 13553 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13808 4060 13820 4069
rect 13775 4032 13820 4060
rect 13541 4023 13599 4029
rect 13808 4023 13820 4032
rect 13814 4020 13820 4023
rect 13872 4020 13878 4072
rect 15010 4020 15016 4072
rect 15068 4020 15074 4072
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 15289 4063 15347 4069
rect 15289 4060 15301 4063
rect 15151 4032 15301 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 15289 4029 15301 4032
rect 15335 4029 15347 4063
rect 15289 4023 15347 4029
rect 17862 4020 17868 4072
rect 17920 4060 17926 4072
rect 17920 4032 17964 4060
rect 17920 4020 17926 4032
rect 18230 4020 18236 4072
rect 18288 4020 18294 4072
rect 18414 4020 18420 4072
rect 18472 4020 18478 4072
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 18800 4069 18828 4100
rect 18966 4088 18972 4140
rect 19024 4088 19030 4140
rect 22738 4128 22744 4140
rect 21836 4100 22744 4128
rect 18693 4063 18751 4069
rect 18693 4060 18705 4063
rect 18656 4032 18705 4060
rect 18656 4020 18662 4032
rect 18693 4029 18705 4032
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 18786 4063 18844 4069
rect 18786 4029 18798 4063
rect 18832 4029 18844 4063
rect 18984 4060 19012 4088
rect 19158 4063 19216 4069
rect 19158 4060 19170 4063
rect 18984 4032 19170 4060
rect 18786 4023 18844 4029
rect 19158 4029 19170 4032
rect 19204 4029 19216 4063
rect 19158 4023 19216 4029
rect 10772 3995 10830 4001
rect 10772 3961 10784 3995
rect 10818 3992 10830 3995
rect 11790 3992 11796 4004
rect 10818 3964 11796 3992
rect 10818 3961 10830 3964
rect 10772 3955 10830 3961
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 15556 3995 15614 4001
rect 15556 3961 15568 3995
rect 15602 3992 15614 3995
rect 16114 3992 16120 4004
rect 15602 3964 16120 3992
rect 15602 3961 15614 3964
rect 15556 3955 15614 3961
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 17589 3995 17647 4001
rect 17589 3961 17601 3995
rect 17635 3961 17647 3995
rect 17589 3955 17647 3961
rect 9217 3927 9275 3933
rect 9217 3893 9229 3927
rect 9263 3893 9275 3927
rect 9217 3887 9275 3893
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9364 3896 9597 3924
rect 9364 3884 9370 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9585 3887 9643 3893
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 12618 3924 12624 3936
rect 11931 3896 12624 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 16758 3884 16764 3936
rect 16816 3884 16822 3936
rect 17604 3924 17632 3955
rect 18966 3952 18972 4004
rect 19024 3952 19030 4004
rect 19058 3952 19064 4004
rect 19116 3952 19122 4004
rect 17954 3924 17960 3936
rect 17604 3896 17960 3924
rect 17954 3884 17960 3896
rect 18012 3924 18018 3936
rect 21836 3933 21864 4100
rect 22738 4088 22744 4100
rect 22796 4088 22802 4140
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 22925 4131 22983 4137
rect 22925 4128 22937 4131
rect 22888 4100 22937 4128
rect 22888 4088 22894 4100
rect 22925 4097 22937 4100
rect 22971 4097 22983 4131
rect 22925 4091 22983 4097
rect 23385 4131 23443 4137
rect 23385 4097 23397 4131
rect 23431 4128 23443 4131
rect 24762 4128 24768 4140
rect 23431 4100 24768 4128
rect 23431 4097 23443 4100
rect 23385 4091 23443 4097
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 26878 4088 26884 4140
rect 26936 4128 26942 4140
rect 26936 4100 27476 4128
rect 26936 4088 26942 4100
rect 21913 4063 21971 4069
rect 21913 4029 21925 4063
rect 21959 4060 21971 4063
rect 22094 4060 22100 4072
rect 21959 4032 22100 4060
rect 21959 4029 21971 4032
rect 21913 4023 21971 4029
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 23750 4020 23756 4072
rect 23808 4060 23814 4072
rect 24029 4063 24087 4069
rect 24029 4060 24041 4063
rect 23808 4032 24041 4060
rect 23808 4020 23814 4032
rect 24029 4029 24041 4032
rect 24075 4060 24087 4063
rect 25222 4060 25228 4072
rect 24075 4032 25228 4060
rect 24075 4029 24087 4032
rect 24029 4023 24087 4029
rect 25222 4020 25228 4032
rect 25280 4020 25286 4072
rect 27246 4020 27252 4072
rect 27304 4020 27310 4072
rect 27448 4069 27476 4100
rect 27433 4063 27491 4069
rect 27433 4029 27445 4063
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 27617 4063 27675 4069
rect 27617 4029 27629 4063
rect 27663 4060 27675 4063
rect 27982 4060 27988 4072
rect 27663 4032 27988 4060
rect 27663 4029 27675 4032
rect 27617 4023 27675 4029
rect 27982 4020 27988 4032
rect 28040 4060 28046 4072
rect 28261 4063 28319 4069
rect 28261 4060 28273 4063
rect 28040 4032 28273 4060
rect 28040 4020 28046 4032
rect 28261 4029 28273 4032
rect 28307 4029 28319 4063
rect 28261 4023 28319 4029
rect 28994 4020 29000 4072
rect 29052 4020 29058 4072
rect 27264 3992 27292 4020
rect 27890 3992 27896 4004
rect 27264 3964 27896 3992
rect 27890 3952 27896 3964
rect 27948 3952 27954 4004
rect 28626 3952 28632 4004
rect 28684 3952 28690 4004
rect 29242 3995 29300 4001
rect 29242 3992 29254 3995
rect 28828 3964 29254 3992
rect 28828 3933 28856 3964
rect 29242 3961 29254 3964
rect 29288 3961 29300 3995
rect 29242 3955 29300 3961
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 18012 3896 21833 3924
rect 18012 3884 18018 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 28813 3927 28871 3933
rect 28813 3893 28825 3927
rect 28859 3893 28871 3927
rect 28813 3887 28871 3893
rect 28902 3884 28908 3936
rect 28960 3924 28966 3936
rect 30377 3927 30435 3933
rect 30377 3924 30389 3927
rect 28960 3896 30389 3924
rect 28960 3884 28966 3896
rect 30377 3893 30389 3896
rect 30423 3893 30435 3927
rect 30377 3887 30435 3893
rect 552 3834 31648 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 12096 3834
rect 12148 3782 12160 3834
rect 12212 3782 12224 3834
rect 12276 3782 12288 3834
rect 12340 3782 12352 3834
rect 12404 3782 19870 3834
rect 19922 3782 19934 3834
rect 19986 3782 19998 3834
rect 20050 3782 20062 3834
rect 20114 3782 20126 3834
rect 20178 3782 27644 3834
rect 27696 3782 27708 3834
rect 27760 3782 27772 3834
rect 27824 3782 27836 3834
rect 27888 3782 27900 3834
rect 27952 3782 31648 3834
rect 552 3760 31648 3782
rect 3145 3723 3203 3729
rect 3145 3689 3157 3723
rect 3191 3720 3203 3723
rect 3326 3720 3332 3732
rect 3191 3692 3332 3720
rect 3191 3689 3203 3692
rect 3145 3683 3203 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 3418 3680 3424 3732
rect 3476 3680 3482 3732
rect 16114 3680 16120 3732
rect 16172 3680 16178 3732
rect 18230 3720 18236 3732
rect 17972 3692 18236 3720
rect 2032 3655 2090 3661
rect 2032 3621 2044 3655
rect 2078 3652 2090 3655
rect 2682 3652 2688 3664
rect 2078 3624 2688 3652
rect 2078 3621 2090 3624
rect 2032 3615 2090 3621
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 5074 3652 5080 3664
rect 4080 3624 5080 3652
rect 1762 3544 1768 3596
rect 1820 3544 1826 3596
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 4080 3593 4108 3624
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 9953 3655 10011 3661
rect 9953 3621 9965 3655
rect 9999 3652 10011 3655
rect 10962 3652 10968 3664
rect 9999 3624 10968 3652
rect 9999 3621 10011 3624
rect 9953 3615 10011 3621
rect 10962 3612 10968 3624
rect 11020 3612 11026 3664
rect 17126 3652 17132 3664
rect 14108 3624 17132 3652
rect 3605 3587 3663 3593
rect 3605 3584 3617 3587
rect 3476 3556 3617 3584
rect 3476 3544 3482 3556
rect 3605 3553 3617 3556
rect 3651 3553 3663 3587
rect 3605 3547 3663 3553
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 4321 3587 4379 3593
rect 4321 3584 4333 3587
rect 4065 3547 4123 3553
rect 4172 3556 4333 3584
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 3835 3488 3924 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 3896 3380 3924 3488
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 4172 3516 4200 3556
rect 4321 3553 4333 3556
rect 4367 3553 4379 3587
rect 4321 3547 4379 3553
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 14108 3593 14136 3624
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 17972 3661 18000 3692
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 18966 3720 18972 3732
rect 18371 3692 18972 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 21542 3680 21548 3732
rect 21600 3720 21606 3732
rect 21821 3723 21879 3729
rect 21821 3720 21833 3723
rect 21600 3692 21833 3720
rect 21600 3680 21606 3692
rect 21821 3689 21833 3692
rect 21867 3720 21879 3723
rect 22370 3720 22376 3732
rect 21867 3692 22376 3720
rect 21867 3689 21879 3692
rect 21821 3683 21879 3689
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 22646 3720 22652 3732
rect 22480 3692 22652 3720
rect 17957 3655 18015 3661
rect 17957 3621 17969 3655
rect 18003 3621 18015 3655
rect 17957 3615 18015 3621
rect 18141 3655 18199 3661
rect 18141 3621 18153 3655
rect 18187 3652 18199 3655
rect 18414 3652 18420 3664
rect 18187 3624 18420 3652
rect 18187 3621 18199 3624
rect 18141 3615 18199 3621
rect 18414 3612 18420 3624
rect 18472 3652 18478 3664
rect 18472 3624 21956 3652
rect 18472 3612 18478 3624
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 8536 3556 14105 3584
rect 8536 3544 8542 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 14277 3587 14335 3593
rect 14277 3553 14289 3587
rect 14323 3584 14335 3587
rect 14918 3584 14924 3596
rect 14323 3556 14924 3584
rect 14323 3553 14335 3556
rect 14277 3547 14335 3553
rect 14918 3544 14924 3556
rect 14976 3544 14982 3596
rect 16298 3544 16304 3596
rect 16356 3544 16362 3596
rect 16482 3544 16488 3596
rect 16540 3544 16546 3596
rect 16577 3587 16635 3593
rect 16577 3553 16589 3587
rect 16623 3584 16635 3587
rect 16758 3584 16764 3596
rect 16623 3556 16764 3584
rect 16623 3553 16635 3556
rect 16577 3547 16635 3553
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 4028 3488 4200 3516
rect 4028 3476 4034 3488
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 7926 3516 7932 3528
rect 5684 3488 7932 3516
rect 5684 3476 5690 3488
rect 7926 3476 7932 3488
rect 7984 3516 7990 3528
rect 8754 3516 8760 3528
rect 7984 3488 8760 3516
rect 7984 3476 7990 3488
rect 8754 3476 8760 3488
rect 8812 3516 8818 3528
rect 10502 3516 10508 3528
rect 8812 3488 10508 3516
rect 8812 3476 8818 3488
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 17144 3516 17172 3612
rect 18506 3544 18512 3596
rect 18564 3544 18570 3596
rect 18601 3587 18659 3593
rect 18601 3553 18613 3587
rect 18647 3584 18659 3587
rect 18874 3584 18880 3596
rect 18647 3556 18880 3584
rect 18647 3553 18659 3556
rect 18601 3547 18659 3553
rect 18874 3544 18880 3556
rect 18932 3584 18938 3596
rect 21928 3593 21956 3624
rect 22094 3612 22100 3664
rect 22152 3612 22158 3664
rect 21729 3587 21787 3593
rect 18932 3556 21680 3584
rect 18932 3544 18938 3556
rect 21542 3516 21548 3528
rect 17144 3488 21548 3516
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 8938 3408 8944 3460
rect 8996 3448 9002 3460
rect 9585 3451 9643 3457
rect 9585 3448 9597 3451
rect 8996 3420 9597 3448
rect 8996 3408 9002 3420
rect 9585 3417 9597 3420
rect 9631 3417 9643 3451
rect 11790 3448 11796 3460
rect 9585 3411 9643 3417
rect 9968 3420 11796 3448
rect 4982 3380 4988 3392
rect 3896 3352 4988 3380
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 5442 3340 5448 3392
rect 5500 3340 5506 3392
rect 8478 3340 8484 3392
rect 8536 3380 8542 3392
rect 9968 3389 9996 3420
rect 11790 3408 11796 3420
rect 11848 3408 11854 3460
rect 9953 3383 10011 3389
rect 9953 3380 9965 3383
rect 8536 3352 9965 3380
rect 8536 3340 8542 3352
rect 9953 3349 9965 3352
rect 9999 3349 10011 3383
rect 9953 3343 10011 3349
rect 10137 3383 10195 3389
rect 10137 3349 10149 3383
rect 10183 3380 10195 3383
rect 11054 3380 11060 3392
rect 10183 3352 11060 3380
rect 10183 3349 10195 3352
rect 10137 3343 10195 3349
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 14277 3383 14335 3389
rect 14277 3349 14289 3383
rect 14323 3380 14335 3383
rect 14366 3380 14372 3392
rect 14323 3352 14372 3380
rect 14323 3349 14335 3352
rect 14277 3343 14335 3349
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 20898 3340 20904 3392
rect 20956 3380 20962 3392
rect 21545 3383 21603 3389
rect 21545 3380 21557 3383
rect 20956 3352 21557 3380
rect 20956 3340 20962 3352
rect 21545 3349 21557 3352
rect 21591 3349 21603 3383
rect 21652 3380 21680 3556
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 21913 3587 21971 3593
rect 21913 3553 21925 3587
rect 21959 3584 21971 3587
rect 22186 3584 22192 3596
rect 21959 3556 22192 3584
rect 21959 3553 21971 3556
rect 21913 3547 21971 3553
rect 21744 3516 21772 3547
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 22480 3593 22508 3692
rect 22646 3680 22652 3692
rect 22704 3720 22710 3732
rect 24670 3720 24676 3732
rect 22704 3692 24676 3720
rect 22704 3680 22710 3692
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 25130 3680 25136 3732
rect 25188 3680 25194 3732
rect 25222 3680 25228 3732
rect 25280 3680 25286 3732
rect 25317 3723 25375 3729
rect 25317 3689 25329 3723
rect 25363 3720 25375 3723
rect 25363 3692 27016 3720
rect 25363 3689 25375 3692
rect 25317 3683 25375 3689
rect 25593 3655 25651 3661
rect 25593 3652 25605 3655
rect 22572 3624 25605 3652
rect 22281 3587 22339 3593
rect 22281 3553 22293 3587
rect 22327 3584 22339 3587
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22327 3556 22477 3584
rect 22327 3553 22339 3556
rect 22281 3547 22339 3553
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 22465 3547 22523 3553
rect 22572 3516 22600 3624
rect 22756 3593 22784 3624
rect 25593 3621 25605 3624
rect 25639 3621 25651 3655
rect 25593 3615 25651 3621
rect 25869 3655 25927 3661
rect 25869 3621 25881 3655
rect 25915 3652 25927 3655
rect 26757 3655 26815 3661
rect 26757 3652 26769 3655
rect 25915 3624 26769 3652
rect 25915 3621 25927 3624
rect 25869 3615 25927 3621
rect 26757 3621 26769 3624
rect 26803 3652 26815 3655
rect 26878 3652 26884 3664
rect 26803 3624 26884 3652
rect 26803 3621 26815 3624
rect 26757 3615 26815 3621
rect 26878 3612 26884 3624
rect 26936 3612 26942 3664
rect 26988 3661 27016 3692
rect 28994 3680 29000 3732
rect 29052 3720 29058 3732
rect 29181 3723 29239 3729
rect 29181 3720 29193 3723
rect 29052 3692 29193 3720
rect 29052 3680 29058 3692
rect 29181 3689 29193 3692
rect 29227 3689 29239 3723
rect 29181 3683 29239 3689
rect 26973 3655 27031 3661
rect 26973 3621 26985 3655
rect 27019 3621 27031 3655
rect 26973 3615 27031 3621
rect 22649 3587 22707 3593
rect 22649 3553 22661 3587
rect 22695 3553 22707 3587
rect 22649 3547 22707 3553
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3553 22799 3587
rect 22741 3547 22799 3553
rect 21744 3488 22600 3516
rect 22664 3516 22692 3547
rect 22830 3544 22836 3596
rect 22888 3584 22894 3596
rect 22925 3587 22983 3593
rect 22925 3584 22937 3587
rect 22888 3556 22937 3584
rect 22888 3544 22894 3556
rect 22925 3553 22937 3556
rect 22971 3553 22983 3587
rect 22925 3547 22983 3553
rect 25501 3587 25559 3593
rect 25501 3553 25513 3587
rect 25547 3584 25559 3587
rect 25777 3587 25835 3593
rect 25777 3584 25789 3587
rect 25547 3556 25789 3584
rect 25547 3553 25559 3556
rect 25501 3547 25559 3553
rect 25777 3553 25789 3556
rect 25823 3553 25835 3587
rect 25777 3547 25835 3553
rect 25961 3587 26019 3593
rect 25961 3553 25973 3587
rect 26007 3553 26019 3587
rect 25961 3547 26019 3553
rect 22664 3488 22876 3516
rect 22370 3448 22376 3460
rect 22204 3420 22376 3448
rect 22204 3380 22232 3420
rect 22370 3408 22376 3420
rect 22428 3408 22434 3460
rect 22848 3392 22876 3488
rect 21652 3352 22232 3380
rect 21545 3343 21603 3349
rect 22646 3340 22652 3392
rect 22704 3340 22710 3392
rect 22830 3340 22836 3392
rect 22888 3340 22894 3392
rect 22940 3380 22968 3547
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 25976 3516 26004 3547
rect 26142 3544 26148 3596
rect 26200 3544 26206 3596
rect 26988 3584 27016 3615
rect 27982 3612 27988 3664
rect 28040 3612 28046 3664
rect 28169 3655 28227 3661
rect 28169 3621 28181 3655
rect 28215 3652 28227 3655
rect 30374 3652 30380 3664
rect 28215 3624 30380 3652
rect 28215 3621 28227 3624
rect 28169 3615 28227 3621
rect 28184 3584 28212 3615
rect 30374 3612 30380 3624
rect 30432 3612 30438 3664
rect 26988 3556 28212 3584
rect 29273 3587 29331 3593
rect 29273 3553 29285 3587
rect 29319 3553 29331 3587
rect 29273 3547 29331 3553
rect 26510 3516 26516 3528
rect 24636 3488 26516 3516
rect 24636 3476 24642 3488
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 28074 3476 28080 3528
rect 28132 3516 28138 3528
rect 29288 3516 29316 3547
rect 28132 3488 29316 3516
rect 28132 3476 28138 3488
rect 24946 3408 24952 3460
rect 25004 3408 25010 3460
rect 27246 3448 27252 3460
rect 26528 3420 27252 3448
rect 26528 3380 26556 3420
rect 22940 3352 26556 3380
rect 26602 3340 26608 3392
rect 26660 3340 26666 3392
rect 26804 3389 26832 3420
rect 27246 3408 27252 3420
rect 27304 3408 27310 3460
rect 26789 3383 26847 3389
rect 26789 3349 26801 3383
rect 26835 3349 26847 3383
rect 26789 3343 26847 3349
rect 28350 3340 28356 3392
rect 28408 3340 28414 3392
rect 552 3290 31648 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 11436 3290
rect 11488 3238 11500 3290
rect 11552 3238 11564 3290
rect 11616 3238 11628 3290
rect 11680 3238 11692 3290
rect 11744 3238 19210 3290
rect 19262 3238 19274 3290
rect 19326 3238 19338 3290
rect 19390 3238 19402 3290
rect 19454 3238 19466 3290
rect 19518 3238 26984 3290
rect 27036 3238 27048 3290
rect 27100 3238 27112 3290
rect 27164 3238 27176 3290
rect 27228 3238 27240 3290
rect 27292 3238 31648 3290
rect 552 3216 31648 3238
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 4154 3176 4160 3188
rect 4111 3148 4160 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 5592 3148 6009 3176
rect 5592 3136 5598 3148
rect 5997 3145 6009 3148
rect 6043 3176 6055 3179
rect 6362 3176 6368 3188
rect 6043 3148 6368 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 9306 3136 9312 3188
rect 9364 3136 9370 3188
rect 10410 3176 10416 3188
rect 9508 3148 10416 3176
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 4982 3108 4988 3120
rect 3099 3080 4988 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1489 2975 1547 2981
rect 1489 2941 1501 2975
rect 1535 2972 1547 2975
rect 1673 2975 1731 2981
rect 1673 2972 1685 2975
rect 1535 2944 1685 2972
rect 1535 2941 1547 2944
rect 1489 2935 1547 2941
rect 1673 2941 1685 2944
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 1940 2975 1998 2981
rect 1940 2941 1952 2975
rect 1986 2972 1998 2975
rect 2222 2972 2228 2984
rect 1986 2944 2228 2972
rect 1986 2941 1998 2944
rect 1940 2935 1998 2941
rect 1412 2904 1440 2935
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 3988 2981 4016 3080
rect 4448 3049 4476 3080
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 7101 3111 7159 3117
rect 7101 3108 7113 3111
rect 6236 3080 7113 3108
rect 6236 3068 6242 3080
rect 7101 3077 7113 3080
rect 7147 3077 7159 3111
rect 7101 3071 7159 3077
rect 9214 3068 9220 3120
rect 9272 3068 9278 3120
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4706 3040 4712 3052
rect 4571 3012 4712 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 2038 2904 2044 2916
rect 1412 2876 2044 2904
rect 2038 2864 2044 2876
rect 2096 2864 2102 2916
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 4264 2904 4292 3003
rect 4706 3000 4712 3012
rect 4764 3040 4770 3052
rect 5442 3040 5448 3052
rect 4764 3012 5448 3040
rect 4764 3000 4770 3012
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3040 6331 3043
rect 8110 3040 8116 3052
rect 6319 3012 7144 3040
rect 6319 3009 6331 3012
rect 6273 3003 6331 3009
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2972 4399 2975
rect 4890 2972 4896 2984
rect 4387 2944 4896 2972
rect 4387 2941 4399 2944
rect 4341 2935 4399 2941
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5399 2944 6316 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5184 2904 5212 2935
rect 3476 2876 5856 2904
rect 3476 2864 3482 2876
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 3510 2836 3516 2848
rect 3375 2808 3516 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5828 2845 5856 2876
rect 6086 2864 6092 2916
rect 6144 2904 6150 2916
rect 6288 2913 6316 2944
rect 6454 2932 6460 2984
rect 6512 2932 6518 2984
rect 6549 2975 6607 2981
rect 6549 2941 6561 2975
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 6181 2907 6239 2913
rect 6181 2904 6193 2907
rect 6144 2876 6193 2904
rect 6144 2864 6150 2876
rect 6181 2873 6193 2876
rect 6227 2873 6239 2907
rect 6181 2867 6239 2873
rect 6273 2907 6331 2913
rect 6273 2873 6285 2907
rect 6319 2873 6331 2907
rect 6564 2904 6592 2935
rect 6730 2932 6736 2984
rect 6788 2932 6794 2984
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 7006 2904 7012 2916
rect 6564 2876 7012 2904
rect 6273 2867 6331 2873
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7116 2904 7144 3012
rect 7208 3012 8116 3040
rect 7208 2981 7236 3012
rect 8110 3000 8116 3012
rect 8168 3040 8174 3052
rect 9030 3040 9036 3052
rect 8168 3012 9036 3040
rect 8168 3000 8174 3012
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9508 3040 9536 3148
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 18785 3179 18843 3185
rect 18785 3145 18797 3179
rect 18831 3176 18843 3179
rect 19058 3176 19064 3188
rect 18831 3148 19064 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 22094 3136 22100 3188
rect 22152 3176 22158 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 22152 3148 22201 3176
rect 22152 3136 22158 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 22189 3139 22247 3145
rect 22278 3136 22284 3188
rect 22336 3136 22342 3188
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 27062 3176 27068 3188
rect 26568 3148 27068 3176
rect 26568 3136 26574 3148
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 28350 3136 28356 3188
rect 28408 3136 28414 3188
rect 30374 3136 30380 3188
rect 30432 3136 30438 3188
rect 10502 3068 10508 3120
rect 10560 3068 10566 3120
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 14090 3108 14096 3120
rect 11848 3080 14096 3108
rect 11848 3068 11854 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 26694 3068 26700 3120
rect 26752 3068 26758 3120
rect 9232 3012 9536 3040
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 8938 2932 8944 2984
rect 8996 2932 9002 2984
rect 9232 2981 9260 3012
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9640 3012 9965 3040
rect 9640 3000 9646 3012
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 13170 3040 13176 3052
rect 12584 3012 13176 3040
rect 12584 3000 12590 3012
rect 13170 3000 13176 3012
rect 13228 3040 13234 3052
rect 15010 3040 15016 3052
rect 13228 3012 15016 3040
rect 13228 3000 13234 3012
rect 10134 2981 10140 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 10112 2975 10140 2981
rect 10112 2941 10124 2975
rect 10112 2935 10140 2941
rect 10134 2932 10140 2935
rect 10192 2932 10198 2984
rect 10226 2932 10232 2984
rect 10284 2932 10290 2984
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2941 11023 2975
rect 10965 2935 11023 2941
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11238 2972 11244 2984
rect 11195 2944 11244 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 8478 2904 8484 2916
rect 7116 2876 8484 2904
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 5994 2845 6000 2848
rect 5261 2839 5319 2845
rect 5261 2836 5273 2839
rect 5224 2808 5273 2836
rect 5224 2796 5230 2808
rect 5261 2805 5273 2808
rect 5307 2805 5319 2839
rect 5261 2799 5319 2805
rect 5813 2839 5871 2845
rect 5813 2805 5825 2839
rect 5859 2805 5871 2839
rect 5813 2799 5871 2805
rect 5981 2839 6000 2845
rect 5981 2805 5993 2839
rect 5981 2799 6000 2805
rect 5994 2796 6000 2799
rect 6052 2796 6058 2848
rect 6825 2839 6883 2845
rect 6825 2805 6837 2839
rect 6871 2836 6883 2839
rect 7098 2836 7104 2848
rect 6871 2808 7104 2836
rect 6871 2805 6883 2808
rect 6825 2799 6883 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 8570 2796 8576 2848
rect 8628 2796 8634 2848
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2836 9091 2839
rect 10042 2836 10048 2848
rect 9079 2808 10048 2836
rect 9079 2805 9091 2808
rect 9033 2799 9091 2805
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 10980 2836 11008 2935
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 11330 2932 11336 2984
rect 11388 2972 11394 2984
rect 12618 2972 12624 2984
rect 11388 2944 12624 2972
rect 11388 2932 11394 2944
rect 12618 2932 12624 2944
rect 12676 2972 12682 2984
rect 13372 2981 13400 3012
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 20714 3040 20720 3052
rect 20548 3012 20720 3040
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12676 2944 12817 2972
rect 12676 2932 12682 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 13357 2975 13415 2981
rect 13357 2941 13369 2975
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 14090 2932 14096 2984
rect 14148 2932 14154 2984
rect 14366 2932 14372 2984
rect 14424 2932 14430 2984
rect 18598 2932 18604 2984
rect 18656 2972 18662 2984
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18656 2944 18705 2972
rect 18656 2932 18662 2944
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 18693 2935 18751 2941
rect 20346 2932 20352 2984
rect 20404 2972 20410 2984
rect 20548 2981 20576 3012
rect 20714 3000 20720 3012
rect 20772 3040 20778 3052
rect 24394 3040 24400 3052
rect 20772 3012 20935 3040
rect 20772 3000 20778 3012
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 20404 2944 20545 2972
rect 20404 2932 20410 2944
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 20625 2975 20683 2981
rect 20625 2941 20637 2975
rect 20671 2972 20683 2975
rect 20809 2975 20867 2981
rect 20809 2972 20821 2975
rect 20671 2944 20821 2972
rect 20671 2941 20683 2944
rect 20625 2935 20683 2941
rect 20809 2941 20821 2944
rect 20855 2941 20867 2975
rect 20907 2972 20935 3012
rect 23584 3012 24400 3040
rect 23584 2972 23612 3012
rect 24394 3000 24400 3012
rect 24452 3000 24458 3052
rect 27430 3040 27436 3052
rect 26988 3012 27436 3040
rect 20907 2944 23612 2972
rect 20809 2935 20867 2941
rect 23658 2932 23664 2984
rect 23716 2932 23722 2984
rect 23845 2975 23903 2981
rect 23845 2941 23857 2975
rect 23891 2941 23903 2975
rect 26602 2972 26608 2984
rect 26560 2947 26608 2972
rect 23845 2935 23903 2941
rect 26559 2941 26608 2947
rect 11256 2904 11284 2932
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 11256 2876 12909 2904
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 13081 2907 13139 2913
rect 13081 2873 13093 2907
rect 13127 2904 13139 2907
rect 13722 2904 13728 2916
rect 13127 2876 13728 2904
rect 13127 2873 13139 2876
rect 13081 2867 13139 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 14108 2904 14136 2932
rect 14826 2904 14832 2916
rect 14108 2876 14832 2904
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 21076 2907 21134 2913
rect 21076 2873 21088 2907
rect 21122 2904 21134 2907
rect 21266 2904 21272 2916
rect 21122 2876 21272 2904
rect 21122 2873 21134 2876
rect 21076 2867 21134 2873
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 22066 2876 22416 2904
rect 11330 2836 11336 2848
rect 10376 2808 11336 2836
rect 10376 2796 10382 2808
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 12492 2808 12817 2836
rect 12492 2796 12498 2808
rect 12805 2805 12817 2808
rect 12851 2805 12863 2839
rect 12805 2799 12863 2805
rect 12986 2796 12992 2848
rect 13044 2836 13050 2848
rect 13265 2839 13323 2845
rect 13265 2836 13277 2839
rect 13044 2808 13277 2836
rect 13044 2796 13050 2808
rect 13265 2805 13277 2808
rect 13311 2805 13323 2839
rect 13265 2799 13323 2805
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 22066 2836 22094 2876
rect 17000 2808 22094 2836
rect 22388 2836 22416 2876
rect 23290 2864 23296 2916
rect 23348 2904 23354 2916
rect 23394 2907 23452 2913
rect 23394 2904 23406 2907
rect 23348 2876 23406 2904
rect 23348 2864 23354 2876
rect 23394 2873 23406 2876
rect 23440 2873 23452 2907
rect 23394 2867 23452 2873
rect 23860 2836 23888 2935
rect 26142 2864 26148 2916
rect 26200 2904 26206 2916
rect 26329 2907 26387 2913
rect 26329 2904 26341 2907
rect 26200 2876 26341 2904
rect 26200 2864 26206 2876
rect 26329 2873 26341 2876
rect 26375 2873 26387 2907
rect 26559 2907 26571 2941
rect 26605 2932 26608 2941
rect 26660 2972 26666 2984
rect 26988 2981 27016 3012
rect 27430 3000 27436 3012
rect 27488 3040 27494 3052
rect 27985 3043 28043 3049
rect 27985 3040 27997 3043
rect 27488 3012 27997 3040
rect 27488 3000 27494 3012
rect 27985 3009 27997 3012
rect 28031 3009 28043 3043
rect 27985 3003 28043 3009
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26660 2944 26985 2972
rect 26660 2932 26666 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 27062 2932 27068 2984
rect 27120 2932 27126 2984
rect 28074 2932 28080 2984
rect 28132 2972 28138 2984
rect 28629 2975 28687 2981
rect 28629 2972 28641 2975
rect 28132 2944 28641 2972
rect 28132 2932 28138 2944
rect 28629 2941 28641 2944
rect 28675 2941 28687 2975
rect 28629 2935 28687 2941
rect 28721 2975 28779 2981
rect 28721 2941 28733 2975
rect 28767 2972 28779 2975
rect 28997 2975 29055 2981
rect 28997 2972 29009 2975
rect 28767 2944 29009 2972
rect 28767 2941 28779 2944
rect 28721 2935 28779 2941
rect 28997 2941 29009 2944
rect 29043 2941 29055 2975
rect 28997 2935 29055 2941
rect 26605 2907 26617 2932
rect 26559 2901 26617 2907
rect 26329 2867 26387 2873
rect 22388 2808 23888 2836
rect 17000 2796 17006 2808
rect 24026 2796 24032 2848
rect 24084 2796 24090 2848
rect 24118 2796 24124 2848
rect 24176 2836 24182 2848
rect 25130 2836 25136 2848
rect 24176 2808 25136 2836
rect 24176 2796 24182 2808
rect 25130 2796 25136 2808
rect 25188 2796 25194 2848
rect 26344 2836 26372 2867
rect 26786 2864 26792 2916
rect 26844 2904 26850 2916
rect 27249 2907 27307 2913
rect 27249 2904 27261 2907
rect 26844 2876 27261 2904
rect 26844 2864 26850 2876
rect 27249 2873 27261 2876
rect 27295 2873 27307 2907
rect 27249 2867 27307 2873
rect 27433 2907 27491 2913
rect 27433 2873 27445 2907
rect 27479 2873 27491 2907
rect 27433 2867 27491 2873
rect 27448 2836 27476 2867
rect 28258 2864 28264 2916
rect 28316 2904 28322 2916
rect 28353 2907 28411 2913
rect 28353 2904 28365 2907
rect 28316 2876 28365 2904
rect 28316 2864 28322 2876
rect 28353 2873 28365 2876
rect 28399 2904 28411 2907
rect 28442 2904 28448 2916
rect 28399 2876 28448 2904
rect 28399 2873 28411 2876
rect 28353 2867 28411 2873
rect 28442 2864 28448 2876
rect 28500 2864 28506 2916
rect 29242 2907 29300 2913
rect 29242 2904 29254 2907
rect 28552 2876 29254 2904
rect 26344 2808 27476 2836
rect 27617 2839 27675 2845
rect 27617 2805 27629 2839
rect 27663 2836 27675 2839
rect 27982 2836 27988 2848
rect 27663 2808 27988 2836
rect 27663 2805 27675 2808
rect 27617 2799 27675 2805
rect 27982 2796 27988 2808
rect 28040 2796 28046 2848
rect 28552 2845 28580 2876
rect 29242 2873 29254 2876
rect 29288 2873 29300 2907
rect 29242 2867 29300 2873
rect 28537 2839 28595 2845
rect 28537 2805 28549 2839
rect 28583 2805 28595 2839
rect 28537 2799 28595 2805
rect 552 2746 31648 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 12096 2746
rect 12148 2694 12160 2746
rect 12212 2694 12224 2746
rect 12276 2694 12288 2746
rect 12340 2694 12352 2746
rect 12404 2694 19870 2746
rect 19922 2694 19934 2746
rect 19986 2694 19998 2746
rect 20050 2694 20062 2746
rect 20114 2694 20126 2746
rect 20178 2694 27644 2746
rect 27696 2694 27708 2746
rect 27760 2694 27772 2746
rect 27824 2694 27836 2746
rect 27888 2694 27900 2746
rect 27952 2694 31648 2746
rect 552 2672 31648 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 3016 2604 3249 2632
rect 3016 2592 3022 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3237 2595 3295 2601
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6454 2632 6460 2644
rect 5951 2604 6460 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 3418 2456 3424 2508
rect 3476 2456 3482 2508
rect 3510 2456 3516 2508
rect 3568 2456 3574 2508
rect 5442 2456 5448 2508
rect 5500 2456 5506 2508
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 5920 2496 5948 2595
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7006 2592 7012 2644
rect 7064 2592 7070 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9582 2632 9588 2644
rect 9171 2604 9588 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10042 2592 10048 2644
rect 10100 2592 10106 2644
rect 10962 2592 10968 2644
rect 11020 2592 11026 2644
rect 12805 2635 12863 2641
rect 12805 2601 12817 2635
rect 12851 2601 12863 2635
rect 12805 2595 12863 2601
rect 6730 2564 6736 2576
rect 6104 2536 6736 2564
rect 5675 2468 5948 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6104 2505 6132 2536
rect 6730 2524 6736 2536
rect 6788 2524 6794 2576
rect 9858 2524 9864 2576
rect 9916 2564 9922 2576
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9916 2536 9965 2564
rect 9916 2524 9922 2536
rect 9953 2533 9965 2536
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 10226 2524 10232 2576
rect 10284 2564 10290 2576
rect 10284 2536 11468 2564
rect 10284 2524 10290 2536
rect 6089 2499 6147 2505
rect 6089 2496 6101 2499
rect 6052 2468 6101 2496
rect 6052 2456 6058 2468
rect 6089 2465 6101 2468
rect 6135 2465 6147 2499
rect 6089 2459 6147 2465
rect 6362 2456 6368 2508
rect 6420 2456 6426 2508
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 11238 2496 11244 2508
rect 9815 2468 11244 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 4062 2428 4068 2440
rect 3283 2400 4068 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 4062 2388 4068 2400
rect 4120 2428 4126 2440
rect 5810 2428 5816 2440
rect 4120 2400 5816 2428
rect 4120 2388 4126 2400
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 6086 2320 6092 2372
rect 6144 2360 6150 2372
rect 6288 2360 6316 2391
rect 7282 2388 7288 2440
rect 7340 2388 7346 2440
rect 7466 2388 7472 2440
rect 7524 2388 7530 2440
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 8036 2400 8217 2428
rect 6822 2360 6828 2372
rect 6144 2332 6828 2360
rect 6144 2320 6150 2332
rect 6822 2320 6828 2332
rect 6880 2360 6886 2372
rect 8036 2360 8064 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8294 2388 8300 2440
rect 8352 2437 8358 2440
rect 8352 2431 8380 2437
rect 8368 2397 8380 2431
rect 8352 2391 8380 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 9122 2428 9128 2440
rect 8527 2400 9128 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8352 2388 8358 2391
rect 9122 2388 9128 2400
rect 9180 2428 9186 2440
rect 9490 2428 9496 2440
rect 9180 2400 9496 2428
rect 9180 2388 9186 2400
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 6880 2332 8064 2360
rect 6880 2320 6886 2332
rect 4706 2252 4712 2304
rect 4764 2292 4770 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 4764 2264 5457 2292
rect 4764 2252 4770 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9398 2292 9404 2304
rect 8996 2264 9404 2292
rect 8996 2252 9002 2264
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 9600 2292 9628 2459
rect 9692 2360 9720 2459
rect 11238 2456 11244 2468
rect 11296 2456 11302 2508
rect 11330 2456 11336 2508
rect 11388 2456 11394 2508
rect 11440 2505 11468 2536
rect 12434 2524 12440 2576
rect 12492 2524 12498 2576
rect 12637 2567 12695 2573
rect 12637 2533 12649 2567
rect 12683 2564 12695 2567
rect 12820 2564 12848 2595
rect 13722 2592 13728 2644
rect 13780 2632 13786 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 13780 2604 14289 2632
rect 13780 2592 13786 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 15010 2592 15016 2644
rect 15068 2592 15074 2644
rect 17218 2632 17224 2644
rect 16776 2604 17224 2632
rect 13142 2567 13200 2573
rect 13142 2564 13154 2567
rect 12683 2536 12756 2564
rect 12820 2536 13154 2564
rect 12683 2533 12695 2536
rect 12637 2527 12695 2533
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 12728 2496 12756 2536
rect 13142 2533 13154 2536
rect 13188 2533 13200 2567
rect 15028 2564 15056 2592
rect 13142 2527 13200 2533
rect 14568 2536 16252 2564
rect 12802 2496 12808 2508
rect 12728 2468 12808 2496
rect 11425 2459 11483 2465
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2496 12955 2499
rect 12986 2496 12992 2508
rect 12943 2468 12992 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 12986 2456 12992 2468
rect 13044 2456 13050 2508
rect 14568 2505 14596 2536
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 15013 2499 15071 2505
rect 15013 2465 15025 2499
rect 15059 2496 15071 2499
rect 15120 2496 15148 2536
rect 15059 2468 15148 2496
rect 15059 2465 15071 2468
rect 15013 2459 15071 2465
rect 15562 2456 15568 2508
rect 15620 2456 15626 2508
rect 16224 2505 16252 2536
rect 16776 2505 16804 2604
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 18325 2635 18383 2641
rect 18325 2601 18337 2635
rect 18371 2632 18383 2635
rect 18874 2632 18880 2644
rect 18371 2604 18880 2632
rect 18371 2601 18383 2604
rect 18325 2595 18383 2601
rect 18874 2592 18880 2604
rect 18932 2632 18938 2644
rect 19521 2635 19579 2641
rect 19521 2632 19533 2635
rect 18932 2604 19533 2632
rect 18932 2592 18938 2604
rect 19521 2601 19533 2604
rect 19567 2632 19579 2635
rect 19702 2632 19708 2644
rect 19567 2604 19708 2632
rect 19567 2601 19579 2604
rect 19521 2595 19579 2601
rect 19702 2592 19708 2604
rect 19760 2592 19766 2644
rect 21266 2592 21272 2644
rect 21324 2592 21330 2644
rect 26694 2632 26700 2644
rect 26068 2604 26700 2632
rect 18233 2567 18291 2573
rect 16868 2536 17816 2564
rect 16868 2505 16896 2536
rect 16209 2499 16267 2505
rect 16209 2465 16221 2499
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2465 17003 2499
rect 16945 2459 17003 2465
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2397 11207 2431
rect 11256 2428 11284 2456
rect 11882 2428 11888 2440
rect 11256 2400 11888 2428
rect 11149 2391 11207 2397
rect 10134 2360 10140 2372
rect 9692 2332 10140 2360
rect 10134 2320 10140 2332
rect 10192 2360 10198 2372
rect 11164 2360 11192 2391
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 16960 2428 16988 2459
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 17092 2468 17141 2496
rect 17092 2456 17098 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 17218 2456 17224 2508
rect 17276 2456 17282 2508
rect 17420 2505 17448 2536
rect 17788 2505 17816 2536
rect 18233 2533 18245 2567
rect 18279 2564 18291 2567
rect 18782 2564 18788 2576
rect 18279 2536 18788 2564
rect 18279 2533 18291 2536
rect 18233 2527 18291 2533
rect 18782 2524 18788 2536
rect 18840 2564 18846 2576
rect 23109 2567 23167 2573
rect 18840 2536 19656 2564
rect 18840 2524 18846 2536
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2465 17463 2499
rect 17405 2459 17463 2465
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18049 2499 18107 2505
rect 18049 2496 18061 2499
rect 17819 2468 18061 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18049 2465 18061 2468
rect 18095 2465 18107 2499
rect 18049 2459 18107 2465
rect 17313 2431 17371 2437
rect 17313 2428 17325 2431
rect 15703 2400 17325 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 17313 2397 17325 2400
rect 17359 2397 17371 2431
rect 17696 2428 17724 2459
rect 18414 2456 18420 2508
rect 18472 2496 18478 2508
rect 18966 2496 18972 2508
rect 18472 2468 18972 2496
rect 18472 2456 18478 2468
rect 18966 2456 18972 2468
rect 19024 2496 19030 2508
rect 19628 2505 19656 2536
rect 21560 2536 22048 2564
rect 19337 2499 19395 2505
rect 19337 2496 19349 2499
rect 19024 2468 19349 2496
rect 19024 2456 19030 2468
rect 19337 2465 19349 2468
rect 19383 2465 19395 2499
rect 19337 2459 19395 2465
rect 19613 2499 19671 2505
rect 19613 2465 19625 2499
rect 19659 2496 19671 2499
rect 20898 2496 20904 2508
rect 19659 2468 20904 2496
rect 19659 2465 19671 2468
rect 19613 2459 19671 2465
rect 20898 2456 20904 2468
rect 20956 2456 20962 2508
rect 21560 2505 21588 2536
rect 21545 2499 21603 2505
rect 21545 2465 21557 2499
rect 21591 2465 21603 2499
rect 21545 2459 21603 2465
rect 21634 2456 21640 2508
rect 21692 2456 21698 2508
rect 22020 2505 22048 2536
rect 23109 2533 23121 2567
rect 23155 2564 23167 2567
rect 24305 2567 24363 2573
rect 23155 2536 24256 2564
rect 23155 2533 23167 2536
rect 23109 2527 23167 2533
rect 21729 2499 21787 2505
rect 21729 2465 21741 2499
rect 21775 2465 21787 2499
rect 21913 2499 21971 2505
rect 21913 2496 21925 2499
rect 21729 2459 21787 2465
rect 21836 2468 21925 2496
rect 18322 2428 18328 2440
rect 17696 2400 18328 2428
rect 17313 2391 17371 2397
rect 18322 2388 18328 2400
rect 18380 2428 18386 2440
rect 20346 2428 20352 2440
rect 18380 2400 20352 2428
rect 18380 2388 18386 2400
rect 20346 2388 20352 2400
rect 20404 2388 20410 2440
rect 10192 2332 12940 2360
rect 10192 2320 10198 2332
rect 10226 2292 10232 2304
rect 9600 2264 10232 2292
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 11790 2252 11796 2304
rect 11848 2292 11854 2304
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 11848 2264 12633 2292
rect 11848 2252 11854 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 12912 2292 12940 2332
rect 14090 2320 14096 2372
rect 14148 2360 14154 2372
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 14148 2332 14473 2360
rect 14148 2320 14154 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 14461 2323 14519 2329
rect 17126 2320 17132 2372
rect 17184 2360 17190 2372
rect 17589 2363 17647 2369
rect 17589 2360 17601 2363
rect 17184 2332 17601 2360
rect 17184 2320 17190 2332
rect 17589 2329 17601 2332
rect 17635 2329 17647 2363
rect 17589 2323 17647 2329
rect 18598 2320 18604 2372
rect 18656 2320 18662 2372
rect 20993 2363 21051 2369
rect 20993 2329 21005 2363
rect 21039 2360 21051 2363
rect 21744 2360 21772 2459
rect 21039 2332 21772 2360
rect 21836 2360 21864 2468
rect 21913 2465 21925 2468
rect 21959 2465 21971 2499
rect 21913 2459 21971 2465
rect 22005 2499 22063 2505
rect 22005 2465 22017 2499
rect 22051 2465 22063 2499
rect 22005 2459 22063 2465
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 22557 2499 22615 2505
rect 22557 2496 22569 2499
rect 22244 2468 22569 2496
rect 22244 2456 22250 2468
rect 22557 2465 22569 2468
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 22646 2456 22652 2508
rect 22704 2496 22710 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 22704 2468 22753 2496
rect 22704 2456 22710 2468
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 22741 2459 22799 2465
rect 23661 2499 23719 2505
rect 23661 2465 23673 2499
rect 23707 2496 23719 2499
rect 23750 2496 23756 2508
rect 23707 2468 23756 2496
rect 23707 2465 23719 2468
rect 23661 2459 23719 2465
rect 23750 2456 23756 2468
rect 23808 2456 23814 2508
rect 23934 2456 23940 2508
rect 23992 2456 23998 2508
rect 24118 2456 24124 2508
rect 24176 2456 24182 2508
rect 23106 2388 23112 2440
rect 23164 2428 23170 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 23164 2400 23489 2428
rect 23164 2388 23170 2400
rect 23477 2397 23489 2400
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 24136 2428 24164 2456
rect 23891 2400 24164 2428
rect 24228 2428 24256 2536
rect 24305 2533 24317 2567
rect 24351 2564 24363 2567
rect 24486 2564 24492 2576
rect 24351 2536 24492 2564
rect 24351 2533 24363 2536
rect 24305 2527 24363 2533
rect 24486 2524 24492 2536
rect 24544 2524 24550 2576
rect 26068 2573 26096 2604
rect 26694 2592 26700 2604
rect 26752 2592 26758 2644
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 28258 2632 28264 2644
rect 26936 2604 28264 2632
rect 26936 2592 26942 2604
rect 28258 2592 28264 2604
rect 28316 2592 28322 2644
rect 24765 2567 24823 2573
rect 24765 2564 24777 2567
rect 24596 2536 24777 2564
rect 24394 2456 24400 2508
rect 24452 2456 24458 2508
rect 24596 2496 24624 2536
rect 24765 2533 24777 2536
rect 24811 2533 24823 2567
rect 24765 2527 24823 2533
rect 26053 2567 26111 2573
rect 26053 2533 26065 2567
rect 26099 2533 26111 2567
rect 26053 2527 26111 2533
rect 26510 2524 26516 2576
rect 26568 2564 26574 2576
rect 27157 2567 27215 2573
rect 27157 2564 27169 2567
rect 26568 2536 27169 2564
rect 26568 2524 26574 2536
rect 27157 2533 27169 2536
rect 27203 2533 27215 2567
rect 27157 2527 27215 2533
rect 27430 2524 27436 2576
rect 27488 2564 27494 2576
rect 27801 2567 27859 2573
rect 27801 2564 27813 2567
rect 27488 2536 27813 2564
rect 27488 2524 27494 2536
rect 27801 2533 27813 2536
rect 27847 2533 27859 2567
rect 27801 2527 27859 2533
rect 24504 2468 24624 2496
rect 24504 2428 24532 2468
rect 24670 2456 24676 2508
rect 24728 2456 24734 2508
rect 24854 2456 24860 2508
rect 24912 2456 24918 2508
rect 24949 2499 25007 2505
rect 24949 2465 24961 2499
rect 24995 2496 25007 2499
rect 25225 2499 25283 2505
rect 25225 2496 25237 2499
rect 24995 2468 25237 2496
rect 24995 2465 25007 2468
rect 24949 2459 25007 2465
rect 25225 2465 25237 2468
rect 25271 2465 25283 2499
rect 25225 2459 25283 2465
rect 24228 2400 24532 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24578 2388 24584 2440
rect 24636 2428 24642 2440
rect 24964 2428 24992 2459
rect 24636 2400 24992 2428
rect 25240 2428 25268 2459
rect 25314 2456 25320 2508
rect 25372 2496 25378 2508
rect 25774 2496 25780 2508
rect 25372 2468 25780 2496
rect 25372 2456 25378 2468
rect 25774 2456 25780 2468
rect 25832 2496 25838 2508
rect 25869 2499 25927 2505
rect 25869 2496 25881 2499
rect 25832 2468 25881 2496
rect 25832 2456 25838 2468
rect 25869 2465 25881 2468
rect 25915 2465 25927 2499
rect 25869 2459 25927 2465
rect 26697 2499 26755 2505
rect 26697 2465 26709 2499
rect 26743 2465 26755 2499
rect 26697 2459 26755 2465
rect 26712 2428 26740 2459
rect 27062 2456 27068 2508
rect 27120 2496 27126 2508
rect 27614 2496 27620 2508
rect 27120 2468 27620 2496
rect 27120 2456 27126 2468
rect 27614 2456 27620 2468
rect 27672 2456 27678 2508
rect 28074 2428 28080 2440
rect 25240 2400 28080 2428
rect 24636 2388 24642 2400
rect 28074 2388 28080 2400
rect 28132 2388 28138 2440
rect 21836 2332 23060 2360
rect 21039 2329 21051 2332
rect 20993 2323 21051 2329
rect 13630 2292 13636 2304
rect 12912 2264 13636 2292
rect 12621 2255 12679 2261
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 15105 2295 15163 2301
rect 15105 2261 15117 2295
rect 15151 2292 15163 2295
rect 15286 2292 15292 2304
rect 15151 2264 15292 2292
rect 15151 2261 15163 2264
rect 15105 2255 15163 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 15746 2252 15752 2304
rect 15804 2292 15810 2304
rect 15841 2295 15899 2301
rect 15841 2292 15853 2295
rect 15804 2264 15853 2292
rect 15804 2252 15810 2264
rect 15841 2261 15853 2264
rect 15887 2261 15899 2295
rect 15841 2255 15899 2261
rect 16298 2252 16304 2304
rect 16356 2252 16362 2304
rect 16482 2252 16488 2304
rect 16540 2252 16546 2304
rect 17862 2252 17868 2304
rect 17920 2252 17926 2304
rect 19058 2252 19064 2304
rect 19116 2292 19122 2304
rect 19153 2295 19211 2301
rect 19153 2292 19165 2295
rect 19116 2264 19165 2292
rect 19116 2252 19122 2264
rect 19153 2261 19165 2264
rect 19199 2261 19211 2295
rect 19153 2255 19211 2261
rect 20070 2252 20076 2304
rect 20128 2292 20134 2304
rect 21836 2292 21864 2332
rect 23032 2304 23060 2332
rect 23290 2320 23296 2372
rect 23348 2320 23354 2372
rect 23658 2320 23664 2372
rect 23716 2360 23722 2372
rect 24489 2363 24547 2369
rect 24489 2360 24501 2363
rect 23716 2332 24501 2360
rect 23716 2320 23722 2332
rect 24489 2329 24501 2332
rect 24535 2329 24547 2363
rect 25130 2360 25136 2372
rect 24489 2323 24547 2329
rect 24596 2332 25136 2360
rect 20128 2264 21864 2292
rect 20128 2252 20134 2264
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 23072 2264 23121 2292
rect 23072 2252 23078 2264
rect 23109 2261 23121 2264
rect 23155 2292 23167 2295
rect 24596 2292 24624 2332
rect 25130 2320 25136 2332
rect 25188 2320 25194 2372
rect 25317 2363 25375 2369
rect 25317 2329 25329 2363
rect 25363 2360 25375 2363
rect 26234 2360 26240 2372
rect 25363 2332 26240 2360
rect 25363 2329 25375 2332
rect 25317 2323 25375 2329
rect 26234 2320 26240 2332
rect 26292 2320 26298 2372
rect 26694 2320 26700 2372
rect 26752 2360 26758 2372
rect 26789 2363 26847 2369
rect 26789 2360 26801 2363
rect 26752 2332 26801 2360
rect 26752 2320 26758 2332
rect 26789 2329 26801 2332
rect 26835 2329 26847 2363
rect 27982 2360 27988 2372
rect 26789 2323 26847 2329
rect 27172 2332 27988 2360
rect 23155 2264 24624 2292
rect 25041 2295 25099 2301
rect 23155 2261 23167 2264
rect 23109 2255 23167 2261
rect 25041 2261 25053 2295
rect 25087 2292 25099 2295
rect 25222 2292 25228 2304
rect 25087 2264 25228 2292
rect 25087 2261 25099 2264
rect 25041 2255 25099 2261
rect 25222 2252 25228 2264
rect 25280 2252 25286 2304
rect 25682 2252 25688 2304
rect 25740 2252 25746 2304
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27172 2301 27200 2332
rect 27982 2320 27988 2332
rect 28040 2320 28046 2372
rect 26605 2295 26663 2301
rect 26605 2292 26617 2295
rect 26476 2264 26617 2292
rect 26476 2252 26482 2264
rect 26605 2261 26617 2264
rect 26651 2261 26663 2295
rect 26605 2255 26663 2261
rect 27157 2295 27215 2301
rect 27157 2261 27169 2295
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27338 2252 27344 2304
rect 27396 2252 27402 2304
rect 27430 2252 27436 2304
rect 27488 2252 27494 2304
rect 552 2202 31648 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 11436 2202
rect 11488 2150 11500 2202
rect 11552 2150 11564 2202
rect 11616 2150 11628 2202
rect 11680 2150 11692 2202
rect 11744 2150 19210 2202
rect 19262 2150 19274 2202
rect 19326 2150 19338 2202
rect 19390 2150 19402 2202
rect 19454 2150 19466 2202
rect 19518 2150 26984 2202
rect 27036 2150 27048 2202
rect 27100 2150 27112 2202
rect 27164 2150 27176 2202
rect 27228 2150 27240 2202
rect 27292 2150 31648 2202
rect 552 2128 31648 2150
rect 6273 2091 6331 2097
rect 6273 2057 6285 2091
rect 6319 2088 6331 2091
rect 6362 2088 6368 2100
rect 6319 2060 6368 2088
rect 6319 2057 6331 2060
rect 6273 2051 6331 2057
rect 6362 2048 6368 2060
rect 6420 2048 6426 2100
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 8018 2088 8024 2100
rect 7340 2060 8024 2088
rect 7340 2048 7346 2060
rect 8018 2048 8024 2060
rect 8076 2088 8082 2100
rect 8389 2091 8447 2097
rect 8389 2088 8401 2091
rect 8076 2060 8401 2088
rect 8076 2048 8082 2060
rect 8389 2057 8401 2060
rect 8435 2057 8447 2091
rect 8389 2051 8447 2057
rect 9953 2091 10011 2097
rect 9953 2057 9965 2091
rect 9999 2088 10011 2091
rect 10226 2088 10232 2100
rect 9999 2060 10232 2088
rect 9999 2057 10011 2060
rect 9953 2051 10011 2057
rect 10226 2048 10232 2060
rect 10284 2048 10290 2100
rect 10410 2048 10416 2100
rect 10468 2088 10474 2100
rect 11609 2091 11667 2097
rect 11609 2088 11621 2091
rect 10468 2060 11621 2088
rect 10468 2048 10474 2060
rect 11609 2057 11621 2060
rect 11655 2057 11667 2091
rect 11609 2051 11667 2057
rect 11882 2048 11888 2100
rect 11940 2088 11946 2100
rect 12342 2088 12348 2100
rect 11940 2060 12348 2088
rect 11940 2048 11946 2060
rect 12342 2048 12348 2060
rect 12400 2088 12406 2100
rect 12400 2060 12848 2088
rect 12400 2048 12406 2060
rect 12621 2023 12679 2029
rect 11348 1992 11928 2020
rect 6822 1912 6828 1964
rect 6880 1952 6886 1964
rect 6917 1955 6975 1961
rect 6917 1952 6929 1955
rect 6880 1924 6929 1952
rect 6880 1912 6886 1924
rect 6917 1921 6929 1924
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 8021 1955 8079 1961
rect 8021 1921 8033 1955
rect 8067 1952 8079 1955
rect 8294 1952 8300 1964
rect 8067 1924 8300 1952
rect 8067 1921 8079 1924
rect 8021 1915 8079 1921
rect 8294 1912 8300 1924
rect 8352 1912 8358 1964
rect 5166 1893 5172 1896
rect 4525 1887 4583 1893
rect 4525 1853 4537 1887
rect 4571 1884 4583 1887
rect 4617 1887 4675 1893
rect 4617 1884 4629 1887
rect 4571 1856 4629 1884
rect 4571 1853 4583 1856
rect 4525 1847 4583 1853
rect 4617 1853 4629 1856
rect 4663 1853 4675 1887
rect 4617 1847 4675 1853
rect 4709 1887 4767 1893
rect 4709 1853 4721 1887
rect 4755 1884 4767 1887
rect 4893 1887 4951 1893
rect 4893 1884 4905 1887
rect 4755 1856 4905 1884
rect 4755 1853 4767 1856
rect 4709 1847 4767 1853
rect 4893 1853 4905 1856
rect 4939 1853 4951 1887
rect 4893 1847 4951 1853
rect 5160 1847 5172 1893
rect 4632 1816 4660 1847
rect 5166 1844 5172 1847
rect 5224 1844 5230 1896
rect 9766 1844 9772 1896
rect 9824 1844 9830 1896
rect 11054 1844 11060 1896
rect 11112 1893 11118 1896
rect 11348 1893 11376 1992
rect 11701 1955 11759 1961
rect 11701 1921 11713 1955
rect 11747 1952 11759 1955
rect 11790 1952 11796 1964
rect 11747 1924 11796 1952
rect 11747 1921 11759 1924
rect 11701 1915 11759 1921
rect 11790 1912 11796 1924
rect 11848 1912 11854 1964
rect 11900 1961 11928 1992
rect 12621 1989 12633 2023
rect 12667 2020 12679 2023
rect 12667 1992 12756 2020
rect 12667 1989 12679 1992
rect 12621 1983 12679 1989
rect 11885 1955 11943 1961
rect 11885 1921 11897 1955
rect 11931 1921 11943 1955
rect 12526 1952 12532 1964
rect 11885 1915 11943 1921
rect 12084 1924 12532 1952
rect 12084 1893 12112 1924
rect 12526 1912 12532 1924
rect 12584 1912 12590 1964
rect 12728 1961 12756 1992
rect 12713 1955 12771 1961
rect 12713 1921 12725 1955
rect 12759 1921 12771 1955
rect 12820 1952 12848 2060
rect 12894 2048 12900 2100
rect 12952 2088 12958 2100
rect 13541 2091 13599 2097
rect 13541 2088 13553 2091
rect 12952 2060 13553 2088
rect 12952 2048 12958 2060
rect 13541 2057 13553 2060
rect 13587 2057 13599 2091
rect 13541 2051 13599 2057
rect 13630 2048 13636 2100
rect 13688 2088 13694 2100
rect 13688 2060 14964 2088
rect 13688 2048 13694 2060
rect 14936 2029 14964 2060
rect 15562 2048 15568 2100
rect 15620 2088 15626 2100
rect 16669 2091 16727 2097
rect 16669 2088 16681 2091
rect 15620 2060 16681 2088
rect 15620 2048 15626 2060
rect 16669 2057 16681 2060
rect 16715 2057 16727 2091
rect 16669 2051 16727 2057
rect 18509 2091 18567 2097
rect 18509 2057 18521 2091
rect 18555 2088 18567 2091
rect 18598 2088 18604 2100
rect 18555 2060 18604 2088
rect 18555 2057 18567 2060
rect 18509 2051 18567 2057
rect 18598 2048 18604 2060
rect 18656 2088 18662 2100
rect 24210 2088 24216 2100
rect 18656 2060 19288 2088
rect 18656 2048 18662 2060
rect 14921 2023 14979 2029
rect 14921 1989 14933 2023
rect 14967 1989 14979 2023
rect 14921 1983 14979 1989
rect 13648 1952 13768 1960
rect 12820 1932 14780 1952
rect 12820 1924 13676 1932
rect 13740 1924 14780 1932
rect 12713 1915 12771 1921
rect 14016 1896 14044 1924
rect 11112 1847 11124 1893
rect 11333 1887 11391 1893
rect 11333 1853 11345 1887
rect 11379 1853 11391 1887
rect 11333 1847 11391 1853
rect 11425 1887 11483 1893
rect 11425 1853 11437 1887
rect 11471 1853 11483 1887
rect 11425 1847 11483 1853
rect 11517 1887 11575 1893
rect 11517 1853 11529 1887
rect 11563 1853 11575 1887
rect 11517 1847 11575 1853
rect 11977 1887 12035 1893
rect 11977 1853 11989 1887
rect 12023 1884 12035 1887
rect 12069 1887 12127 1893
rect 12069 1884 12081 1887
rect 12023 1856 12081 1884
rect 12023 1853 12035 1856
rect 11977 1847 12035 1853
rect 12069 1853 12081 1856
rect 12115 1853 12127 1887
rect 12069 1847 12127 1853
rect 11112 1844 11118 1847
rect 5074 1816 5080 1828
rect 4632 1788 5080 1816
rect 5074 1776 5080 1788
rect 5132 1776 5138 1828
rect 6086 1776 6092 1828
rect 6144 1816 6150 1828
rect 6365 1819 6423 1825
rect 6365 1816 6377 1819
rect 6144 1788 6377 1816
rect 6144 1776 6150 1788
rect 6365 1785 6377 1788
rect 6411 1785 6423 1819
rect 6365 1779 6423 1785
rect 8846 1776 8852 1828
rect 8904 1816 8910 1828
rect 9502 1819 9560 1825
rect 9502 1816 9514 1819
rect 8904 1788 9514 1816
rect 8904 1776 8910 1788
rect 9502 1785 9514 1788
rect 9548 1785 9560 1819
rect 9502 1779 9560 1785
rect 10594 1776 10600 1828
rect 10652 1816 10658 1828
rect 11440 1816 11468 1847
rect 10652 1788 11468 1816
rect 10652 1776 10658 1788
rect 4246 1708 4252 1760
rect 4304 1748 4310 1760
rect 4433 1751 4491 1757
rect 4433 1748 4445 1751
rect 4304 1720 4445 1748
rect 4304 1708 4310 1720
rect 4433 1717 4445 1720
rect 4479 1717 4491 1751
rect 4433 1711 4491 1717
rect 7098 1708 7104 1760
rect 7156 1748 7162 1760
rect 7377 1751 7435 1757
rect 7377 1748 7389 1751
rect 7156 1720 7389 1748
rect 7156 1708 7162 1720
rect 7377 1717 7389 1720
rect 7423 1717 7435 1751
rect 7377 1711 7435 1717
rect 9398 1708 9404 1760
rect 9456 1748 9462 1760
rect 11532 1748 11560 1847
rect 12342 1844 12348 1896
rect 12400 1844 12406 1896
rect 12621 1887 12679 1893
rect 12621 1853 12633 1887
rect 12667 1884 12679 1887
rect 13630 1884 13636 1896
rect 12667 1856 13636 1884
rect 12667 1853 12679 1856
rect 12621 1847 12679 1853
rect 13630 1844 13636 1856
rect 13688 1844 13694 1896
rect 13722 1844 13728 1896
rect 13780 1844 13786 1896
rect 13998 1844 14004 1896
rect 14056 1844 14062 1896
rect 14645 1887 14703 1893
rect 14645 1853 14657 1887
rect 14691 1853 14703 1887
rect 14752 1884 14780 1924
rect 14826 1912 14832 1964
rect 14884 1912 14890 1964
rect 15286 1912 15292 1964
rect 15344 1912 15350 1964
rect 16574 1912 16580 1964
rect 16632 1952 16638 1964
rect 16761 1955 16819 1961
rect 16761 1952 16773 1955
rect 16632 1924 16773 1952
rect 16632 1912 16638 1924
rect 16761 1921 16773 1924
rect 16807 1952 16819 1955
rect 17034 1952 17040 1964
rect 16807 1924 17040 1952
rect 16807 1921 16819 1924
rect 16761 1915 16819 1921
rect 17034 1912 17040 1924
rect 17092 1912 17098 1964
rect 17126 1912 17132 1964
rect 17184 1912 17190 1964
rect 19260 1961 19288 2060
rect 22756 2060 24216 2088
rect 20070 2020 20076 2032
rect 19628 1992 20076 2020
rect 19245 1955 19303 1961
rect 19245 1921 19257 1955
rect 19291 1921 19303 1955
rect 19245 1915 19303 1921
rect 15013 1887 15071 1893
rect 15013 1884 15025 1887
rect 14752 1856 15025 1884
rect 14645 1847 14703 1853
rect 15013 1853 15025 1856
rect 15059 1853 15071 1887
rect 15013 1847 15071 1853
rect 15105 1887 15163 1893
rect 15105 1853 15117 1887
rect 15151 1886 15163 1887
rect 15151 1858 15240 1886
rect 15151 1853 15163 1858
rect 15105 1847 15163 1853
rect 14093 1819 14151 1825
rect 14093 1816 14105 1819
rect 13280 1788 14105 1816
rect 9456 1720 11560 1748
rect 9456 1708 9462 1720
rect 11974 1708 11980 1760
rect 12032 1748 12038 1760
rect 12161 1751 12219 1757
rect 12161 1748 12173 1751
rect 12032 1720 12173 1748
rect 12032 1708 12038 1720
rect 12161 1717 12173 1720
rect 12207 1717 12219 1751
rect 12161 1711 12219 1717
rect 12437 1751 12495 1757
rect 12437 1717 12449 1751
rect 12483 1748 12495 1751
rect 13280 1748 13308 1788
rect 14093 1785 14105 1788
rect 14139 1785 14151 1819
rect 14093 1779 14151 1785
rect 12483 1720 13308 1748
rect 12483 1717 12495 1720
rect 12437 1711 12495 1717
rect 13354 1708 13360 1760
rect 13412 1708 13418 1760
rect 13722 1708 13728 1760
rect 13780 1748 13786 1760
rect 13909 1751 13967 1757
rect 13909 1748 13921 1751
rect 13780 1720 13921 1748
rect 13780 1708 13786 1720
rect 13909 1717 13921 1720
rect 13955 1748 13967 1751
rect 14660 1748 14688 1847
rect 15212 1748 15240 1858
rect 16942 1844 16948 1896
rect 17000 1844 17006 1896
rect 17052 1884 17080 1912
rect 19150 1884 19156 1896
rect 17052 1856 19156 1884
rect 19150 1844 19156 1856
rect 19208 1884 19214 1896
rect 19628 1884 19656 1992
rect 20070 1980 20076 1992
rect 20128 1980 20134 2032
rect 20438 2020 20444 2032
rect 20272 1992 20444 2020
rect 20272 1952 20300 1992
rect 20438 1980 20444 1992
rect 20496 1980 20502 2032
rect 19812 1924 20300 1952
rect 19208 1856 19656 1884
rect 19208 1844 19214 1856
rect 19702 1844 19708 1896
rect 19760 1844 19766 1896
rect 19812 1893 19840 1924
rect 19797 1887 19855 1893
rect 19797 1853 19809 1887
rect 19843 1853 19855 1887
rect 19797 1847 19855 1853
rect 19889 1887 19947 1893
rect 19889 1853 19901 1887
rect 19935 1853 19947 1887
rect 19889 1847 19947 1853
rect 15562 1825 15568 1828
rect 15556 1779 15568 1825
rect 15562 1776 15568 1779
rect 15620 1776 15626 1828
rect 17396 1819 17454 1825
rect 17396 1785 17408 1819
rect 17442 1816 17454 1819
rect 17678 1816 17684 1828
rect 17442 1788 17684 1816
rect 17442 1785 17454 1788
rect 17396 1779 17454 1785
rect 17678 1776 17684 1788
rect 17736 1776 17742 1828
rect 17954 1776 17960 1828
rect 18012 1816 18018 1828
rect 18693 1819 18751 1825
rect 18693 1816 18705 1819
rect 18012 1788 18705 1816
rect 18012 1776 18018 1788
rect 18693 1785 18705 1788
rect 18739 1785 18751 1819
rect 18693 1779 18751 1785
rect 18782 1776 18788 1828
rect 18840 1816 18846 1828
rect 19812 1816 19840 1847
rect 18840 1788 19840 1816
rect 19904 1816 19932 1847
rect 20070 1844 20076 1896
rect 20128 1844 20134 1896
rect 20346 1844 20352 1896
rect 20404 1844 20410 1896
rect 20438 1844 20444 1896
rect 20496 1844 20502 1896
rect 22756 1893 22784 2060
rect 24210 2048 24216 2060
rect 24268 2048 24274 2100
rect 24486 2088 24492 2100
rect 24320 2060 24492 2088
rect 24026 2020 24032 2032
rect 23032 1992 24032 2020
rect 20625 1887 20683 1893
rect 20625 1853 20637 1887
rect 20671 1884 20683 1887
rect 20809 1887 20867 1893
rect 20809 1884 20821 1887
rect 20671 1856 20821 1884
rect 20671 1853 20683 1856
rect 20625 1847 20683 1853
rect 20809 1853 20821 1856
rect 20855 1853 20867 1887
rect 20809 1847 20867 1853
rect 21361 1887 21419 1893
rect 21361 1853 21373 1887
rect 21407 1853 21419 1887
rect 21361 1847 21419 1853
rect 22741 1887 22799 1893
rect 22741 1853 22753 1887
rect 22787 1853 22799 1887
rect 22741 1847 22799 1853
rect 20533 1819 20591 1825
rect 20533 1816 20545 1819
rect 19904 1788 20545 1816
rect 18840 1776 18846 1788
rect 20533 1785 20545 1788
rect 20579 1785 20591 1819
rect 21376 1816 21404 1847
rect 22830 1844 22836 1896
rect 22888 1844 22894 1896
rect 23032 1893 23060 1992
rect 24026 1980 24032 1992
rect 24084 1980 24090 2032
rect 24320 2020 24348 2060
rect 24486 2048 24492 2060
rect 24544 2088 24550 2100
rect 24544 2060 25360 2088
rect 24544 2048 24550 2060
rect 25332 2029 25360 2060
rect 25682 2048 25688 2100
rect 25740 2048 25746 2100
rect 26142 2048 26148 2100
rect 26200 2088 26206 2100
rect 26200 2060 27384 2088
rect 26200 2048 26206 2060
rect 24127 1992 24348 2020
rect 25317 2023 25375 2029
rect 23750 1912 23756 1964
rect 23808 1952 23814 1964
rect 24127 1952 24155 1992
rect 25317 1989 25329 2023
rect 25363 2020 25375 2023
rect 25961 2023 26019 2029
rect 25961 2020 25973 2023
rect 25363 1992 25973 2020
rect 25363 1989 25375 1992
rect 25317 1983 25375 1989
rect 25961 1989 25973 1992
rect 26007 1989 26019 2023
rect 27356 2020 27384 2060
rect 27614 2048 27620 2100
rect 27672 2088 27678 2100
rect 27801 2091 27859 2097
rect 27801 2088 27813 2091
rect 27672 2060 27813 2088
rect 27672 2048 27678 2060
rect 27801 2057 27813 2060
rect 27847 2057 27859 2091
rect 27801 2051 27859 2057
rect 28902 2020 28908 2032
rect 27356 1992 28908 2020
rect 25961 1983 26019 1989
rect 28902 1980 28908 1992
rect 28960 1980 28966 2032
rect 23808 1924 24155 1952
rect 23808 1912 23814 1924
rect 25222 1912 25228 1964
rect 25280 1912 25286 1964
rect 26418 1912 26424 1964
rect 26476 1912 26482 1964
rect 23017 1887 23075 1893
rect 23017 1853 23029 1887
rect 23063 1853 23075 1887
rect 23017 1847 23075 1853
rect 23106 1844 23112 1896
rect 23164 1844 23170 1896
rect 23198 1844 23204 1896
rect 23256 1844 23262 1896
rect 24670 1884 24676 1896
rect 23308 1856 24676 1884
rect 20533 1779 20591 1785
rect 20640 1788 21404 1816
rect 20640 1760 20668 1788
rect 22370 1776 22376 1828
rect 22428 1816 22434 1828
rect 22848 1816 22876 1844
rect 23308 1816 23336 1856
rect 24670 1844 24676 1856
rect 24728 1844 24734 1896
rect 25130 1844 25136 1896
rect 25188 1884 25194 1896
rect 26510 1884 26516 1896
rect 25188 1856 26516 1884
rect 25188 1844 25194 1856
rect 25700 1825 25728 1856
rect 26510 1844 26516 1856
rect 26568 1844 26574 1896
rect 28074 1844 28080 1896
rect 28132 1844 28138 1896
rect 22428 1788 22784 1816
rect 22848 1788 23336 1816
rect 23477 1819 23535 1825
rect 22428 1776 22434 1788
rect 15470 1748 15476 1760
rect 13955 1720 15476 1748
rect 13955 1717 13967 1720
rect 13909 1711 13967 1717
rect 15470 1708 15476 1720
rect 15528 1708 15534 1760
rect 19426 1708 19432 1760
rect 19484 1708 19490 1760
rect 19610 1708 19616 1760
rect 19668 1748 19674 1760
rect 20257 1751 20315 1757
rect 20257 1748 20269 1751
rect 19668 1720 20269 1748
rect 19668 1708 19674 1720
rect 20257 1717 20269 1720
rect 20303 1717 20315 1751
rect 20257 1711 20315 1717
rect 20622 1708 20628 1760
rect 20680 1708 20686 1760
rect 22646 1708 22652 1760
rect 22704 1708 22710 1760
rect 22756 1748 22784 1788
rect 23477 1785 23489 1819
rect 23523 1816 23535 1819
rect 24958 1819 25016 1825
rect 24958 1816 24970 1819
rect 23523 1788 24970 1816
rect 23523 1785 23535 1788
rect 23477 1779 23535 1785
rect 24958 1785 24970 1788
rect 25004 1785 25016 1819
rect 24958 1779 25016 1785
rect 25685 1819 25743 1825
rect 25685 1785 25697 1819
rect 25731 1785 25743 1819
rect 25685 1779 25743 1785
rect 25774 1776 25780 1828
rect 25832 1816 25838 1828
rect 26329 1819 26387 1825
rect 26329 1816 26341 1819
rect 25832 1788 26341 1816
rect 25832 1776 25838 1788
rect 26329 1785 26341 1788
rect 26375 1785 26387 1819
rect 26329 1779 26387 1785
rect 26688 1819 26746 1825
rect 26688 1785 26700 1819
rect 26734 1816 26746 1819
rect 26970 1816 26976 1828
rect 26734 1788 26976 1816
rect 26734 1785 26746 1788
rect 26688 1779 26746 1785
rect 26970 1776 26976 1788
rect 27028 1776 27034 1828
rect 23198 1748 23204 1760
rect 22756 1720 23204 1748
rect 23198 1708 23204 1720
rect 23256 1748 23262 1760
rect 23845 1751 23903 1757
rect 23845 1748 23857 1751
rect 23256 1720 23857 1748
rect 23256 1708 23262 1720
rect 23845 1717 23857 1720
rect 23891 1748 23903 1751
rect 24854 1748 24860 1760
rect 23891 1720 24860 1748
rect 23891 1717 23903 1720
rect 23845 1711 23903 1717
rect 24854 1708 24860 1720
rect 24912 1708 24918 1760
rect 25866 1708 25872 1760
rect 25924 1708 25930 1760
rect 26129 1751 26187 1757
rect 26129 1717 26141 1751
rect 26175 1748 26187 1751
rect 26418 1748 26424 1760
rect 26175 1720 26424 1748
rect 26175 1717 26187 1720
rect 26129 1711 26187 1717
rect 26418 1708 26424 1720
rect 26476 1748 26482 1760
rect 26786 1748 26792 1760
rect 26476 1720 26792 1748
rect 26476 1708 26482 1720
rect 26786 1708 26792 1720
rect 26844 1708 26850 1760
rect 27982 1708 27988 1760
rect 28040 1708 28046 1760
rect 552 1658 31648 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 12096 1658
rect 12148 1606 12160 1658
rect 12212 1606 12224 1658
rect 12276 1606 12288 1658
rect 12340 1606 12352 1658
rect 12404 1606 19870 1658
rect 19922 1606 19934 1658
rect 19986 1606 19998 1658
rect 20050 1606 20062 1658
rect 20114 1606 20126 1658
rect 20178 1606 27644 1658
rect 27696 1606 27708 1658
rect 27760 1606 27772 1658
rect 27824 1606 27836 1658
rect 27888 1606 27900 1658
rect 27952 1606 31648 1658
rect 552 1584 31648 1606
rect 5629 1547 5687 1553
rect 5629 1513 5641 1547
rect 5675 1544 5687 1547
rect 6822 1544 6828 1556
rect 5675 1516 6828 1544
rect 5675 1513 5687 1516
rect 5629 1507 5687 1513
rect 6822 1504 6828 1516
rect 6880 1504 6886 1556
rect 7561 1547 7619 1553
rect 7561 1513 7573 1547
rect 7607 1544 7619 1547
rect 7929 1547 7987 1553
rect 7929 1544 7941 1547
rect 7607 1516 7941 1544
rect 7607 1513 7619 1516
rect 7561 1507 7619 1513
rect 7929 1513 7941 1516
rect 7975 1544 7987 1547
rect 8294 1544 8300 1556
rect 7975 1516 8300 1544
rect 7975 1513 7987 1516
rect 7929 1507 7987 1513
rect 8294 1504 8300 1516
rect 8352 1504 8358 1556
rect 8846 1504 8852 1556
rect 8904 1504 8910 1556
rect 10594 1544 10600 1556
rect 8956 1516 10600 1544
rect 4516 1479 4574 1485
rect 4516 1445 4528 1479
rect 4562 1476 4574 1479
rect 4706 1476 4712 1488
rect 4562 1448 4712 1476
rect 4562 1445 4574 1448
rect 4516 1439 4574 1445
rect 4706 1436 4712 1448
rect 4764 1436 4770 1488
rect 6448 1479 6506 1485
rect 6448 1445 6460 1479
rect 6494 1476 6506 1479
rect 7006 1476 7012 1488
rect 6494 1448 7012 1476
rect 6494 1445 6506 1448
rect 6448 1439 6506 1445
rect 7006 1436 7012 1448
rect 7064 1436 7070 1488
rect 8018 1436 8024 1488
rect 8076 1436 8082 1488
rect 8662 1436 8668 1488
rect 8720 1436 8726 1488
rect 4246 1368 4252 1420
rect 4304 1368 4310 1420
rect 6086 1368 6092 1420
rect 6144 1368 6150 1420
rect 7837 1411 7895 1417
rect 7837 1377 7849 1411
rect 7883 1408 7895 1411
rect 8386 1408 8392 1420
rect 7883 1380 8392 1408
rect 7883 1377 7895 1380
rect 7837 1371 7895 1377
rect 8386 1368 8392 1380
rect 8444 1408 8450 1420
rect 8846 1408 8852 1420
rect 8444 1380 8852 1408
rect 8444 1368 8450 1380
rect 8846 1368 8852 1380
rect 8904 1368 8910 1420
rect 5810 1300 5816 1352
rect 5868 1300 5874 1352
rect 6178 1300 6184 1352
rect 6236 1300 6242 1352
rect 7190 1300 7196 1352
rect 7248 1340 7254 1352
rect 8297 1343 8355 1349
rect 8297 1340 8309 1343
rect 7248 1312 8309 1340
rect 7248 1300 7254 1312
rect 8297 1309 8309 1312
rect 8343 1309 8355 1343
rect 8297 1303 8355 1309
rect 5442 1232 5448 1284
rect 5500 1272 5506 1284
rect 5905 1275 5963 1281
rect 5905 1272 5917 1275
rect 5500 1244 5917 1272
rect 5500 1232 5506 1244
rect 5905 1241 5917 1244
rect 5951 1241 5963 1275
rect 5905 1235 5963 1241
rect 7466 1232 7472 1284
rect 7524 1272 7530 1284
rect 8205 1275 8263 1281
rect 8205 1272 8217 1275
rect 7524 1244 8217 1272
rect 7524 1232 7530 1244
rect 8205 1241 8217 1244
rect 8251 1272 8263 1275
rect 8956 1272 8984 1516
rect 10594 1504 10600 1516
rect 10652 1544 10658 1556
rect 10689 1547 10747 1553
rect 10689 1544 10701 1547
rect 10652 1516 10701 1544
rect 10652 1504 10658 1516
rect 10689 1513 10701 1516
rect 10735 1513 10747 1547
rect 10689 1507 10747 1513
rect 12529 1547 12587 1553
rect 12529 1513 12541 1547
rect 12575 1544 12587 1547
rect 12575 1516 13492 1544
rect 12575 1513 12587 1516
rect 12529 1507 12587 1513
rect 9214 1436 9220 1488
rect 9272 1476 9278 1488
rect 9554 1479 9612 1485
rect 9554 1476 9566 1479
rect 9272 1448 9566 1476
rect 9272 1436 9278 1448
rect 9554 1445 9566 1448
rect 9600 1445 9612 1479
rect 9554 1439 9612 1445
rect 12069 1479 12127 1485
rect 12069 1445 12081 1479
rect 12115 1476 12127 1479
rect 12618 1476 12624 1488
rect 12115 1448 12624 1476
rect 12115 1445 12127 1448
rect 12069 1439 12127 1445
rect 12618 1436 12624 1448
rect 12676 1436 12682 1488
rect 12888 1479 12946 1485
rect 12888 1445 12900 1479
rect 12934 1476 12946 1479
rect 13354 1476 13360 1488
rect 12934 1448 13360 1476
rect 12934 1445 12946 1448
rect 12888 1439 12946 1445
rect 13354 1436 13360 1448
rect 13412 1436 13418 1488
rect 13464 1476 13492 1516
rect 13998 1504 14004 1556
rect 14056 1504 14062 1556
rect 15470 1504 15476 1556
rect 15528 1504 15534 1556
rect 15562 1504 15568 1556
rect 15620 1504 15626 1556
rect 17218 1504 17224 1556
rect 17276 1544 17282 1556
rect 17589 1547 17647 1553
rect 17589 1544 17601 1547
rect 17276 1516 17601 1544
rect 17276 1504 17282 1516
rect 17589 1513 17601 1516
rect 17635 1513 17647 1547
rect 17589 1507 17647 1513
rect 17678 1504 17684 1556
rect 17736 1504 17742 1556
rect 19058 1504 19064 1556
rect 19116 1544 19122 1556
rect 19153 1547 19211 1553
rect 19153 1544 19165 1547
rect 19116 1516 19165 1544
rect 19116 1504 19122 1516
rect 19153 1513 19165 1516
rect 19199 1513 19211 1547
rect 19153 1507 19211 1513
rect 19702 1504 19708 1556
rect 19760 1544 19766 1556
rect 20622 1544 20628 1556
rect 19760 1516 20628 1544
rect 19760 1504 19766 1516
rect 20622 1504 20628 1516
rect 20680 1544 20686 1556
rect 20993 1547 21051 1553
rect 20993 1544 21005 1547
rect 20680 1516 21005 1544
rect 20680 1504 20686 1516
rect 20993 1513 21005 1516
rect 21039 1513 21051 1547
rect 20993 1507 21051 1513
rect 23014 1504 23020 1556
rect 23072 1504 23078 1556
rect 23201 1547 23259 1553
rect 23201 1513 23213 1547
rect 23247 1513 23259 1547
rect 23201 1507 23259 1513
rect 16482 1485 16488 1488
rect 14338 1479 14396 1485
rect 14338 1476 14350 1479
rect 13464 1448 14350 1476
rect 14338 1445 14350 1448
rect 14384 1445 14396 1479
rect 16476 1476 16488 1485
rect 16443 1448 16488 1476
rect 14338 1439 14396 1445
rect 16476 1439 16488 1448
rect 16482 1436 16488 1439
rect 16540 1436 16546 1488
rect 17862 1436 17868 1488
rect 17920 1476 17926 1488
rect 17920 1448 18184 1476
rect 17920 1436 17926 1448
rect 9030 1368 9036 1420
rect 9088 1368 9094 1420
rect 11974 1368 11980 1420
rect 12032 1408 12038 1420
rect 12636 1408 12664 1436
rect 13722 1408 13728 1420
rect 12032 1380 12434 1408
rect 12636 1380 13728 1408
rect 12032 1368 12038 1380
rect 9125 1343 9183 1349
rect 9125 1309 9137 1343
rect 9171 1340 9183 1343
rect 9309 1343 9367 1349
rect 9309 1340 9321 1343
rect 9171 1312 9321 1340
rect 9171 1309 9183 1312
rect 9125 1303 9183 1309
rect 9309 1309 9321 1312
rect 9355 1309 9367 1343
rect 12406 1340 12434 1380
rect 13722 1368 13728 1380
rect 13780 1368 13786 1420
rect 14090 1368 14096 1420
rect 14148 1368 14154 1420
rect 15746 1368 15752 1420
rect 15804 1368 15810 1420
rect 16209 1411 16267 1417
rect 16209 1377 16221 1411
rect 16255 1408 16267 1411
rect 16298 1408 16304 1420
rect 16255 1380 16304 1408
rect 16255 1377 16267 1380
rect 16209 1371 16267 1377
rect 16298 1368 16304 1380
rect 16356 1368 16362 1420
rect 17954 1368 17960 1420
rect 18012 1368 18018 1420
rect 18156 1417 18184 1448
rect 19426 1436 19432 1488
rect 19484 1476 19490 1488
rect 19858 1479 19916 1485
rect 19858 1476 19870 1479
rect 19484 1448 19870 1476
rect 19484 1436 19490 1448
rect 19858 1445 19870 1448
rect 19904 1445 19916 1479
rect 23216 1476 23244 1507
rect 24118 1504 24124 1556
rect 24176 1544 24182 1556
rect 24673 1547 24731 1553
rect 24673 1544 24685 1547
rect 24176 1516 24685 1544
rect 24176 1504 24182 1516
rect 24673 1513 24685 1516
rect 24719 1513 24731 1547
rect 24673 1507 24731 1513
rect 24857 1547 24915 1553
rect 24857 1513 24869 1547
rect 24903 1544 24915 1547
rect 25774 1544 25780 1556
rect 24903 1516 25780 1544
rect 24903 1513 24915 1516
rect 24857 1507 24915 1513
rect 25774 1504 25780 1516
rect 25832 1504 25838 1556
rect 26789 1547 26847 1553
rect 26789 1513 26801 1547
rect 26835 1544 26847 1547
rect 26878 1544 26884 1556
rect 26835 1516 26884 1544
rect 26835 1513 26847 1516
rect 26789 1507 26847 1513
rect 23538 1479 23596 1485
rect 23538 1476 23550 1479
rect 23216 1448 23550 1476
rect 19858 1439 19916 1445
rect 23538 1445 23550 1448
rect 23584 1445 23596 1479
rect 23538 1439 23596 1445
rect 25866 1436 25872 1488
rect 25924 1476 25930 1488
rect 25970 1479 26028 1485
rect 25970 1476 25982 1479
rect 25924 1448 25982 1476
rect 25924 1436 25930 1448
rect 25970 1445 25982 1448
rect 26016 1445 26028 1479
rect 25970 1439 26028 1445
rect 18049 1411 18107 1417
rect 18049 1377 18061 1411
rect 18095 1377 18107 1411
rect 18049 1371 18107 1377
rect 18141 1411 18199 1417
rect 18141 1377 18153 1411
rect 18187 1377 18199 1411
rect 18141 1371 18199 1377
rect 18325 1411 18383 1417
rect 18325 1377 18337 1411
rect 18371 1408 18383 1411
rect 19150 1408 19156 1420
rect 18371 1380 19156 1408
rect 18371 1377 18383 1380
rect 18325 1371 18383 1377
rect 12621 1343 12679 1349
rect 12621 1340 12633 1343
rect 12406 1312 12633 1340
rect 9309 1303 9367 1309
rect 12621 1309 12633 1312
rect 12667 1309 12679 1343
rect 12621 1303 12679 1309
rect 15933 1343 15991 1349
rect 15933 1309 15945 1343
rect 15979 1340 15991 1343
rect 18064 1340 18092 1371
rect 19150 1368 19156 1380
rect 19208 1368 19214 1420
rect 19610 1368 19616 1420
rect 19668 1368 19674 1420
rect 22646 1368 22652 1420
rect 22704 1408 22710 1420
rect 23293 1411 23351 1417
rect 23293 1408 23305 1411
rect 22704 1380 23305 1408
rect 22704 1368 22710 1380
rect 23293 1377 23305 1380
rect 23339 1377 23351 1411
rect 23293 1371 23351 1377
rect 24026 1368 24032 1420
rect 24084 1408 24090 1420
rect 26804 1408 26832 1507
rect 26878 1504 26884 1516
rect 26936 1504 26942 1556
rect 26970 1504 26976 1556
rect 27028 1504 27034 1556
rect 27338 1504 27344 1556
rect 27396 1544 27402 1556
rect 27396 1516 28120 1544
rect 27396 1504 27402 1516
rect 27982 1476 27988 1488
rect 27724 1448 27988 1476
rect 27724 1408 27752 1448
rect 27982 1436 27988 1448
rect 28040 1436 28046 1488
rect 24084 1380 26832 1408
rect 27632 1380 27752 1408
rect 27792 1411 27850 1417
rect 24084 1368 24090 1380
rect 18690 1340 18696 1352
rect 15979 1312 16252 1340
rect 18064 1312 18696 1340
rect 15979 1309 15991 1312
rect 15933 1303 15991 1309
rect 8251 1244 8984 1272
rect 8251 1241 8263 1244
rect 8205 1235 8263 1241
rect 11790 1232 11796 1284
rect 11848 1272 11854 1284
rect 12345 1275 12403 1281
rect 12345 1272 12357 1275
rect 11848 1244 12357 1272
rect 11848 1232 11854 1244
rect 12345 1241 12357 1244
rect 12391 1241 12403 1275
rect 12345 1235 12403 1241
rect 5994 1164 6000 1216
rect 6052 1204 6058 1216
rect 7653 1207 7711 1213
rect 7653 1204 7665 1207
rect 6052 1176 7665 1204
rect 6052 1164 6058 1176
rect 7653 1173 7665 1176
rect 7699 1173 7711 1207
rect 7653 1167 7711 1173
rect 8570 1164 8576 1216
rect 8628 1204 8634 1216
rect 8665 1207 8723 1213
rect 8665 1204 8677 1207
rect 8628 1176 8677 1204
rect 8628 1164 8634 1176
rect 8665 1173 8677 1176
rect 8711 1173 8723 1207
rect 16224 1204 16252 1312
rect 18690 1300 18696 1312
rect 18748 1340 18754 1352
rect 18785 1343 18843 1349
rect 18785 1340 18797 1343
rect 18748 1312 18797 1340
rect 18748 1300 18754 1312
rect 18785 1309 18797 1312
rect 18831 1309 18843 1343
rect 18785 1303 18843 1309
rect 26234 1300 26240 1352
rect 26292 1300 26298 1352
rect 26418 1300 26424 1352
rect 26476 1300 26482 1352
rect 27525 1343 27583 1349
rect 27525 1309 27537 1343
rect 27571 1340 27583 1343
rect 27632 1340 27660 1380
rect 27792 1377 27804 1411
rect 27838 1408 27850 1411
rect 28092 1408 28120 1516
rect 28902 1504 28908 1556
rect 28960 1504 28966 1556
rect 27838 1380 28120 1408
rect 27838 1377 27850 1380
rect 27792 1371 27850 1377
rect 27571 1312 27660 1340
rect 27571 1309 27583 1312
rect 27525 1303 27583 1309
rect 22649 1275 22707 1281
rect 22649 1241 22661 1275
rect 22695 1272 22707 1275
rect 23106 1272 23112 1284
rect 22695 1244 23112 1272
rect 22695 1241 22707 1244
rect 22649 1235 22707 1241
rect 23106 1232 23112 1244
rect 23164 1232 23170 1284
rect 16574 1204 16580 1216
rect 16224 1176 16580 1204
rect 8665 1167 8723 1173
rect 16574 1164 16580 1176
rect 16632 1164 16638 1216
rect 19150 1164 19156 1216
rect 19208 1164 19214 1216
rect 19337 1207 19395 1213
rect 19337 1173 19349 1207
rect 19383 1204 19395 1207
rect 19610 1204 19616 1216
rect 19383 1176 19616 1204
rect 19383 1173 19395 1176
rect 19337 1167 19395 1173
rect 19610 1164 19616 1176
rect 19668 1164 19674 1216
rect 23017 1207 23075 1213
rect 23017 1173 23029 1207
rect 23063 1204 23075 1207
rect 23934 1204 23940 1216
rect 23063 1176 23940 1204
rect 23063 1173 23075 1176
rect 23017 1167 23075 1173
rect 23934 1164 23940 1176
rect 23992 1164 23998 1216
rect 26789 1207 26847 1213
rect 26789 1173 26801 1207
rect 26835 1204 26847 1207
rect 27430 1204 27436 1216
rect 26835 1176 27436 1204
rect 26835 1173 26847 1176
rect 26789 1167 26847 1173
rect 27430 1164 27436 1176
rect 27488 1164 27494 1216
rect 552 1114 31648 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 11436 1114
rect 11488 1062 11500 1114
rect 11552 1062 11564 1114
rect 11616 1062 11628 1114
rect 11680 1062 11692 1114
rect 11744 1062 19210 1114
rect 19262 1062 19274 1114
rect 19326 1062 19338 1114
rect 19390 1062 19402 1114
rect 19454 1062 19466 1114
rect 19518 1062 26984 1114
rect 27036 1062 27048 1114
rect 27100 1062 27112 1114
rect 27164 1062 27176 1114
rect 27228 1062 27240 1114
rect 27292 1062 31648 1114
rect 552 1040 31648 1062
rect 6914 960 6920 1012
rect 6972 960 6978 1012
rect 7009 1003 7067 1009
rect 7009 969 7021 1003
rect 7055 1000 7067 1003
rect 7190 1000 7196 1012
rect 7055 972 7196 1000
rect 7055 969 7067 972
rect 7009 963 7067 969
rect 7190 960 7196 972
rect 7248 960 7254 1012
rect 7377 1003 7435 1009
rect 7377 969 7389 1003
rect 7423 1000 7435 1003
rect 8018 1000 8024 1012
rect 7423 972 8024 1000
rect 7423 969 7435 972
rect 7377 963 7435 969
rect 8018 960 8024 972
rect 8076 960 8082 1012
rect 8662 960 8668 1012
rect 8720 1000 8726 1012
rect 8849 1003 8907 1009
rect 8849 1000 8861 1003
rect 8720 972 8861 1000
rect 8720 960 8726 972
rect 8849 969 8861 972
rect 8895 969 8907 1003
rect 8849 963 8907 969
rect 9033 1003 9091 1009
rect 9033 969 9045 1003
rect 9079 1000 9091 1003
rect 9766 1000 9772 1012
rect 9079 972 9772 1000
rect 9079 969 9091 972
rect 9033 963 9091 969
rect 9766 960 9772 972
rect 9824 960 9830 1012
rect 18690 960 18696 1012
rect 18748 960 18754 1012
rect 18874 960 18880 1012
rect 18932 960 18938 1012
rect 8036 932 8064 960
rect 8036 904 8708 932
rect 5810 824 5816 876
rect 5868 864 5874 876
rect 6825 867 6883 873
rect 6825 864 6837 867
rect 5868 836 6837 864
rect 5868 824 5874 836
rect 6825 833 6837 836
rect 6871 864 6883 867
rect 8570 864 8576 876
rect 6871 836 8576 864
rect 6871 833 6883 836
rect 6825 827 6883 833
rect 8570 824 8576 836
rect 8628 824 8634 876
rect 7098 756 7104 808
rect 7156 756 7162 808
rect 8386 796 8392 808
rect 7392 768 8392 796
rect 7392 737 7420 768
rect 8386 756 8392 768
rect 8444 756 8450 808
rect 8680 805 8708 904
rect 8665 799 8723 805
rect 8665 765 8677 799
rect 8711 765 8723 799
rect 8665 759 8723 765
rect 8941 799 8999 805
rect 8941 765 8953 799
rect 8987 796 8999 799
rect 9030 796 9036 808
rect 8987 768 9036 796
rect 8987 765 8999 768
rect 8941 759 8999 765
rect 9030 756 9036 768
rect 9088 756 9094 808
rect 18322 756 18328 808
rect 18380 756 18386 808
rect 19610 805 19616 808
rect 18417 799 18475 805
rect 18417 765 18429 799
rect 18463 796 18475 799
rect 19337 799 19395 805
rect 19337 796 19349 799
rect 18463 768 19349 796
rect 18463 765 18475 768
rect 18417 759 18475 765
rect 19337 765 19349 768
rect 19383 765 19395 799
rect 19604 796 19616 805
rect 19571 768 19616 796
rect 19337 759 19395 765
rect 19604 759 19616 768
rect 19610 756 19616 759
rect 19668 756 19674 808
rect 7361 731 7420 737
rect 7361 697 7373 731
rect 7407 700 7420 731
rect 7407 697 7419 700
rect 7361 691 7419 697
rect 7466 688 7472 740
rect 7524 728 7530 740
rect 18874 737 18880 740
rect 7561 731 7619 737
rect 7561 728 7573 731
rect 7524 700 7573 728
rect 7524 688 7530 700
rect 7561 697 7573 700
rect 7607 728 7619 731
rect 8481 731 8539 737
rect 8481 728 8493 731
rect 7607 700 8493 728
rect 7607 697 7619 700
rect 7561 691 7619 697
rect 8481 697 8493 700
rect 8527 697 8539 731
rect 8481 691 8539 697
rect 18861 731 18880 737
rect 18861 697 18873 731
rect 18861 691 18880 697
rect 18874 688 18880 691
rect 18932 688 18938 740
rect 18966 688 18972 740
rect 19024 728 19030 740
rect 19061 731 19119 737
rect 19061 728 19073 731
rect 19024 700 19073 728
rect 19024 688 19030 700
rect 19061 697 19073 700
rect 19107 697 19119 731
rect 19061 691 19119 697
rect 19076 660 19104 691
rect 20717 663 20775 669
rect 20717 660 20729 663
rect 19076 632 20729 660
rect 20717 629 20729 632
rect 20763 629 20775 663
rect 20717 623 20775 629
rect 552 570 31648 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 12096 570
rect 12148 518 12160 570
rect 12212 518 12224 570
rect 12276 518 12288 570
rect 12340 518 12352 570
rect 12404 518 19870 570
rect 19922 518 19934 570
rect 19986 518 19998 570
rect 20050 518 20062 570
rect 20114 518 20126 570
rect 20178 518 27644 570
rect 27696 518 27708 570
rect 27760 518 27772 570
rect 27824 518 27836 570
rect 27888 518 27900 570
rect 27952 518 31648 570
rect 552 496 31648 518
<< via1 >>
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 11436 21734 11488 21786
rect 11500 21734 11552 21786
rect 11564 21734 11616 21786
rect 11628 21734 11680 21786
rect 11692 21734 11744 21786
rect 19210 21734 19262 21786
rect 19274 21734 19326 21786
rect 19338 21734 19390 21786
rect 19402 21734 19454 21786
rect 19466 21734 19518 21786
rect 26984 21734 27036 21786
rect 27048 21734 27100 21786
rect 27112 21734 27164 21786
rect 27176 21734 27228 21786
rect 27240 21734 27292 21786
rect 6092 21675 6144 21684
rect 6092 21641 6101 21675
rect 6101 21641 6135 21675
rect 6135 21641 6144 21675
rect 6092 21632 6144 21641
rect 8024 21675 8076 21684
rect 8024 21641 8033 21675
rect 8033 21641 8067 21675
rect 8067 21641 8076 21675
rect 8024 21632 8076 21641
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 8668 21675 8720 21684
rect 8668 21641 8677 21675
rect 8677 21641 8711 21675
rect 8711 21641 8720 21675
rect 8668 21632 8720 21641
rect 11796 21632 11848 21684
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12992 21675 13044 21684
rect 12992 21641 13001 21675
rect 13001 21641 13035 21675
rect 13035 21641 13044 21675
rect 12992 21632 13044 21641
rect 18788 21632 18840 21684
rect 29276 21632 29328 21684
rect 1400 21428 1452 21480
rect 2964 21471 3016 21480
rect 2964 21437 2973 21471
rect 2973 21437 3007 21471
rect 3007 21437 3016 21471
rect 2964 21428 3016 21437
rect 4160 21428 4212 21480
rect 5356 21428 5408 21480
rect 7196 21496 7248 21548
rect 13912 21496 13964 21548
rect 23664 21496 23716 21548
rect 3148 21360 3200 21412
rect 6920 21428 6972 21480
rect 12808 21428 12860 21480
rect 19616 21428 19668 21480
rect 20628 21428 20680 21480
rect 7012 21403 7064 21412
rect 7012 21369 7021 21403
rect 7021 21369 7055 21403
rect 7055 21369 7064 21403
rect 7012 21360 7064 21369
rect 14648 21360 14700 21412
rect 17868 21403 17920 21412
rect 17868 21369 17877 21403
rect 17877 21369 17911 21403
rect 17911 21369 17920 21403
rect 17868 21360 17920 21369
rect 18052 21403 18104 21412
rect 18052 21369 18077 21403
rect 18077 21369 18104 21403
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 23848 21471 23900 21480
rect 23848 21437 23857 21471
rect 23857 21437 23891 21471
rect 23891 21437 23900 21471
rect 23848 21428 23900 21437
rect 24400 21471 24452 21480
rect 24400 21437 24409 21471
rect 24409 21437 24443 21471
rect 24443 21437 24452 21471
rect 24400 21428 24452 21437
rect 26424 21471 26476 21480
rect 26424 21437 26433 21471
rect 26433 21437 26467 21471
rect 26467 21437 26476 21471
rect 26424 21428 26476 21437
rect 26700 21471 26752 21480
rect 26700 21437 26709 21471
rect 26709 21437 26743 21471
rect 26743 21437 26752 21471
rect 26700 21428 26752 21437
rect 27344 21428 27396 21480
rect 27712 21471 27764 21480
rect 27712 21437 27721 21471
rect 27721 21437 27755 21471
rect 27755 21437 27764 21471
rect 27712 21428 27764 21437
rect 28264 21471 28316 21480
rect 28264 21437 28273 21471
rect 28273 21437 28307 21471
rect 28307 21437 28316 21471
rect 28264 21428 28316 21437
rect 29000 21471 29052 21480
rect 29000 21437 29009 21471
rect 29009 21437 29043 21471
rect 29043 21437 29052 21471
rect 29000 21428 29052 21437
rect 18052 21360 18104 21369
rect 24676 21360 24728 21412
rect 25136 21360 25188 21412
rect 1952 21292 2004 21344
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 5264 21335 5316 21344
rect 5264 21301 5273 21335
rect 5273 21301 5307 21335
rect 5307 21301 5316 21335
rect 5264 21292 5316 21301
rect 6644 21335 6696 21344
rect 6644 21301 6653 21335
rect 6653 21301 6687 21335
rect 6687 21301 6696 21335
rect 6644 21292 6696 21301
rect 6828 21335 6880 21344
rect 6828 21301 6837 21335
rect 6837 21301 6871 21335
rect 6871 21301 6880 21335
rect 6828 21292 6880 21301
rect 12624 21292 12676 21344
rect 12992 21292 13044 21344
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 14004 21292 14056 21301
rect 16856 21292 16908 21344
rect 18236 21335 18288 21344
rect 18236 21301 18245 21335
rect 18245 21301 18279 21335
rect 18279 21301 18288 21335
rect 18236 21292 18288 21301
rect 21272 21292 21324 21344
rect 21824 21292 21876 21344
rect 22376 21335 22428 21344
rect 22376 21301 22385 21335
rect 22385 21301 22419 21335
rect 22419 21301 22428 21335
rect 22376 21292 22428 21301
rect 24032 21335 24084 21344
rect 24032 21301 24041 21335
rect 24041 21301 24075 21335
rect 24075 21301 24084 21335
rect 24032 21292 24084 21301
rect 24584 21335 24636 21344
rect 24584 21301 24593 21335
rect 24593 21301 24627 21335
rect 24627 21301 24636 21335
rect 24584 21292 24636 21301
rect 26056 21335 26108 21344
rect 26056 21301 26065 21335
rect 26065 21301 26099 21335
rect 26099 21301 26108 21335
rect 26056 21292 26108 21301
rect 27068 21292 27120 21344
rect 27344 21335 27396 21344
rect 27344 21301 27353 21335
rect 27353 21301 27387 21335
rect 27387 21301 27396 21335
rect 27344 21292 27396 21301
rect 30104 21292 30156 21344
rect 30380 21335 30432 21344
rect 30380 21301 30389 21335
rect 30389 21301 30423 21335
rect 30423 21301 30432 21335
rect 30380 21292 30432 21301
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 12096 21190 12148 21242
rect 12160 21190 12212 21242
rect 12224 21190 12276 21242
rect 12288 21190 12340 21242
rect 12352 21190 12404 21242
rect 19870 21190 19922 21242
rect 19934 21190 19986 21242
rect 19998 21190 20050 21242
rect 20062 21190 20114 21242
rect 20126 21190 20178 21242
rect 27644 21190 27696 21242
rect 27708 21190 27760 21242
rect 27772 21190 27824 21242
rect 27836 21190 27888 21242
rect 27900 21190 27952 21242
rect 2964 21088 3016 21140
rect 6828 21088 6880 21140
rect 7196 21131 7248 21140
rect 7196 21097 7205 21131
rect 7205 21097 7239 21131
rect 7239 21097 7248 21131
rect 7196 21088 7248 21097
rect 8116 21088 8168 21140
rect 6644 21020 6696 21072
rect 1952 20995 2004 21004
rect 1952 20961 1961 20995
rect 1961 20961 1995 20995
rect 1995 20961 2004 20995
rect 1952 20952 2004 20961
rect 2504 20952 2556 21004
rect 3516 20952 3568 21004
rect 4068 20952 4120 21004
rect 4160 20995 4212 21004
rect 4160 20961 4169 20995
rect 4169 20961 4203 20995
rect 4203 20961 4212 20995
rect 4160 20952 4212 20961
rect 4712 20995 4764 21004
rect 4712 20961 4721 20995
rect 4721 20961 4755 20995
rect 4755 20961 4764 20995
rect 4712 20952 4764 20961
rect 4896 20995 4948 21004
rect 4896 20961 4905 20995
rect 4905 20961 4939 20995
rect 4939 20961 4948 20995
rect 4896 20952 4948 20961
rect 5264 20952 5316 21004
rect 6920 20952 6972 21004
rect 8576 21131 8628 21140
rect 8576 21097 8585 21131
rect 8585 21097 8619 21131
rect 8619 21097 8628 21131
rect 8576 21088 8628 21097
rect 8944 21131 8996 21140
rect 8944 21097 8953 21131
rect 8953 21097 8987 21131
rect 8987 21097 8996 21131
rect 8944 21088 8996 21097
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 17868 21088 17920 21140
rect 18052 21088 18104 21140
rect 19524 21088 19576 21140
rect 22192 21088 22244 21140
rect 25136 21131 25188 21140
rect 25136 21097 25145 21131
rect 25145 21097 25179 21131
rect 25179 21097 25188 21131
rect 25136 21088 25188 21097
rect 27344 21088 27396 21140
rect 9404 20952 9456 21004
rect 9496 20995 9548 21004
rect 9496 20961 9505 20995
rect 9505 20961 9539 20995
rect 9539 20961 9548 20995
rect 9496 20952 9548 20961
rect 18236 21020 18288 21072
rect 9680 20952 9732 21004
rect 11244 20995 11296 21004
rect 11244 20961 11253 20995
rect 11253 20961 11287 20995
rect 11287 20961 11296 20995
rect 11244 20952 11296 20961
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 16856 20995 16908 21004
rect 16856 20961 16865 20995
rect 16865 20961 16899 20995
rect 16899 20961 16908 20995
rect 16856 20952 16908 20961
rect 17132 20995 17184 21004
rect 17132 20961 17166 20995
rect 17166 20961 17184 20995
rect 17132 20952 17184 20961
rect 18328 20952 18380 21004
rect 19064 20952 19116 21004
rect 8852 20884 8904 20936
rect 12900 20927 12952 20936
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 14832 20927 14884 20936
rect 14832 20893 14841 20927
rect 14841 20893 14875 20927
rect 14875 20893 14884 20927
rect 14832 20884 14884 20893
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 18696 20884 18748 20936
rect 3240 20816 3292 20868
rect 13636 20816 13688 20868
rect 17868 20816 17920 20868
rect 19524 20995 19576 21004
rect 19524 20961 19533 20995
rect 19533 20961 19567 20995
rect 19567 20961 19576 20995
rect 19524 20952 19576 20961
rect 19708 20995 19760 21004
rect 24032 21020 24084 21072
rect 30380 21088 30432 21140
rect 19708 20961 19753 20995
rect 19753 20961 19760 20995
rect 19708 20952 19760 20961
rect 20628 20952 20680 21004
rect 21272 20995 21324 21004
rect 21272 20961 21281 20995
rect 21281 20961 21315 20995
rect 21315 20961 21324 20995
rect 21272 20952 21324 20961
rect 19984 20884 20036 20936
rect 20720 20884 20772 20936
rect 21824 20952 21876 21004
rect 25320 20995 25372 21004
rect 25320 20961 25329 20995
rect 25329 20961 25363 20995
rect 25363 20961 25372 20995
rect 25320 20952 25372 20961
rect 25504 20995 25556 21004
rect 25504 20961 25513 20995
rect 25513 20961 25547 20995
rect 25547 20961 25556 20995
rect 25504 20952 25556 20961
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 25872 20884 25924 20936
rect 27068 20952 27120 21004
rect 29184 21020 29236 21072
rect 19800 20816 19852 20868
rect 29460 20816 29512 20868
rect 3332 20791 3384 20800
rect 3332 20757 3341 20791
rect 3341 20757 3375 20791
rect 3375 20757 3384 20791
rect 3332 20748 3384 20757
rect 4804 20791 4856 20800
rect 4804 20757 4813 20791
rect 4813 20757 4847 20791
rect 4847 20757 4856 20791
rect 4804 20748 4856 20757
rect 7840 20791 7892 20800
rect 7840 20757 7849 20791
rect 7849 20757 7883 20791
rect 7883 20757 7892 20791
rect 7840 20748 7892 20757
rect 8208 20791 8260 20800
rect 8208 20757 8217 20791
rect 8217 20757 8251 20791
rect 8251 20757 8260 20791
rect 8208 20748 8260 20757
rect 11060 20748 11112 20800
rect 13268 20748 13320 20800
rect 14188 20791 14240 20800
rect 14188 20757 14197 20791
rect 14197 20757 14231 20791
rect 14231 20757 14240 20791
rect 14188 20748 14240 20757
rect 15200 20748 15252 20800
rect 18052 20748 18104 20800
rect 18512 20748 18564 20800
rect 20996 20791 21048 20800
rect 20996 20757 21005 20791
rect 21005 20757 21039 20791
rect 21039 20757 21048 20791
rect 20996 20748 21048 20757
rect 25320 20748 25372 20800
rect 25964 20748 26016 20800
rect 28356 20791 28408 20800
rect 28356 20757 28365 20791
rect 28365 20757 28399 20791
rect 28399 20757 28408 20791
rect 28356 20748 28408 20757
rect 29368 20748 29420 20800
rect 30012 20748 30064 20800
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 11436 20646 11488 20698
rect 11500 20646 11552 20698
rect 11564 20646 11616 20698
rect 11628 20646 11680 20698
rect 11692 20646 11744 20698
rect 19210 20646 19262 20698
rect 19274 20646 19326 20698
rect 19338 20646 19390 20698
rect 19402 20646 19454 20698
rect 19466 20646 19518 20698
rect 26984 20646 27036 20698
rect 27048 20646 27100 20698
rect 27112 20646 27164 20698
rect 27176 20646 27228 20698
rect 27240 20646 27292 20698
rect 1400 20544 1452 20596
rect 4160 20544 4212 20596
rect 4896 20544 4948 20596
rect 6920 20544 6972 20596
rect 3240 20451 3292 20460
rect 3240 20417 3249 20451
rect 3249 20417 3283 20451
rect 3283 20417 3292 20451
rect 3240 20408 3292 20417
rect 1308 20383 1360 20392
rect 1308 20349 1317 20383
rect 1317 20349 1351 20383
rect 1351 20349 1360 20383
rect 1308 20340 1360 20349
rect 3884 20340 3936 20392
rect 9680 20544 9732 20596
rect 12900 20544 12952 20596
rect 14556 20544 14608 20596
rect 14832 20544 14884 20596
rect 9404 20476 9456 20528
rect 5448 20340 5500 20392
rect 9588 20408 9640 20460
rect 9956 20408 10008 20460
rect 6920 20340 6972 20392
rect 8116 20383 8168 20392
rect 8116 20349 8125 20383
rect 8125 20349 8159 20383
rect 8159 20349 8168 20383
rect 8116 20340 8168 20349
rect 8300 20340 8352 20392
rect 12624 20408 12676 20460
rect 13176 20408 13228 20460
rect 2320 20272 2372 20324
rect 3056 20272 3108 20324
rect 5908 20315 5960 20324
rect 5908 20281 5942 20315
rect 5942 20281 5960 20315
rect 5908 20272 5960 20281
rect 6736 20272 6788 20324
rect 2780 20204 2832 20256
rect 3608 20204 3660 20256
rect 3976 20204 4028 20256
rect 6092 20204 6144 20256
rect 9496 20272 9548 20324
rect 9128 20204 9180 20256
rect 9588 20204 9640 20256
rect 9956 20272 10008 20324
rect 12992 20340 13044 20392
rect 13452 20476 13504 20528
rect 13912 20476 13964 20528
rect 14280 20476 14332 20528
rect 14648 20476 14700 20528
rect 16488 20544 16540 20596
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 17776 20544 17828 20596
rect 18512 20544 18564 20596
rect 18788 20544 18840 20596
rect 18972 20544 19024 20596
rect 19984 20544 20036 20596
rect 20904 20544 20956 20596
rect 21548 20544 21600 20596
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 15476 20476 15528 20528
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 18696 20519 18748 20528
rect 18696 20485 18705 20519
rect 18705 20485 18739 20519
rect 18739 20485 18748 20519
rect 18696 20476 18748 20485
rect 19708 20476 19760 20528
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16212 20451 16264 20460
rect 16212 20417 16246 20451
rect 16246 20417 16264 20451
rect 16212 20408 16264 20417
rect 12808 20272 12860 20324
rect 13636 20272 13688 20324
rect 13820 20272 13872 20324
rect 14280 20340 14332 20392
rect 16396 20383 16448 20392
rect 16396 20349 16405 20383
rect 16405 20349 16439 20383
rect 16439 20349 16448 20383
rect 16396 20340 16448 20349
rect 17868 20408 17920 20460
rect 18880 20408 18932 20460
rect 19064 20408 19116 20460
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 18144 20383 18196 20392
rect 18144 20349 18153 20383
rect 18153 20349 18187 20383
rect 18187 20349 18196 20383
rect 18144 20340 18196 20349
rect 15292 20272 15344 20324
rect 17960 20272 18012 20324
rect 18512 20272 18564 20324
rect 20352 20340 20404 20392
rect 20536 20340 20588 20392
rect 10140 20204 10192 20256
rect 11980 20247 12032 20256
rect 11980 20213 11989 20247
rect 11989 20213 12023 20247
rect 12023 20213 12032 20247
rect 11980 20204 12032 20213
rect 12532 20247 12584 20256
rect 12532 20213 12541 20247
rect 12541 20213 12575 20247
rect 12575 20213 12584 20247
rect 12532 20204 12584 20213
rect 14188 20204 14240 20256
rect 15200 20204 15252 20256
rect 19156 20204 19208 20256
rect 20720 20383 20772 20392
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 21088 20408 21140 20460
rect 20996 20340 21048 20392
rect 21272 20340 21324 20392
rect 21548 20340 21600 20392
rect 23664 20408 23716 20460
rect 25872 20544 25924 20596
rect 23388 20383 23440 20392
rect 23388 20349 23397 20383
rect 23397 20349 23431 20383
rect 23431 20349 23440 20383
rect 23388 20340 23440 20349
rect 21916 20204 21968 20256
rect 22928 20247 22980 20256
rect 22928 20213 22937 20247
rect 22937 20213 22971 20247
rect 22971 20213 22980 20247
rect 22928 20204 22980 20213
rect 24584 20272 24636 20324
rect 25964 20340 26016 20392
rect 29000 20383 29052 20392
rect 29000 20349 29009 20383
rect 29009 20349 29043 20383
rect 29043 20349 29052 20383
rect 29000 20340 29052 20349
rect 29276 20383 29328 20392
rect 29276 20349 29310 20383
rect 29310 20349 29328 20383
rect 29276 20340 29328 20349
rect 25412 20204 25464 20256
rect 26608 20204 26660 20256
rect 26700 20204 26752 20256
rect 29092 20204 29144 20256
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 12096 20102 12148 20154
rect 12160 20102 12212 20154
rect 12224 20102 12276 20154
rect 12288 20102 12340 20154
rect 12352 20102 12404 20154
rect 19870 20102 19922 20154
rect 19934 20102 19986 20154
rect 19998 20102 20050 20154
rect 20062 20102 20114 20154
rect 20126 20102 20178 20154
rect 27644 20102 27696 20154
rect 27708 20102 27760 20154
rect 27772 20102 27824 20154
rect 27836 20102 27888 20154
rect 27900 20102 27952 20154
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 2780 20000 2832 20052
rect 3056 20000 3108 20052
rect 3148 20000 3200 20052
rect 2044 19907 2096 19916
rect 2044 19873 2053 19907
rect 2053 19873 2087 19907
rect 2087 19873 2096 19907
rect 2044 19864 2096 19873
rect 2872 19932 2924 19984
rect 4804 19932 4856 19984
rect 5448 20043 5500 20052
rect 5448 20009 5457 20043
rect 5457 20009 5491 20043
rect 5491 20009 5500 20043
rect 5448 20000 5500 20009
rect 5908 20000 5960 20052
rect 2136 19703 2188 19712
rect 2136 19669 2145 19703
rect 2145 19669 2179 19703
rect 2179 19669 2188 19703
rect 2136 19660 2188 19669
rect 3516 19864 3568 19916
rect 3884 19907 3936 19916
rect 3884 19873 3893 19907
rect 3893 19873 3927 19907
rect 3927 19873 3936 19907
rect 3884 19864 3936 19873
rect 3976 19907 4028 19916
rect 3976 19873 3985 19907
rect 3985 19873 4019 19907
rect 4019 19873 4028 19907
rect 3976 19864 4028 19873
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 5356 19907 5408 19916
rect 5356 19873 5365 19907
rect 5365 19873 5399 19907
rect 5399 19873 5408 19907
rect 5356 19864 5408 19873
rect 5816 19864 5868 19916
rect 6092 19907 6144 19916
rect 6092 19873 6101 19907
rect 6101 19873 6135 19907
rect 6135 19873 6144 19907
rect 6092 19864 6144 19873
rect 6276 19907 6328 19916
rect 6276 19873 6285 19907
rect 6285 19873 6319 19907
rect 6319 19873 6328 19907
rect 6276 19864 6328 19873
rect 7012 20000 7064 20052
rect 9680 20000 9732 20052
rect 14648 20000 14700 20052
rect 8852 19932 8904 19984
rect 3148 19796 3200 19848
rect 7012 19796 7064 19848
rect 8024 19728 8076 19780
rect 3148 19660 3200 19712
rect 3240 19703 3292 19712
rect 3240 19669 3249 19703
rect 3249 19669 3283 19703
rect 3283 19669 3292 19703
rect 3240 19660 3292 19669
rect 3516 19660 3568 19712
rect 4160 19660 4212 19712
rect 5080 19660 5132 19712
rect 9128 19907 9180 19916
rect 9128 19873 9137 19907
rect 9137 19873 9171 19907
rect 9171 19873 9180 19907
rect 9128 19864 9180 19873
rect 9864 19864 9916 19916
rect 11980 19864 12032 19916
rect 15200 19932 15252 19984
rect 12532 19907 12584 19916
rect 12532 19873 12541 19907
rect 12541 19873 12575 19907
rect 12575 19873 12584 19907
rect 12532 19864 12584 19873
rect 14832 19864 14884 19916
rect 18052 20000 18104 20052
rect 18144 20000 18196 20052
rect 19340 20000 19392 20052
rect 20628 20000 20680 20052
rect 20720 20000 20772 20052
rect 21272 20043 21324 20052
rect 21272 20009 21281 20043
rect 21281 20009 21315 20043
rect 21315 20009 21324 20043
rect 21272 20000 21324 20009
rect 21916 20000 21968 20052
rect 22100 20000 22152 20052
rect 22468 20000 22520 20052
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 15568 19864 15620 19916
rect 16304 19864 16356 19916
rect 17960 19864 18012 19916
rect 18788 19864 18840 19916
rect 19064 19864 19116 19916
rect 19340 19864 19392 19916
rect 19616 19907 19668 19916
rect 19616 19873 19625 19907
rect 19625 19873 19659 19907
rect 19659 19873 19668 19907
rect 19616 19864 19668 19873
rect 11244 19728 11296 19780
rect 14280 19728 14332 19780
rect 15292 19771 15344 19780
rect 15292 19737 15301 19771
rect 15301 19737 15335 19771
rect 15335 19737 15344 19771
rect 15292 19728 15344 19737
rect 16028 19728 16080 19780
rect 20444 19796 20496 19848
rect 21088 19907 21140 19916
rect 21088 19873 21097 19907
rect 21097 19873 21131 19907
rect 21131 19873 21140 19907
rect 21088 19864 21140 19873
rect 21180 19864 21232 19916
rect 21640 19907 21692 19916
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 22928 19932 22980 19984
rect 21824 19864 21876 19916
rect 22192 19907 22244 19916
rect 22192 19873 22201 19907
rect 22201 19873 22235 19907
rect 22235 19873 22244 19907
rect 22192 19864 22244 19873
rect 16856 19728 16908 19780
rect 18696 19728 18748 19780
rect 18880 19728 18932 19780
rect 19800 19728 19852 19780
rect 22100 19796 22152 19848
rect 21088 19728 21140 19780
rect 23388 19864 23440 19916
rect 24860 19907 24912 19916
rect 24860 19873 24869 19907
rect 24869 19873 24903 19907
rect 24903 19873 24912 19907
rect 24860 19864 24912 19873
rect 24952 19907 25004 19916
rect 24952 19873 24961 19907
rect 24961 19873 24995 19907
rect 24995 19873 25004 19907
rect 24952 19864 25004 19873
rect 26332 20000 26384 20052
rect 25504 19932 25556 19984
rect 10876 19660 10928 19712
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 15476 19660 15528 19712
rect 16488 19660 16540 19712
rect 16580 19703 16632 19712
rect 16580 19669 16589 19703
rect 16589 19669 16623 19703
rect 16623 19669 16632 19703
rect 16580 19660 16632 19669
rect 16764 19703 16816 19712
rect 16764 19669 16773 19703
rect 16773 19669 16807 19703
rect 16807 19669 16816 19703
rect 16764 19660 16816 19669
rect 18052 19660 18104 19712
rect 19708 19703 19760 19712
rect 19708 19669 19717 19703
rect 19717 19669 19751 19703
rect 19751 19669 19760 19703
rect 19708 19660 19760 19669
rect 20352 19660 20404 19712
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 25320 19907 25372 19916
rect 25320 19873 25329 19907
rect 25329 19873 25363 19907
rect 25363 19873 25372 19907
rect 25320 19864 25372 19873
rect 25412 19864 25464 19916
rect 25964 19864 26016 19916
rect 26608 20000 26660 20052
rect 26700 19975 26752 19984
rect 26700 19941 26709 19975
rect 26709 19941 26743 19975
rect 26743 19941 26752 19975
rect 26700 19932 26752 19941
rect 26516 19864 26568 19916
rect 26792 19907 26844 19916
rect 26792 19873 26801 19907
rect 26801 19873 26835 19907
rect 26835 19873 26844 19907
rect 26792 19864 26844 19873
rect 28356 20000 28408 20052
rect 29092 19975 29144 19984
rect 29092 19941 29101 19975
rect 29101 19941 29135 19975
rect 29135 19941 29144 19975
rect 29092 19932 29144 19941
rect 30104 19975 30156 19984
rect 30104 19941 30113 19975
rect 30113 19941 30147 19975
rect 30147 19941 30156 19975
rect 30104 19932 30156 19941
rect 27988 19864 28040 19916
rect 28172 19907 28224 19916
rect 28172 19873 28181 19907
rect 28181 19873 28215 19907
rect 28215 19873 28224 19907
rect 28172 19864 28224 19873
rect 29368 19907 29420 19916
rect 25504 19771 25556 19780
rect 25504 19737 25513 19771
rect 25513 19737 25547 19771
rect 25547 19737 25556 19771
rect 25504 19728 25556 19737
rect 29368 19873 29376 19907
rect 29376 19873 29410 19907
rect 29410 19873 29420 19907
rect 29368 19864 29420 19873
rect 29460 19907 29512 19916
rect 29460 19873 29469 19907
rect 29469 19873 29503 19907
rect 29503 19873 29512 19907
rect 29460 19864 29512 19873
rect 29736 19907 29788 19916
rect 29736 19873 29745 19907
rect 29745 19873 29779 19907
rect 29779 19873 29788 19907
rect 29736 19864 29788 19873
rect 25596 19703 25648 19712
rect 25596 19669 25605 19703
rect 25605 19669 25639 19703
rect 25639 19669 25648 19703
rect 25596 19660 25648 19669
rect 26240 19660 26292 19712
rect 27712 19703 27764 19712
rect 27712 19669 27721 19703
rect 27721 19669 27755 19703
rect 27755 19669 27764 19703
rect 27712 19660 27764 19669
rect 29092 19660 29144 19712
rect 30196 19660 30248 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 11436 19558 11488 19610
rect 11500 19558 11552 19610
rect 11564 19558 11616 19610
rect 11628 19558 11680 19610
rect 11692 19558 11744 19610
rect 19210 19558 19262 19610
rect 19274 19558 19326 19610
rect 19338 19558 19390 19610
rect 19402 19558 19454 19610
rect 19466 19558 19518 19610
rect 26984 19558 27036 19610
rect 27048 19558 27100 19610
rect 27112 19558 27164 19610
rect 27176 19558 27228 19610
rect 27240 19558 27292 19610
rect 3240 19456 3292 19508
rect 4068 19456 4120 19508
rect 7564 19456 7616 19508
rect 9588 19456 9640 19508
rect 9956 19499 10008 19508
rect 9956 19465 9965 19499
rect 9965 19465 9999 19499
rect 9999 19465 10008 19499
rect 9956 19456 10008 19465
rect 11980 19456 12032 19508
rect 14280 19456 14332 19508
rect 16304 19499 16356 19508
rect 16304 19465 16313 19499
rect 16313 19465 16347 19499
rect 16347 19465 16356 19499
rect 16304 19456 16356 19465
rect 16580 19456 16632 19508
rect 17040 19456 17092 19508
rect 18788 19499 18840 19508
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 2044 19388 2096 19440
rect 4712 19388 4764 19440
rect 7932 19388 7984 19440
rect 1400 19252 1452 19304
rect 2136 19252 2188 19304
rect 3332 19320 3384 19372
rect 4068 19320 4120 19372
rect 2964 19295 3016 19304
rect 2964 19261 2973 19295
rect 2973 19261 3007 19295
rect 3007 19261 3016 19295
rect 2964 19252 3016 19261
rect 3240 19295 3292 19304
rect 3240 19261 3249 19295
rect 3249 19261 3283 19295
rect 3283 19261 3292 19295
rect 3240 19252 3292 19261
rect 5080 19320 5132 19372
rect 5724 19252 5776 19304
rect 2504 19227 2556 19236
rect 2504 19193 2513 19227
rect 2513 19193 2547 19227
rect 2547 19193 2556 19227
rect 2504 19184 2556 19193
rect 4068 19184 4120 19236
rect 6920 19184 6972 19236
rect 15844 19388 15896 19440
rect 1584 19116 1636 19168
rect 3332 19116 3384 19168
rect 4804 19116 4856 19168
rect 7564 19116 7616 19168
rect 7748 19227 7800 19236
rect 7748 19193 7757 19227
rect 7757 19193 7791 19227
rect 7791 19193 7800 19227
rect 7748 19184 7800 19193
rect 8024 19252 8076 19304
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 8576 19295 8628 19304
rect 8576 19261 8585 19295
rect 8585 19261 8619 19295
rect 8619 19261 8628 19295
rect 8576 19252 8628 19261
rect 8668 19252 8720 19304
rect 9220 19252 9272 19304
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 10324 19295 10376 19304
rect 10324 19261 10333 19295
rect 10333 19261 10367 19295
rect 10367 19261 10376 19295
rect 10324 19252 10376 19261
rect 8944 19184 8996 19236
rect 14096 19320 14148 19372
rect 14924 19320 14976 19372
rect 15936 19320 15988 19372
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 10692 19297 10744 19304
rect 10692 19263 10701 19297
rect 10701 19263 10735 19297
rect 10735 19263 10744 19297
rect 10692 19252 10744 19263
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 15016 19295 15068 19304
rect 15016 19261 15025 19295
rect 15025 19261 15059 19295
rect 15059 19261 15068 19295
rect 15016 19252 15068 19261
rect 16948 19320 17000 19372
rect 16304 19252 16356 19304
rect 10508 19184 10560 19236
rect 13912 19184 13964 19236
rect 16028 19184 16080 19236
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 17500 19320 17552 19372
rect 20536 19456 20588 19508
rect 21640 19456 21692 19508
rect 25596 19456 25648 19508
rect 25964 19456 26016 19508
rect 26792 19456 26844 19508
rect 28172 19456 28224 19508
rect 20444 19388 20496 19440
rect 19708 19320 19760 19372
rect 20628 19320 20680 19372
rect 24860 19388 24912 19440
rect 27712 19388 27764 19440
rect 14004 19116 14056 19168
rect 15660 19116 15712 19168
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 18144 19295 18196 19304
rect 18144 19261 18153 19295
rect 18153 19261 18187 19295
rect 18187 19261 18196 19295
rect 18144 19252 18196 19261
rect 17224 19227 17276 19236
rect 17224 19193 17233 19227
rect 17233 19193 17267 19227
rect 17267 19193 17276 19227
rect 17224 19184 17276 19193
rect 17316 19184 17368 19236
rect 18328 19252 18380 19304
rect 21088 19252 21140 19304
rect 21548 19295 21600 19304
rect 21548 19261 21557 19295
rect 21557 19261 21591 19295
rect 21591 19261 21600 19295
rect 21548 19252 21600 19261
rect 25688 19252 25740 19304
rect 25872 19320 25924 19372
rect 25964 19252 26016 19304
rect 26332 19320 26384 19372
rect 29184 19388 29236 19440
rect 27344 19252 27396 19304
rect 29000 19295 29052 19304
rect 29000 19261 29009 19295
rect 29009 19261 29043 19295
rect 29043 19261 29052 19295
rect 29000 19252 29052 19261
rect 26056 19227 26108 19236
rect 26056 19193 26065 19227
rect 26065 19193 26099 19227
rect 26099 19193 26108 19227
rect 26056 19184 26108 19193
rect 28448 19227 28500 19236
rect 28448 19193 28457 19227
rect 28457 19193 28491 19227
rect 28491 19193 28500 19227
rect 28448 19184 28500 19193
rect 29552 19227 29604 19236
rect 29552 19193 29586 19227
rect 29586 19193 29604 19227
rect 29552 19184 29604 19193
rect 17132 19116 17184 19168
rect 18972 19116 19024 19168
rect 24952 19116 25004 19168
rect 25320 19116 25372 19168
rect 26240 19116 26292 19168
rect 26424 19116 26476 19168
rect 26884 19116 26936 19168
rect 29000 19116 29052 19168
rect 29368 19116 29420 19168
rect 29460 19116 29512 19168
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 12096 19014 12148 19066
rect 12160 19014 12212 19066
rect 12224 19014 12276 19066
rect 12288 19014 12340 19066
rect 12352 19014 12404 19066
rect 19870 19014 19922 19066
rect 19934 19014 19986 19066
rect 19998 19014 20050 19066
rect 20062 19014 20114 19066
rect 20126 19014 20178 19066
rect 27644 19014 27696 19066
rect 27708 19014 27760 19066
rect 27772 19014 27824 19066
rect 27836 19014 27888 19066
rect 27900 19014 27952 19066
rect 3240 18912 3292 18964
rect 5724 18912 5776 18964
rect 8392 18912 8444 18964
rect 9128 18912 9180 18964
rect 9312 18912 9364 18964
rect 10508 18912 10560 18964
rect 10600 18912 10652 18964
rect 3148 18844 3200 18896
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 3332 18819 3384 18828
rect 3332 18785 3341 18819
rect 3341 18785 3375 18819
rect 3375 18785 3384 18819
rect 3332 18776 3384 18785
rect 3424 18819 3476 18828
rect 3424 18785 3433 18819
rect 3433 18785 3467 18819
rect 3467 18785 3476 18819
rect 3424 18776 3476 18785
rect 8944 18844 8996 18896
rect 4068 18776 4120 18828
rect 5908 18776 5960 18828
rect 6460 18776 6512 18828
rect 7748 18776 7800 18828
rect 9036 18776 9088 18828
rect 9312 18819 9364 18828
rect 9312 18785 9321 18819
rect 9321 18785 9355 18819
rect 9355 18785 9364 18819
rect 9312 18776 9364 18785
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 4252 18640 4304 18692
rect 4988 18751 5040 18760
rect 4988 18717 4997 18751
rect 4997 18717 5031 18751
rect 5031 18717 5040 18751
rect 4988 18708 5040 18717
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 6920 18708 6972 18760
rect 10232 18844 10284 18896
rect 10324 18844 10376 18896
rect 11060 18844 11112 18896
rect 14740 18912 14792 18964
rect 15200 18912 15252 18964
rect 15752 18912 15804 18964
rect 16488 18912 16540 18964
rect 16672 18912 16724 18964
rect 18144 18912 18196 18964
rect 9772 18776 9824 18828
rect 10508 18819 10560 18828
rect 10508 18785 10517 18819
rect 10517 18785 10551 18819
rect 10551 18785 10560 18819
rect 10508 18776 10560 18785
rect 11152 18819 11204 18828
rect 11152 18785 11161 18819
rect 11161 18785 11195 18819
rect 11195 18785 11204 18819
rect 11152 18776 11204 18785
rect 11796 18776 11848 18828
rect 11980 18776 12032 18828
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10692 18708 10744 18760
rect 12440 18776 12492 18828
rect 12624 18844 12676 18896
rect 13820 18844 13872 18896
rect 12808 18819 12860 18828
rect 12808 18785 12817 18819
rect 12817 18785 12851 18819
rect 12851 18785 12860 18819
rect 12808 18776 12860 18785
rect 13728 18776 13780 18828
rect 14924 18776 14976 18828
rect 15568 18819 15620 18828
rect 15568 18785 15577 18819
rect 15577 18785 15611 18819
rect 15611 18785 15620 18819
rect 15568 18776 15620 18785
rect 15936 18776 15988 18828
rect 17040 18844 17092 18896
rect 21088 18844 21140 18896
rect 12992 18708 13044 18760
rect 14556 18708 14608 18760
rect 15660 18708 15712 18760
rect 16488 18819 16540 18828
rect 16488 18785 16497 18819
rect 16497 18785 16531 18819
rect 16531 18785 16540 18819
rect 16488 18776 16540 18785
rect 17224 18776 17276 18828
rect 18696 18819 18748 18828
rect 18696 18785 18705 18819
rect 18705 18785 18739 18819
rect 18739 18785 18748 18819
rect 18696 18776 18748 18785
rect 18788 18776 18840 18828
rect 19064 18776 19116 18828
rect 20628 18776 20680 18828
rect 16764 18708 16816 18760
rect 24860 18912 24912 18964
rect 25688 18912 25740 18964
rect 27988 18912 28040 18964
rect 28080 18912 28132 18964
rect 22376 18887 22428 18896
rect 22376 18853 22394 18887
rect 22394 18853 22428 18887
rect 22376 18844 22428 18853
rect 22008 18776 22060 18828
rect 28724 18844 28776 18896
rect 29552 18912 29604 18964
rect 8852 18640 8904 18692
rect 9496 18640 9548 18692
rect 4160 18572 4212 18624
rect 4804 18572 4856 18624
rect 5172 18615 5224 18624
rect 5172 18581 5181 18615
rect 5181 18581 5215 18615
rect 5215 18581 5224 18615
rect 5172 18572 5224 18581
rect 6000 18615 6052 18624
rect 6000 18581 6009 18615
rect 6009 18581 6043 18615
rect 6043 18581 6052 18615
rect 6000 18572 6052 18581
rect 8576 18572 8628 18624
rect 10232 18615 10284 18624
rect 10232 18581 10241 18615
rect 10241 18581 10275 18615
rect 10275 18581 10284 18615
rect 10232 18572 10284 18581
rect 13084 18640 13136 18692
rect 16948 18640 17000 18692
rect 11980 18572 12032 18624
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 15844 18572 15896 18624
rect 16120 18572 16172 18624
rect 17040 18572 17092 18624
rect 19064 18572 19116 18624
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 21364 18572 21416 18624
rect 23480 18708 23532 18760
rect 24032 18751 24084 18760
rect 24032 18717 24041 18751
rect 24041 18717 24075 18751
rect 24075 18717 24084 18751
rect 24032 18708 24084 18717
rect 26424 18819 26476 18828
rect 26424 18785 26433 18819
rect 26433 18785 26467 18819
rect 26467 18785 26476 18819
rect 26424 18776 26476 18785
rect 26516 18776 26568 18828
rect 24860 18751 24912 18760
rect 24860 18717 24878 18751
rect 24878 18717 24912 18751
rect 24860 18708 24912 18717
rect 24952 18751 25004 18760
rect 24952 18717 24961 18751
rect 24961 18717 24995 18751
rect 24995 18717 25004 18751
rect 24952 18708 25004 18717
rect 25872 18751 25924 18760
rect 25872 18717 25881 18751
rect 25881 18717 25915 18751
rect 25915 18717 25924 18751
rect 25872 18708 25924 18717
rect 28816 18819 28868 18828
rect 28816 18785 28825 18819
rect 28825 18785 28859 18819
rect 28859 18785 28868 18819
rect 28816 18776 28868 18785
rect 29460 18844 29512 18896
rect 29000 18819 29052 18828
rect 29000 18785 29009 18819
rect 29009 18785 29043 18819
rect 29043 18785 29052 18819
rect 29000 18776 29052 18785
rect 29368 18819 29420 18828
rect 29368 18785 29377 18819
rect 29377 18785 29411 18819
rect 29411 18785 29420 18819
rect 29368 18776 29420 18785
rect 29184 18708 29236 18760
rect 29644 18819 29696 18828
rect 29644 18785 29678 18819
rect 29678 18785 29696 18819
rect 29644 18776 29696 18785
rect 30196 18776 30248 18828
rect 25228 18683 25280 18692
rect 25228 18649 25237 18683
rect 25237 18649 25271 18683
rect 25271 18649 25280 18683
rect 25228 18640 25280 18649
rect 27712 18572 27764 18624
rect 28356 18572 28408 18624
rect 28724 18572 28776 18624
rect 31024 18615 31076 18624
rect 31024 18581 31033 18615
rect 31033 18581 31067 18615
rect 31067 18581 31076 18615
rect 31024 18572 31076 18581
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 11436 18470 11488 18522
rect 11500 18470 11552 18522
rect 11564 18470 11616 18522
rect 11628 18470 11680 18522
rect 11692 18470 11744 18522
rect 19210 18470 19262 18522
rect 19274 18470 19326 18522
rect 19338 18470 19390 18522
rect 19402 18470 19454 18522
rect 19466 18470 19518 18522
rect 26984 18470 27036 18522
rect 27048 18470 27100 18522
rect 27112 18470 27164 18522
rect 27176 18470 27228 18522
rect 27240 18470 27292 18522
rect 4988 18368 5040 18420
rect 5172 18411 5224 18420
rect 5172 18377 5181 18411
rect 5181 18377 5215 18411
rect 5215 18377 5224 18411
rect 5172 18368 5224 18377
rect 6276 18368 6328 18420
rect 8024 18368 8076 18420
rect 9864 18368 9916 18420
rect 3240 18164 3292 18216
rect 3516 18207 3568 18216
rect 3516 18173 3525 18207
rect 3525 18173 3559 18207
rect 3559 18173 3568 18207
rect 3516 18164 3568 18173
rect 3884 18164 3936 18216
rect 4068 18232 4120 18284
rect 4804 18164 4856 18216
rect 4988 18207 5040 18216
rect 4988 18173 4997 18207
rect 4997 18173 5031 18207
rect 5031 18173 5040 18207
rect 4988 18164 5040 18173
rect 9036 18300 9088 18352
rect 9312 18300 9364 18352
rect 10048 18368 10100 18420
rect 5356 18164 5408 18216
rect 2780 18096 2832 18148
rect 3424 18096 3476 18148
rect 4252 18096 4304 18148
rect 5816 18232 5868 18284
rect 6000 18207 6052 18216
rect 6000 18173 6009 18207
rect 6009 18173 6043 18207
rect 6043 18173 6052 18207
rect 6000 18164 6052 18173
rect 6184 18164 6236 18216
rect 6460 18207 6512 18216
rect 6460 18173 6469 18207
rect 6469 18173 6503 18207
rect 6503 18173 6512 18207
rect 6460 18164 6512 18173
rect 8944 18232 8996 18284
rect 9220 18232 9272 18284
rect 3240 18028 3292 18080
rect 5632 18096 5684 18148
rect 8300 18164 8352 18216
rect 9956 18232 10008 18284
rect 10508 18300 10560 18352
rect 10140 18232 10192 18284
rect 4804 18028 4856 18080
rect 5172 18028 5224 18080
rect 6184 18028 6236 18080
rect 6460 18028 6512 18080
rect 6828 18028 6880 18080
rect 8668 18028 8720 18080
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 9496 18071 9548 18080
rect 9496 18037 9505 18071
rect 9505 18037 9539 18071
rect 9539 18037 9548 18071
rect 9496 18028 9548 18037
rect 9864 18139 9916 18148
rect 9864 18105 9873 18139
rect 9873 18105 9907 18139
rect 9907 18105 9916 18139
rect 9864 18096 9916 18105
rect 10600 18207 10652 18216
rect 10600 18173 10609 18207
rect 10609 18173 10643 18207
rect 10643 18173 10652 18207
rect 10600 18164 10652 18173
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 10784 18207 10836 18216
rect 10784 18173 10793 18207
rect 10793 18173 10827 18207
rect 10827 18173 10836 18207
rect 10784 18164 10836 18173
rect 10876 18164 10928 18216
rect 15476 18300 15528 18352
rect 15568 18300 15620 18352
rect 18972 18300 19024 18352
rect 20628 18411 20680 18420
rect 20628 18377 20637 18411
rect 20637 18377 20671 18411
rect 20671 18377 20680 18411
rect 20628 18368 20680 18377
rect 24584 18368 24636 18420
rect 25780 18368 25832 18420
rect 26516 18368 26568 18420
rect 28816 18411 28868 18420
rect 28816 18377 28825 18411
rect 28825 18377 28859 18411
rect 28859 18377 28868 18411
rect 28816 18368 28868 18377
rect 20904 18300 20956 18352
rect 22008 18300 22060 18352
rect 28356 18300 28408 18352
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 11612 18164 11664 18216
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 14188 18232 14240 18284
rect 13360 18164 13412 18216
rect 13912 18164 13964 18216
rect 15936 18232 15988 18284
rect 15016 18139 15068 18148
rect 15016 18105 15025 18139
rect 15025 18105 15059 18139
rect 15059 18105 15068 18139
rect 15016 18096 15068 18105
rect 15752 18207 15804 18216
rect 15752 18173 15761 18207
rect 15761 18173 15795 18207
rect 15795 18173 15804 18207
rect 15752 18164 15804 18173
rect 15844 18207 15896 18216
rect 15844 18173 15853 18207
rect 15853 18173 15887 18207
rect 15887 18173 15896 18207
rect 17040 18232 17092 18284
rect 15844 18164 15896 18173
rect 16212 18164 16264 18216
rect 16304 18207 16356 18216
rect 16304 18173 16313 18207
rect 16313 18173 16347 18207
rect 16347 18173 16356 18207
rect 16304 18164 16356 18173
rect 16488 18207 16540 18216
rect 16488 18173 16497 18207
rect 16497 18173 16531 18207
rect 16531 18173 16540 18207
rect 16488 18164 16540 18173
rect 16856 18164 16908 18216
rect 18880 18164 18932 18216
rect 18972 18207 19024 18216
rect 18972 18173 18981 18207
rect 18981 18173 19015 18207
rect 19015 18173 19024 18207
rect 18972 18164 19024 18173
rect 19340 18164 19392 18216
rect 9956 18071 10008 18080
rect 9956 18037 9965 18071
rect 9965 18037 9999 18071
rect 9999 18037 10008 18071
rect 9956 18028 10008 18037
rect 10140 18028 10192 18080
rect 12624 18071 12676 18080
rect 12624 18037 12633 18071
rect 12633 18037 12667 18071
rect 12667 18037 12676 18071
rect 12624 18028 12676 18037
rect 13636 18028 13688 18080
rect 15660 18028 15712 18080
rect 15844 18028 15896 18080
rect 17316 18096 17368 18148
rect 19524 18139 19576 18148
rect 19524 18105 19558 18139
rect 19558 18105 19576 18139
rect 19524 18096 19576 18105
rect 19616 18096 19668 18148
rect 19800 18096 19852 18148
rect 20628 18096 20680 18148
rect 21364 18164 21416 18216
rect 21824 18164 21876 18216
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 18696 18028 18748 18080
rect 19064 18028 19116 18080
rect 19432 18028 19484 18080
rect 20444 18028 20496 18080
rect 23480 18207 23532 18216
rect 23480 18173 23489 18207
rect 23489 18173 23523 18207
rect 23523 18173 23532 18207
rect 23480 18164 23532 18173
rect 24400 18164 24452 18216
rect 25504 18207 25556 18216
rect 25504 18173 25513 18207
rect 25513 18173 25547 18207
rect 25547 18173 25556 18207
rect 25504 18164 25556 18173
rect 25596 18164 25648 18216
rect 25780 18207 25832 18216
rect 25780 18173 25789 18207
rect 25789 18173 25823 18207
rect 25823 18173 25832 18207
rect 25780 18164 25832 18173
rect 25872 18207 25924 18216
rect 25872 18173 25881 18207
rect 25881 18173 25915 18207
rect 25915 18173 25924 18207
rect 25872 18164 25924 18173
rect 28080 18232 28132 18284
rect 24124 18139 24176 18148
rect 24124 18105 24158 18139
rect 24158 18105 24176 18139
rect 24124 18096 24176 18105
rect 24860 18096 24912 18148
rect 26700 18207 26752 18216
rect 26700 18173 26709 18207
rect 26709 18173 26743 18207
rect 26743 18173 26752 18207
rect 26700 18164 26752 18173
rect 26884 18207 26936 18216
rect 26884 18173 26893 18207
rect 26893 18173 26927 18207
rect 26927 18173 26936 18207
rect 26884 18164 26936 18173
rect 27988 18207 28040 18216
rect 27988 18173 27997 18207
rect 27997 18173 28031 18207
rect 28031 18173 28040 18207
rect 27988 18164 28040 18173
rect 28172 18164 28224 18216
rect 28448 18232 28500 18284
rect 26792 18096 26844 18148
rect 27712 18096 27764 18148
rect 28540 18207 28592 18216
rect 28540 18173 28549 18207
rect 28549 18173 28583 18207
rect 28583 18173 28592 18207
rect 28540 18164 28592 18173
rect 29644 18368 29696 18420
rect 29368 18300 29420 18352
rect 29552 18275 29604 18284
rect 29552 18241 29561 18275
rect 29561 18241 29595 18275
rect 29595 18241 29604 18275
rect 29552 18232 29604 18241
rect 29000 18096 29052 18148
rect 29092 18096 29144 18148
rect 30380 18164 30432 18216
rect 31024 18164 31076 18216
rect 22284 18028 22336 18080
rect 23296 18028 23348 18080
rect 24952 18028 25004 18080
rect 25136 18028 25188 18080
rect 28080 18028 28132 18080
rect 29276 18028 29328 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 12096 17926 12148 17978
rect 12160 17926 12212 17978
rect 12224 17926 12276 17978
rect 12288 17926 12340 17978
rect 12352 17926 12404 17978
rect 19870 17926 19922 17978
rect 19934 17926 19986 17978
rect 19998 17926 20050 17978
rect 20062 17926 20114 17978
rect 20126 17926 20178 17978
rect 27644 17926 27696 17978
rect 27708 17926 27760 17978
rect 27772 17926 27824 17978
rect 27836 17926 27888 17978
rect 27900 17926 27952 17978
rect 3424 17824 3476 17876
rect 3884 17824 3936 17876
rect 5724 17824 5776 17876
rect 6000 17824 6052 17876
rect 2688 17731 2740 17740
rect 2688 17697 2697 17731
rect 2697 17697 2731 17731
rect 2731 17697 2740 17731
rect 2688 17688 2740 17697
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 4160 17756 4212 17808
rect 4988 17756 5040 17808
rect 3056 17731 3108 17740
rect 3056 17697 3065 17731
rect 3065 17697 3099 17731
rect 3099 17697 3108 17731
rect 3056 17688 3108 17697
rect 3884 17731 3936 17740
rect 3884 17697 3893 17731
rect 3893 17697 3927 17731
rect 3927 17697 3936 17731
rect 3884 17688 3936 17697
rect 4068 17688 4120 17740
rect 4528 17688 4580 17740
rect 5540 17756 5592 17808
rect 6460 17756 6512 17808
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 6644 17756 6696 17808
rect 2412 17527 2464 17536
rect 2412 17493 2421 17527
rect 2421 17493 2455 17527
rect 2455 17493 2464 17527
rect 2412 17484 2464 17493
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 4160 17620 4212 17629
rect 5172 17731 5224 17740
rect 5172 17697 5181 17731
rect 5181 17697 5215 17731
rect 5215 17697 5224 17731
rect 5172 17688 5224 17697
rect 5264 17731 5316 17740
rect 5264 17697 5273 17731
rect 5273 17697 5307 17731
rect 5307 17697 5316 17731
rect 5264 17688 5316 17697
rect 5448 17731 5500 17740
rect 5448 17697 5457 17731
rect 5457 17697 5491 17731
rect 5491 17697 5500 17731
rect 5448 17688 5500 17697
rect 3240 17552 3292 17604
rect 4068 17552 4120 17604
rect 4160 17484 4212 17536
rect 5356 17620 5408 17672
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 6184 17731 6236 17740
rect 6184 17697 6193 17731
rect 6193 17697 6227 17731
rect 6227 17697 6236 17731
rect 6184 17688 6236 17697
rect 6368 17688 6420 17740
rect 5816 17620 5868 17672
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 6736 17731 6788 17740
rect 6736 17697 6745 17731
rect 6745 17697 6779 17731
rect 6779 17697 6788 17731
rect 6736 17688 6788 17697
rect 8760 17756 8812 17808
rect 7104 17688 7156 17740
rect 8576 17731 8628 17740
rect 8576 17697 8585 17731
rect 8585 17697 8619 17731
rect 8619 17697 8628 17731
rect 8576 17688 8628 17697
rect 8668 17731 8720 17740
rect 8668 17697 8677 17731
rect 8677 17697 8711 17731
rect 8711 17697 8720 17731
rect 8668 17688 8720 17697
rect 9680 17756 9732 17808
rect 9864 17824 9916 17876
rect 9864 17688 9916 17740
rect 10232 17824 10284 17876
rect 10692 17824 10744 17876
rect 11152 17824 11204 17876
rect 11612 17824 11664 17876
rect 12440 17824 12492 17876
rect 15016 17824 15068 17876
rect 15936 17824 15988 17876
rect 17132 17824 17184 17876
rect 19340 17824 19392 17876
rect 10048 17620 10100 17672
rect 11336 17731 11388 17740
rect 11336 17697 11345 17731
rect 11345 17697 11379 17731
rect 11379 17697 11388 17731
rect 11336 17688 11388 17697
rect 12716 17756 12768 17808
rect 13636 17799 13688 17808
rect 13636 17765 13645 17799
rect 13645 17765 13679 17799
rect 13679 17765 13688 17799
rect 13636 17756 13688 17765
rect 12072 17688 12124 17740
rect 12532 17688 12584 17740
rect 10600 17620 10652 17672
rect 11612 17663 11664 17672
rect 11612 17629 11621 17663
rect 11621 17629 11655 17663
rect 11655 17629 11664 17663
rect 11612 17620 11664 17629
rect 14464 17731 14516 17740
rect 14464 17697 14473 17731
rect 14473 17697 14507 17731
rect 14507 17697 14516 17731
rect 14464 17688 14516 17697
rect 14556 17620 14608 17672
rect 5264 17552 5316 17604
rect 10508 17552 10560 17604
rect 13360 17595 13412 17604
rect 13360 17561 13369 17595
rect 13369 17561 13403 17595
rect 13403 17561 13412 17595
rect 13360 17552 13412 17561
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 15200 17688 15252 17740
rect 16212 17756 16264 17808
rect 15568 17731 15620 17740
rect 15568 17697 15577 17731
rect 15577 17697 15611 17731
rect 15611 17697 15620 17731
rect 15568 17688 15620 17697
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 16028 17688 16080 17740
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 18420 17688 18472 17740
rect 19432 17756 19484 17808
rect 19524 17799 19576 17808
rect 19524 17765 19533 17799
rect 19533 17765 19567 17799
rect 19567 17765 19576 17799
rect 19524 17756 19576 17765
rect 20628 17756 20680 17808
rect 22560 17799 22612 17808
rect 16764 17620 16816 17672
rect 18144 17620 18196 17672
rect 19064 17731 19116 17740
rect 19064 17697 19073 17731
rect 19073 17697 19107 17731
rect 19107 17697 19116 17731
rect 19064 17688 19116 17697
rect 18972 17620 19024 17672
rect 19248 17731 19300 17740
rect 19248 17697 19257 17731
rect 19257 17697 19291 17731
rect 19291 17697 19300 17731
rect 19248 17688 19300 17697
rect 19616 17688 19668 17740
rect 19708 17688 19760 17740
rect 20720 17731 20772 17740
rect 20720 17697 20729 17731
rect 20729 17697 20763 17731
rect 20763 17697 20772 17731
rect 20720 17688 20772 17697
rect 21088 17688 21140 17740
rect 22560 17765 22569 17799
rect 22569 17765 22603 17799
rect 22603 17765 22612 17799
rect 22560 17756 22612 17765
rect 22192 17731 22244 17740
rect 22192 17697 22201 17731
rect 22201 17697 22235 17731
rect 22235 17697 22244 17731
rect 22192 17688 22244 17697
rect 23940 17824 23992 17876
rect 24124 17824 24176 17876
rect 24860 17824 24912 17876
rect 20812 17620 20864 17672
rect 21272 17552 21324 17604
rect 22560 17620 22612 17672
rect 24124 17688 24176 17740
rect 24400 17731 24452 17740
rect 24400 17697 24409 17731
rect 24409 17697 24443 17731
rect 24443 17697 24452 17731
rect 24400 17688 24452 17697
rect 24308 17552 24360 17604
rect 4344 17484 4396 17536
rect 5540 17484 5592 17536
rect 6276 17484 6328 17536
rect 6920 17484 6972 17536
rect 9588 17484 9640 17536
rect 11336 17484 11388 17536
rect 14372 17484 14424 17536
rect 14924 17484 14976 17536
rect 15200 17527 15252 17536
rect 15200 17493 15209 17527
rect 15209 17493 15243 17527
rect 15243 17493 15252 17527
rect 15200 17484 15252 17493
rect 18696 17484 18748 17536
rect 22008 17484 22060 17536
rect 22928 17484 22980 17536
rect 23204 17484 23256 17536
rect 24676 17731 24728 17740
rect 24676 17697 24685 17731
rect 24685 17697 24719 17731
rect 24719 17697 24728 17731
rect 24676 17688 24728 17697
rect 24768 17688 24820 17740
rect 25412 17756 25464 17808
rect 26056 17756 26108 17808
rect 26148 17731 26200 17740
rect 26148 17697 26157 17731
rect 26157 17697 26191 17731
rect 26191 17697 26200 17731
rect 26148 17688 26200 17697
rect 26240 17731 26292 17740
rect 26240 17697 26249 17731
rect 26249 17697 26283 17731
rect 26283 17697 26292 17731
rect 26240 17688 26292 17697
rect 26700 17824 26752 17876
rect 27344 17756 27396 17808
rect 28540 17824 28592 17876
rect 28080 17756 28132 17808
rect 29000 17867 29052 17876
rect 29000 17833 29009 17867
rect 29009 17833 29043 17867
rect 29043 17833 29052 17867
rect 29000 17824 29052 17833
rect 29460 17824 29512 17876
rect 30288 17824 30340 17876
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 25780 17620 25832 17672
rect 28356 17731 28408 17740
rect 28356 17697 28365 17731
rect 28365 17697 28399 17731
rect 28399 17697 28408 17731
rect 28356 17688 28408 17697
rect 28540 17731 28592 17740
rect 28540 17697 28549 17731
rect 28549 17697 28583 17731
rect 28583 17697 28592 17731
rect 28540 17688 28592 17697
rect 28632 17731 28684 17740
rect 28632 17697 28641 17731
rect 28641 17697 28675 17731
rect 28675 17697 28684 17731
rect 28632 17688 28684 17697
rect 28724 17731 28776 17740
rect 28724 17697 28733 17731
rect 28733 17697 28767 17731
rect 28767 17697 28776 17731
rect 28724 17688 28776 17697
rect 29276 17756 29328 17808
rect 30012 17688 30064 17740
rect 30196 17688 30248 17740
rect 28172 17620 28224 17672
rect 29552 17620 29604 17672
rect 28080 17552 28132 17604
rect 28448 17552 28500 17604
rect 28724 17552 28776 17604
rect 25228 17484 25280 17536
rect 27620 17484 27672 17536
rect 30472 17484 30524 17536
rect 30564 17484 30616 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 11436 17382 11488 17434
rect 11500 17382 11552 17434
rect 11564 17382 11616 17434
rect 11628 17382 11680 17434
rect 11692 17382 11744 17434
rect 19210 17382 19262 17434
rect 19274 17382 19326 17434
rect 19338 17382 19390 17434
rect 19402 17382 19454 17434
rect 19466 17382 19518 17434
rect 26984 17382 27036 17434
rect 27048 17382 27100 17434
rect 27112 17382 27164 17434
rect 27176 17382 27228 17434
rect 27240 17382 27292 17434
rect 3516 17280 3568 17332
rect 4068 17280 4120 17332
rect 5172 17280 5224 17332
rect 6000 17280 6052 17332
rect 2688 17144 2740 17196
rect 3884 17212 3936 17264
rect 6368 17212 6420 17264
rect 2412 17076 2464 17128
rect 4160 17076 4212 17128
rect 4528 17076 4580 17128
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 4804 17076 4856 17085
rect 4988 17119 5040 17128
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 1400 17008 1452 17060
rect 2688 17008 2740 17060
rect 4712 17008 4764 17060
rect 5264 17119 5316 17128
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 5448 17119 5500 17128
rect 5448 17085 5457 17119
rect 5457 17085 5491 17119
rect 5491 17085 5500 17119
rect 5448 17076 5500 17085
rect 6184 17144 6236 17196
rect 6000 17119 6052 17128
rect 6000 17085 6009 17119
rect 6009 17085 6043 17119
rect 6043 17085 6052 17119
rect 6000 17076 6052 17085
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 6276 17119 6328 17128
rect 6276 17085 6285 17119
rect 6285 17085 6319 17119
rect 6319 17085 6328 17119
rect 6276 17076 6328 17085
rect 8300 17280 8352 17332
rect 8300 17144 8352 17196
rect 9864 17255 9916 17264
rect 9864 17221 9873 17255
rect 9873 17221 9907 17255
rect 9907 17221 9916 17255
rect 9864 17212 9916 17221
rect 11336 17280 11388 17332
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 11152 17212 11204 17264
rect 9956 17144 10008 17196
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 3884 16940 3936 16992
rect 4344 16940 4396 16992
rect 5172 16940 5224 16992
rect 5632 17008 5684 17060
rect 5908 17008 5960 17060
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 10048 17076 10100 17128
rect 6736 17008 6788 17060
rect 9404 17008 9456 17060
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 10416 17076 10468 17128
rect 10600 17119 10652 17128
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 11152 17119 11204 17128
rect 11152 17085 11161 17119
rect 11161 17085 11195 17119
rect 11195 17085 11204 17119
rect 11152 17076 11204 17085
rect 12624 17076 12676 17128
rect 13728 17119 13780 17128
rect 13728 17085 13737 17119
rect 13737 17085 13771 17119
rect 13771 17085 13780 17119
rect 13728 17076 13780 17085
rect 13912 17076 13964 17128
rect 11704 17008 11756 17060
rect 15936 17280 15988 17332
rect 16212 17280 16264 17332
rect 20720 17280 20772 17332
rect 23664 17280 23716 17332
rect 24032 17280 24084 17332
rect 25596 17280 25648 17332
rect 25780 17280 25832 17332
rect 26148 17280 26200 17332
rect 28356 17280 28408 17332
rect 30380 17280 30432 17332
rect 14832 17255 14884 17264
rect 14832 17221 14841 17255
rect 14841 17221 14875 17255
rect 14875 17221 14884 17255
rect 14832 17212 14884 17221
rect 14280 17144 14332 17196
rect 14188 17119 14240 17128
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 16304 17076 16356 17128
rect 16948 17076 17000 17128
rect 17776 17076 17828 17128
rect 19432 17212 19484 17264
rect 20260 17255 20312 17264
rect 20260 17221 20269 17255
rect 20269 17221 20303 17255
rect 20303 17221 20312 17255
rect 20260 17212 20312 17221
rect 29552 17212 29604 17264
rect 30288 17212 30340 17264
rect 18604 17144 18656 17196
rect 15936 17008 15988 17060
rect 11612 16940 11664 16992
rect 16764 17008 16816 17060
rect 18696 17119 18748 17128
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 19064 17119 19116 17128
rect 19064 17085 19073 17119
rect 19073 17085 19107 17119
rect 19107 17085 19116 17119
rect 19064 17076 19116 17085
rect 19616 17119 19668 17128
rect 19616 17085 19625 17119
rect 19625 17085 19659 17119
rect 19659 17085 19668 17119
rect 19616 17076 19668 17085
rect 19156 17008 19208 17060
rect 18880 16940 18932 16992
rect 19432 16983 19484 16992
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 19616 16940 19668 16992
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 21088 17187 21140 17196
rect 21088 17153 21106 17187
rect 21106 17153 21140 17187
rect 21088 17144 21140 17153
rect 21456 17187 21508 17196
rect 21456 17153 21465 17187
rect 21465 17153 21499 17187
rect 21499 17153 21508 17187
rect 21456 17144 21508 17153
rect 22560 17144 22612 17196
rect 24952 17144 25004 17196
rect 25964 17144 26016 17196
rect 26148 17144 26200 17196
rect 26792 17144 26844 17196
rect 19800 17076 19852 17128
rect 21180 17119 21232 17128
rect 21180 17085 21189 17119
rect 21189 17085 21223 17119
rect 21223 17085 21232 17119
rect 21180 17076 21232 17085
rect 20352 17008 20404 17060
rect 21456 16940 21508 16992
rect 23296 17119 23348 17128
rect 23296 17085 23314 17119
rect 23314 17085 23348 17119
rect 23296 17076 23348 17085
rect 23480 17076 23532 17128
rect 22284 16940 22336 16992
rect 24492 17119 24544 17128
rect 24492 17085 24501 17119
rect 24501 17085 24535 17119
rect 24535 17085 24544 17119
rect 24492 17076 24544 17085
rect 24768 17076 24820 17128
rect 25872 17076 25924 17128
rect 27344 17076 27396 17128
rect 27988 17144 28040 17196
rect 27620 17119 27672 17128
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 25136 17008 25188 17060
rect 25596 17008 25648 17060
rect 27896 17119 27948 17128
rect 27896 17085 27905 17119
rect 27905 17085 27939 17119
rect 27939 17085 27948 17119
rect 27896 17076 27948 17085
rect 24676 16940 24728 16992
rect 24860 16983 24912 16992
rect 24860 16949 24869 16983
rect 24869 16949 24903 16983
rect 24903 16949 24912 16983
rect 24860 16940 24912 16949
rect 25228 16983 25280 16992
rect 25228 16949 25237 16983
rect 25237 16949 25271 16983
rect 25271 16949 25280 16983
rect 25228 16940 25280 16949
rect 27988 17051 28040 17060
rect 27988 17017 27997 17051
rect 27997 17017 28031 17051
rect 28031 17017 28040 17051
rect 27988 17008 28040 17017
rect 28172 17051 28224 17060
rect 28172 17017 28181 17051
rect 28181 17017 28215 17051
rect 28215 17017 28224 17051
rect 28172 17008 28224 17017
rect 28816 17144 28868 17196
rect 30196 17144 30248 17196
rect 30472 17212 30524 17264
rect 28908 17076 28960 17128
rect 29092 17076 29144 17128
rect 29184 17119 29236 17128
rect 29184 17085 29193 17119
rect 29193 17085 29227 17119
rect 29227 17085 29236 17119
rect 29184 17076 29236 17085
rect 29276 17119 29328 17128
rect 29276 17085 29285 17119
rect 29285 17085 29319 17119
rect 29319 17085 29328 17119
rect 29276 17076 29328 17085
rect 28448 17051 28500 17060
rect 28448 17017 28457 17051
rect 28457 17017 28491 17051
rect 28491 17017 28500 17051
rect 28448 17008 28500 17017
rect 28632 17051 28684 17060
rect 28632 17017 28641 17051
rect 28641 17017 28675 17051
rect 28675 17017 28684 17051
rect 28632 17008 28684 17017
rect 30564 17119 30616 17128
rect 30564 17085 30573 17119
rect 30573 17085 30607 17119
rect 30607 17085 30616 17119
rect 30564 17076 30616 17085
rect 30748 17119 30800 17128
rect 30748 17085 30757 17119
rect 30757 17085 30791 17119
rect 30791 17085 30800 17119
rect 30748 17076 30800 17085
rect 28540 16940 28592 16992
rect 30012 17008 30064 17060
rect 30196 16940 30248 16992
rect 31208 16983 31260 16992
rect 31208 16949 31217 16983
rect 31217 16949 31251 16983
rect 31251 16949 31260 16983
rect 31208 16940 31260 16949
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 12096 16838 12148 16890
rect 12160 16838 12212 16890
rect 12224 16838 12276 16890
rect 12288 16838 12340 16890
rect 12352 16838 12404 16890
rect 19870 16838 19922 16890
rect 19934 16838 19986 16890
rect 19998 16838 20050 16890
rect 20062 16838 20114 16890
rect 20126 16838 20178 16890
rect 27644 16838 27696 16890
rect 27708 16838 27760 16890
rect 27772 16838 27824 16890
rect 27836 16838 27888 16890
rect 27900 16838 27952 16890
rect 3240 16736 3292 16788
rect 4068 16736 4120 16788
rect 4160 16779 4212 16788
rect 4160 16745 4169 16779
rect 4169 16745 4203 16779
rect 4203 16745 4212 16779
rect 4160 16736 4212 16745
rect 5356 16736 5408 16788
rect 6276 16736 6328 16788
rect 2688 16600 2740 16652
rect 2964 16600 3016 16652
rect 3424 16600 3476 16652
rect 4712 16668 4764 16720
rect 2780 16464 2832 16516
rect 4160 16600 4212 16652
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 4804 16600 4856 16652
rect 4896 16600 4948 16652
rect 5264 16600 5316 16652
rect 3884 16532 3936 16584
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 5908 16668 5960 16720
rect 6368 16668 6420 16720
rect 6736 16736 6788 16788
rect 9772 16736 9824 16788
rect 10416 16736 10468 16788
rect 10876 16736 10928 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 16304 16736 16356 16788
rect 19064 16736 19116 16788
rect 19156 16779 19208 16788
rect 19156 16745 19165 16779
rect 19165 16745 19199 16779
rect 19199 16745 19208 16779
rect 19156 16736 19208 16745
rect 19524 16736 19576 16788
rect 20996 16736 21048 16788
rect 22652 16779 22704 16788
rect 22652 16745 22661 16779
rect 22661 16745 22695 16779
rect 22695 16745 22704 16779
rect 22652 16736 22704 16745
rect 25780 16736 25832 16788
rect 29736 16736 29788 16788
rect 30104 16736 30156 16788
rect 30748 16736 30800 16788
rect 6552 16668 6604 16720
rect 11796 16668 11848 16720
rect 13728 16668 13780 16720
rect 14832 16668 14884 16720
rect 19708 16668 19760 16720
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 1952 16396 2004 16448
rect 4252 16396 4304 16448
rect 5356 16464 5408 16516
rect 6736 16600 6788 16652
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 11060 16600 11112 16652
rect 11152 16643 11204 16652
rect 11152 16609 11161 16643
rect 11161 16609 11195 16643
rect 11195 16609 11204 16643
rect 11152 16600 11204 16609
rect 11244 16600 11296 16652
rect 11612 16643 11664 16652
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 12440 16600 12492 16652
rect 17132 16600 17184 16652
rect 17684 16600 17736 16652
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 9772 16575 9824 16584
rect 9772 16541 9790 16575
rect 9790 16541 9824 16575
rect 9772 16532 9824 16541
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 10416 16532 10468 16584
rect 10508 16532 10560 16584
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 10968 16464 11020 16516
rect 11428 16507 11480 16516
rect 11428 16473 11437 16507
rect 11437 16473 11471 16507
rect 11471 16473 11480 16507
rect 11428 16464 11480 16473
rect 18144 16643 18196 16652
rect 18144 16609 18153 16643
rect 18153 16609 18187 16643
rect 18187 16609 18196 16643
rect 18144 16600 18196 16609
rect 18512 16600 18564 16652
rect 18972 16600 19024 16652
rect 19524 16600 19576 16652
rect 19892 16668 19944 16720
rect 22192 16668 22244 16720
rect 23664 16668 23716 16720
rect 24860 16668 24912 16720
rect 30012 16668 30064 16720
rect 30196 16711 30248 16720
rect 30196 16677 30214 16711
rect 30214 16677 30248 16711
rect 30196 16668 30248 16677
rect 20076 16643 20128 16652
rect 20076 16609 20085 16643
rect 20085 16609 20119 16643
rect 20119 16609 20128 16643
rect 20076 16600 20128 16609
rect 20352 16600 20404 16652
rect 21364 16600 21416 16652
rect 22928 16643 22980 16652
rect 22928 16609 22937 16643
rect 22937 16609 22971 16643
rect 22971 16609 22980 16643
rect 22928 16600 22980 16609
rect 23020 16643 23072 16652
rect 23020 16609 23029 16643
rect 23029 16609 23063 16643
rect 23063 16609 23072 16643
rect 23020 16600 23072 16609
rect 23204 16643 23256 16652
rect 23204 16609 23213 16643
rect 23213 16609 23247 16643
rect 23247 16609 23256 16643
rect 23204 16600 23256 16609
rect 23480 16600 23532 16652
rect 6000 16396 6052 16448
rect 17500 16439 17552 16448
rect 17500 16405 17509 16439
rect 17509 16405 17543 16439
rect 17543 16405 17552 16439
rect 17500 16396 17552 16405
rect 17684 16396 17736 16448
rect 19064 16464 19116 16516
rect 19432 16464 19484 16516
rect 19708 16464 19760 16516
rect 22468 16532 22520 16584
rect 24032 16643 24084 16652
rect 24032 16609 24041 16643
rect 24041 16609 24075 16643
rect 24075 16609 24084 16643
rect 24032 16600 24084 16609
rect 24124 16643 24176 16652
rect 24124 16609 24133 16643
rect 24133 16609 24167 16643
rect 24167 16609 24176 16643
rect 24124 16600 24176 16609
rect 25228 16600 25280 16652
rect 26700 16643 26752 16652
rect 26700 16609 26709 16643
rect 26709 16609 26743 16643
rect 26743 16609 26752 16643
rect 26700 16600 26752 16609
rect 27896 16600 27948 16652
rect 22560 16464 22612 16516
rect 20260 16396 20312 16448
rect 23388 16464 23440 16516
rect 24492 16464 24544 16516
rect 24768 16464 24820 16516
rect 28448 16532 28500 16584
rect 28632 16643 28684 16652
rect 28632 16609 28641 16643
rect 28641 16609 28675 16643
rect 28675 16609 28684 16643
rect 28632 16600 28684 16609
rect 28724 16643 28776 16652
rect 28724 16609 28733 16643
rect 28733 16609 28767 16643
rect 28767 16609 28776 16643
rect 28724 16600 28776 16609
rect 28816 16643 28868 16652
rect 28816 16609 28825 16643
rect 28825 16609 28859 16643
rect 28859 16609 28868 16643
rect 28816 16600 28868 16609
rect 28908 16600 28960 16652
rect 31208 16600 31260 16652
rect 27344 16464 27396 16516
rect 27620 16464 27672 16516
rect 25964 16396 26016 16448
rect 27528 16396 27580 16448
rect 29000 16396 29052 16448
rect 30288 16396 30340 16448
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 11436 16294 11488 16346
rect 11500 16294 11552 16346
rect 11564 16294 11616 16346
rect 11628 16294 11680 16346
rect 11692 16294 11744 16346
rect 19210 16294 19262 16346
rect 19274 16294 19326 16346
rect 19338 16294 19390 16346
rect 19402 16294 19454 16346
rect 19466 16294 19518 16346
rect 26984 16294 27036 16346
rect 27048 16294 27100 16346
rect 27112 16294 27164 16346
rect 27176 16294 27228 16346
rect 27240 16294 27292 16346
rect 4896 16192 4948 16244
rect 2688 16124 2740 16176
rect 4712 16124 4764 16176
rect 5172 16192 5224 16244
rect 9496 16192 9548 16244
rect 17224 16192 17276 16244
rect 18420 16235 18472 16244
rect 18420 16201 18429 16235
rect 18429 16201 18463 16235
rect 18463 16201 18472 16235
rect 18420 16192 18472 16201
rect 19064 16235 19116 16244
rect 19064 16201 19073 16235
rect 19073 16201 19107 16235
rect 19107 16201 19116 16235
rect 19064 16192 19116 16201
rect 19524 16192 19576 16244
rect 20168 16192 20220 16244
rect 20628 16192 20680 16244
rect 5816 16124 5868 16176
rect 8576 16124 8628 16176
rect 11060 16124 11112 16176
rect 17684 16124 17736 16176
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 1952 16031 2004 16040
rect 1952 15997 1986 16031
rect 1986 15997 2004 16031
rect 1952 15988 2004 15997
rect 4160 15988 4212 16040
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 6552 15988 6604 16040
rect 8024 16031 8076 16040
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 9312 16031 9364 16040
rect 9312 15997 9321 16031
rect 9321 15997 9355 16031
rect 9355 15997 9364 16031
rect 9312 15988 9364 15997
rect 9956 16056 10008 16108
rect 10232 16056 10284 16108
rect 9496 16031 9548 16040
rect 9496 15997 9505 16031
rect 9505 15997 9539 16031
rect 9539 15997 9548 16031
rect 9496 15988 9548 15997
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 9772 15988 9824 16040
rect 10968 15988 11020 16040
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 5540 15920 5592 15972
rect 5724 15920 5776 15972
rect 6644 15963 6696 15972
rect 6644 15929 6653 15963
rect 6653 15929 6687 15963
rect 6687 15929 6696 15963
rect 6644 15920 6696 15929
rect 13268 15988 13320 16040
rect 19524 16099 19576 16108
rect 19524 16065 19533 16099
rect 19533 16065 19567 16099
rect 19567 16065 19576 16099
rect 19524 16056 19576 16065
rect 20352 16124 20404 16176
rect 21088 16124 21140 16176
rect 19708 16056 19760 16108
rect 20720 16056 20772 16108
rect 14004 16031 14056 16040
rect 14004 15997 14013 16031
rect 14013 15997 14047 16031
rect 14047 15997 14056 16031
rect 14004 15988 14056 15997
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 17592 15988 17644 16040
rect 17776 16031 17828 16040
rect 17776 15997 17785 16031
rect 17785 15997 17819 16031
rect 17819 15997 17828 16031
rect 17776 15988 17828 15997
rect 17868 15988 17920 16040
rect 19892 16031 19944 16040
rect 19892 15997 19901 16031
rect 19901 15997 19935 16031
rect 19935 15997 19944 16031
rect 19892 15988 19944 15997
rect 22284 16192 22336 16244
rect 23388 16192 23440 16244
rect 25136 16192 25188 16244
rect 25504 16192 25556 16244
rect 29184 16192 29236 16244
rect 21824 16124 21876 16176
rect 24124 16124 24176 16176
rect 26148 16124 26200 16176
rect 22008 16031 22060 16040
rect 22008 15997 22017 16031
rect 22017 15997 22051 16031
rect 22051 15997 22060 16031
rect 22008 15988 22060 15997
rect 22100 15988 22152 16040
rect 14924 15920 14976 15972
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 7288 15852 7340 15904
rect 8116 15895 8168 15904
rect 8116 15861 8125 15895
rect 8125 15861 8159 15895
rect 8159 15861 8168 15895
rect 8116 15852 8168 15861
rect 9036 15895 9088 15904
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 9312 15852 9364 15904
rect 10324 15852 10376 15904
rect 11888 15852 11940 15904
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 17224 15895 17276 15904
rect 17224 15861 17233 15895
rect 17233 15861 17267 15895
rect 17267 15861 17276 15895
rect 17224 15852 17276 15861
rect 17776 15852 17828 15904
rect 18144 15963 18196 15972
rect 18144 15929 18153 15963
rect 18153 15929 18187 15963
rect 18187 15929 18196 15963
rect 18144 15920 18196 15929
rect 20076 15920 20128 15972
rect 22560 15988 22612 16040
rect 22652 15988 22704 16040
rect 23664 15988 23716 16040
rect 24768 15988 24820 16040
rect 25228 16056 25280 16108
rect 18420 15852 18472 15904
rect 18696 15852 18748 15904
rect 21272 15852 21324 15904
rect 21732 15895 21784 15904
rect 21732 15861 21741 15895
rect 21741 15861 21775 15895
rect 21775 15861 21784 15895
rect 21732 15852 21784 15861
rect 22468 15920 22520 15972
rect 23480 15920 23532 15972
rect 24952 15920 25004 15972
rect 22376 15852 22428 15904
rect 22928 15895 22980 15904
rect 22928 15861 22937 15895
rect 22937 15861 22971 15895
rect 22971 15861 22980 15895
rect 22928 15852 22980 15861
rect 23388 15852 23440 15904
rect 25412 15920 25464 15972
rect 25780 16031 25832 16040
rect 25780 15997 25789 16031
rect 25789 15997 25823 16031
rect 25823 15997 25832 16031
rect 25780 15988 25832 15997
rect 26056 16031 26108 16040
rect 26056 15997 26065 16031
rect 26065 15997 26099 16031
rect 26099 15997 26108 16031
rect 26056 15988 26108 15997
rect 26700 15920 26752 15972
rect 27344 15920 27396 15972
rect 26240 15852 26292 15904
rect 27620 16031 27672 16040
rect 27620 15997 27629 16031
rect 27629 15997 27663 16031
rect 27663 15997 27672 16031
rect 27620 15988 27672 15997
rect 27804 16031 27856 16040
rect 27804 15997 27813 16031
rect 27813 15997 27847 16031
rect 27847 15997 27856 16031
rect 27804 15988 27856 15997
rect 28172 16056 28224 16108
rect 29552 16099 29604 16108
rect 29552 16065 29561 16099
rect 29561 16065 29595 16099
rect 29595 16065 29604 16099
rect 29552 16056 29604 16065
rect 28632 15988 28684 16040
rect 28540 15920 28592 15972
rect 30012 16031 30064 16040
rect 30012 15997 30021 16031
rect 30021 15997 30055 16031
rect 30055 15997 30064 16031
rect 30012 15988 30064 15997
rect 28080 15852 28132 15904
rect 28172 15895 28224 15904
rect 28172 15861 28181 15895
rect 28181 15861 28215 15895
rect 28215 15861 28224 15895
rect 28172 15852 28224 15861
rect 28908 15852 28960 15904
rect 29828 15852 29880 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 12096 15750 12148 15802
rect 12160 15750 12212 15802
rect 12224 15750 12276 15802
rect 12288 15750 12340 15802
rect 12352 15750 12404 15802
rect 19870 15750 19922 15802
rect 19934 15750 19986 15802
rect 19998 15750 20050 15802
rect 20062 15750 20114 15802
rect 20126 15750 20178 15802
rect 27644 15750 27696 15802
rect 27708 15750 27760 15802
rect 27772 15750 27824 15802
rect 27836 15750 27888 15802
rect 27900 15750 27952 15802
rect 2688 15691 2740 15700
rect 2688 15657 2697 15691
rect 2697 15657 2731 15691
rect 2731 15657 2740 15691
rect 2688 15648 2740 15657
rect 6000 15648 6052 15700
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 9772 15648 9824 15700
rect 10416 15648 10468 15700
rect 1400 15580 1452 15632
rect 1308 15555 1360 15564
rect 1308 15521 1317 15555
rect 1317 15521 1351 15555
rect 1351 15521 1360 15555
rect 1308 15512 1360 15521
rect 5540 15580 5592 15632
rect 5724 15580 5776 15632
rect 6644 15580 6696 15632
rect 11152 15648 11204 15700
rect 14004 15648 14056 15700
rect 14188 15648 14240 15700
rect 17776 15648 17828 15700
rect 12440 15580 12492 15632
rect 13084 15580 13136 15632
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 8116 15512 8168 15564
rect 9036 15555 9088 15564
rect 9036 15521 9070 15555
rect 9070 15521 9088 15555
rect 9036 15512 9088 15521
rect 9864 15512 9916 15564
rect 3056 15444 3108 15496
rect 4068 15444 4120 15496
rect 7104 15444 7156 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10876 15512 10928 15564
rect 11060 15512 11112 15564
rect 11888 15512 11940 15564
rect 13544 15512 13596 15564
rect 15568 15580 15620 15632
rect 17500 15623 17552 15632
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 14004 15555 14056 15564
rect 14004 15521 14013 15555
rect 14013 15521 14047 15555
rect 14047 15521 14056 15555
rect 14004 15512 14056 15521
rect 14096 15555 14148 15564
rect 14096 15521 14105 15555
rect 14105 15521 14139 15555
rect 14139 15521 14148 15555
rect 14096 15512 14148 15521
rect 12532 15444 12584 15496
rect 13728 15444 13780 15496
rect 14832 15555 14884 15564
rect 14832 15521 14841 15555
rect 14841 15521 14875 15555
rect 14875 15521 14884 15555
rect 14832 15512 14884 15521
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 16764 15555 16816 15564
rect 16764 15521 16772 15555
rect 16772 15521 16806 15555
rect 16806 15521 16816 15555
rect 16764 15512 16816 15521
rect 15752 15444 15804 15496
rect 11244 15376 11296 15428
rect 14096 15376 14148 15428
rect 1400 15351 1452 15360
rect 1400 15317 1409 15351
rect 1409 15317 1443 15351
rect 1443 15317 1452 15351
rect 1400 15308 1452 15317
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 10416 15351 10468 15360
rect 10416 15317 10425 15351
rect 10425 15317 10459 15351
rect 10459 15317 10468 15351
rect 10416 15308 10468 15317
rect 10968 15308 11020 15360
rect 14372 15308 14424 15360
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 17040 15512 17092 15564
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 17500 15589 17534 15623
rect 17534 15589 17552 15623
rect 17500 15580 17552 15589
rect 18328 15580 18380 15632
rect 18512 15580 18564 15632
rect 20720 15648 20772 15700
rect 21364 15648 21416 15700
rect 18788 15580 18840 15632
rect 19616 15580 19668 15632
rect 20260 15580 20312 15632
rect 21732 15648 21784 15700
rect 22100 15648 22152 15700
rect 22468 15648 22520 15700
rect 24308 15648 24360 15700
rect 18052 15512 18104 15564
rect 18236 15512 18288 15564
rect 19708 15555 19760 15564
rect 19708 15521 19717 15555
rect 19717 15521 19751 15555
rect 19751 15521 19760 15555
rect 19708 15512 19760 15521
rect 20444 15555 20496 15564
rect 20444 15521 20453 15555
rect 20453 15521 20487 15555
rect 20487 15521 20496 15555
rect 20444 15512 20496 15521
rect 20996 15512 21048 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 22284 15580 22336 15632
rect 18328 15376 18380 15428
rect 19984 15376 20036 15428
rect 17960 15308 18012 15360
rect 19708 15308 19760 15360
rect 21088 15444 21140 15496
rect 20904 15376 20956 15428
rect 21824 15444 21876 15496
rect 23940 15555 23992 15564
rect 23940 15521 23949 15555
rect 23949 15521 23983 15555
rect 23983 15521 23992 15555
rect 27436 15580 27488 15632
rect 27804 15580 27856 15632
rect 23940 15512 23992 15521
rect 22284 15444 22336 15496
rect 23204 15444 23256 15496
rect 24400 15512 24452 15564
rect 24952 15512 25004 15564
rect 24584 15444 24636 15496
rect 26700 15512 26752 15564
rect 26792 15512 26844 15564
rect 27528 15512 27580 15564
rect 27896 15555 27948 15564
rect 27896 15521 27905 15555
rect 27905 15521 27939 15555
rect 27939 15521 27948 15555
rect 27896 15512 27948 15521
rect 28172 15512 28224 15564
rect 28908 15648 28960 15700
rect 29000 15648 29052 15700
rect 30288 15648 30340 15700
rect 29276 15512 29328 15564
rect 29828 15555 29880 15564
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 30748 15512 30800 15564
rect 22652 15376 22704 15428
rect 27804 15376 27856 15428
rect 27988 15376 28040 15428
rect 23296 15308 23348 15360
rect 24032 15308 24084 15360
rect 24860 15308 24912 15360
rect 28448 15308 28500 15360
rect 29184 15308 29236 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 11436 15206 11488 15258
rect 11500 15206 11552 15258
rect 11564 15206 11616 15258
rect 11628 15206 11680 15258
rect 11692 15206 11744 15258
rect 19210 15206 19262 15258
rect 19274 15206 19326 15258
rect 19338 15206 19390 15258
rect 19402 15206 19454 15258
rect 19466 15206 19518 15258
rect 26984 15206 27036 15258
rect 27048 15206 27100 15258
rect 27112 15206 27164 15258
rect 27176 15206 27228 15258
rect 27240 15206 27292 15258
rect 9864 15104 9916 15156
rect 9956 15104 10008 15156
rect 11612 15104 11664 15156
rect 5632 15036 5684 15088
rect 1400 14968 1452 15020
rect 3332 14968 3384 15020
rect 1308 14943 1360 14952
rect 1308 14909 1317 14943
rect 1317 14909 1351 14943
rect 1351 14909 1360 14943
rect 1308 14900 1360 14909
rect 3516 14900 3568 14952
rect 3976 14943 4028 14952
rect 3976 14909 3985 14943
rect 3985 14909 4019 14943
rect 4019 14909 4028 14943
rect 3976 14900 4028 14909
rect 4804 14968 4856 15020
rect 1492 14764 1544 14816
rect 4160 14832 4212 14884
rect 4620 14900 4672 14952
rect 4896 14900 4948 14952
rect 5540 14900 5592 14952
rect 5172 14832 5224 14884
rect 6828 14875 6880 14884
rect 6828 14841 6846 14875
rect 6846 14841 6880 14875
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 9956 14968 10008 15020
rect 13728 15104 13780 15156
rect 14004 15147 14056 15156
rect 14004 15113 14013 15147
rect 14013 15113 14047 15147
rect 14047 15113 14056 15147
rect 14004 15104 14056 15113
rect 16672 15147 16724 15156
rect 16672 15113 16681 15147
rect 16681 15113 16715 15147
rect 16715 15113 16724 15147
rect 16672 15104 16724 15113
rect 16948 15104 17000 15156
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 9496 14943 9548 14952
rect 9496 14909 9505 14943
rect 9505 14909 9539 14943
rect 9539 14909 9548 14943
rect 9496 14900 9548 14909
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 11060 14900 11112 14952
rect 11612 14943 11664 14952
rect 11612 14909 11621 14943
rect 11621 14909 11655 14943
rect 11655 14909 11664 14943
rect 11612 14900 11664 14909
rect 11796 14900 11848 14952
rect 6828 14832 6880 14841
rect 4712 14764 4764 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 6552 14764 6604 14816
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 9680 14764 9732 14816
rect 11980 14900 12032 14952
rect 13452 14968 13504 15020
rect 13728 14968 13780 15020
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 18144 15104 18196 15156
rect 19248 15104 19300 15156
rect 19616 15104 19668 15156
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 13268 14900 13320 14952
rect 13636 14943 13688 14952
rect 13636 14909 13645 14943
rect 13645 14909 13679 14943
rect 13679 14909 13688 14943
rect 14372 14943 14424 14952
rect 13636 14900 13688 14909
rect 13176 14832 13228 14884
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 13820 14875 13872 14884
rect 13820 14841 13829 14875
rect 13829 14841 13863 14875
rect 13863 14841 13872 14875
rect 13820 14832 13872 14841
rect 14372 14909 14406 14943
rect 14406 14909 14424 14943
rect 14372 14900 14424 14909
rect 14464 14832 14516 14884
rect 14188 14764 14240 14816
rect 16948 14900 17000 14952
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 18144 14968 18196 15020
rect 18972 15036 19024 15088
rect 20720 15104 20772 15156
rect 21364 15147 21416 15156
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 23204 15104 23256 15156
rect 23664 15104 23716 15156
rect 25412 15104 25464 15156
rect 25504 15104 25556 15156
rect 27896 15104 27948 15156
rect 15752 14807 15804 14816
rect 15752 14773 15761 14807
rect 15761 14773 15795 14807
rect 15795 14773 15804 14807
rect 15752 14764 15804 14773
rect 17500 14832 17552 14884
rect 18604 14900 18656 14952
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 18788 14943 18840 14952
rect 18788 14909 18798 14943
rect 18798 14909 18832 14943
rect 18832 14909 18840 14943
rect 18788 14900 18840 14909
rect 18972 14900 19024 14952
rect 19984 15036 20036 15088
rect 23480 15036 23532 15088
rect 19248 14968 19300 15020
rect 19340 14900 19392 14952
rect 22744 14968 22796 15020
rect 21088 14943 21140 14952
rect 21088 14909 21097 14943
rect 21097 14909 21131 14943
rect 21131 14909 21140 14943
rect 21088 14900 21140 14909
rect 21364 14943 21416 14952
rect 21364 14909 21373 14943
rect 21373 14909 21407 14943
rect 21407 14909 21416 14943
rect 21364 14900 21416 14909
rect 16948 14764 17000 14816
rect 17684 14764 17736 14816
rect 17960 14764 18012 14816
rect 19156 14764 19208 14816
rect 20628 14832 20680 14884
rect 20996 14832 21048 14884
rect 22100 14900 22152 14952
rect 23664 14943 23716 14952
rect 23664 14909 23673 14943
rect 23673 14909 23707 14943
rect 23707 14909 23716 14943
rect 23664 14900 23716 14909
rect 24032 14943 24084 14952
rect 24032 14909 24041 14943
rect 24041 14909 24075 14943
rect 24075 14909 24084 14943
rect 24032 14900 24084 14909
rect 24216 14900 24268 14952
rect 25596 15036 25648 15088
rect 26240 15036 26292 15088
rect 28724 15104 28776 15156
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 20720 14764 20772 14816
rect 23480 14875 23532 14884
rect 23480 14841 23489 14875
rect 23489 14841 23523 14875
rect 23523 14841 23532 14875
rect 23480 14832 23532 14841
rect 23756 14832 23808 14884
rect 21548 14764 21600 14816
rect 22652 14764 22704 14816
rect 23388 14764 23440 14816
rect 23572 14764 23624 14816
rect 24952 14943 25004 14952
rect 24952 14909 24961 14943
rect 24961 14909 24995 14943
rect 24995 14909 25004 14943
rect 24952 14900 25004 14909
rect 25504 14968 25556 15020
rect 25228 14900 25280 14952
rect 25044 14764 25096 14816
rect 25320 14807 25372 14816
rect 25320 14773 25329 14807
rect 25329 14773 25363 14807
rect 25363 14773 25372 14807
rect 25320 14764 25372 14773
rect 25504 14764 25556 14816
rect 25872 14943 25924 14952
rect 25872 14909 25881 14943
rect 25881 14909 25915 14943
rect 25915 14909 25924 14943
rect 25872 14900 25924 14909
rect 26056 14943 26108 14952
rect 26056 14909 26065 14943
rect 26065 14909 26099 14943
rect 26099 14909 26108 14943
rect 26056 14900 26108 14909
rect 26700 14943 26752 14952
rect 26700 14909 26709 14943
rect 26709 14909 26743 14943
rect 26743 14909 26752 14943
rect 28172 14968 28224 15020
rect 26700 14900 26752 14909
rect 27436 14900 27488 14952
rect 27528 14943 27580 14952
rect 27528 14909 27537 14943
rect 27537 14909 27571 14943
rect 27571 14909 27580 14943
rect 27528 14900 27580 14909
rect 28264 14900 28316 14952
rect 29000 15036 29052 15088
rect 28540 14943 28592 14952
rect 28540 14909 28549 14943
rect 28549 14909 28583 14943
rect 28583 14909 28592 14943
rect 28540 14900 28592 14909
rect 28816 14943 28868 14952
rect 28816 14909 28825 14943
rect 28825 14909 28859 14943
rect 28859 14909 28868 14943
rect 28816 14900 28868 14909
rect 25964 14764 26016 14816
rect 29092 14900 29144 14952
rect 29460 14968 29512 15020
rect 29552 14900 29604 14952
rect 29736 14943 29788 14952
rect 29736 14909 29745 14943
rect 29745 14909 29779 14943
rect 29779 14909 29788 14943
rect 29736 14900 29788 14909
rect 30748 14900 30800 14952
rect 26608 14764 26660 14816
rect 27436 14764 27488 14816
rect 28908 14764 28960 14816
rect 29644 14807 29696 14816
rect 29644 14773 29653 14807
rect 29653 14773 29687 14807
rect 29687 14773 29696 14807
rect 29644 14764 29696 14773
rect 30104 14764 30156 14816
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 12096 14662 12148 14714
rect 12160 14662 12212 14714
rect 12224 14662 12276 14714
rect 12288 14662 12340 14714
rect 12352 14662 12404 14714
rect 19870 14662 19922 14714
rect 19934 14662 19986 14714
rect 19998 14662 20050 14714
rect 20062 14662 20114 14714
rect 20126 14662 20178 14714
rect 27644 14662 27696 14714
rect 27708 14662 27760 14714
rect 27772 14662 27824 14714
rect 27836 14662 27888 14714
rect 27900 14662 27952 14714
rect 4804 14560 4856 14612
rect 5356 14560 5408 14612
rect 1584 14492 1636 14544
rect 2964 14492 3016 14544
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2780 14424 2832 14476
rect 3424 14492 3476 14544
rect 3976 14492 4028 14544
rect 4068 14492 4120 14544
rect 3516 14356 3568 14408
rect 4068 14356 4120 14408
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 7104 14424 7156 14476
rect 6552 14356 6604 14408
rect 9036 14492 9088 14544
rect 11612 14492 11664 14544
rect 12900 14560 12952 14612
rect 14832 14560 14884 14612
rect 13360 14492 13412 14544
rect 17592 14560 17644 14612
rect 17684 14560 17736 14612
rect 8852 14424 8904 14476
rect 3056 14331 3108 14340
rect 3056 14297 3065 14331
rect 3065 14297 3099 14331
rect 3099 14297 3108 14331
rect 3056 14288 3108 14297
rect 4988 14288 5040 14340
rect 5356 14288 5408 14340
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 11796 14424 11848 14476
rect 12624 14424 12676 14476
rect 12992 14424 13044 14476
rect 13636 14467 13688 14476
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 13820 14424 13872 14476
rect 14556 14424 14608 14476
rect 10508 14288 10560 14340
rect 13084 14356 13136 14408
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 12532 14331 12584 14340
rect 12532 14297 12541 14331
rect 12541 14297 12575 14331
rect 12575 14297 12584 14331
rect 12532 14288 12584 14297
rect 15752 14424 15804 14476
rect 16580 14356 16632 14408
rect 17224 14424 17276 14476
rect 17500 14424 17552 14476
rect 17960 14424 18012 14476
rect 19708 14560 19760 14612
rect 18512 14492 18564 14544
rect 19616 14492 19668 14544
rect 19892 14492 19944 14544
rect 20536 14492 20588 14544
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 18236 14424 18288 14476
rect 18604 14467 18656 14476
rect 18604 14433 18613 14467
rect 18613 14433 18647 14467
rect 18647 14433 18656 14467
rect 18604 14424 18656 14433
rect 18512 14356 18564 14408
rect 20260 14467 20312 14476
rect 20260 14433 20269 14467
rect 20269 14433 20303 14467
rect 20303 14433 20312 14467
rect 20260 14424 20312 14433
rect 21548 14560 21600 14612
rect 21088 14492 21140 14544
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 21364 14424 21416 14476
rect 22744 14535 22796 14544
rect 22744 14501 22753 14535
rect 22753 14501 22787 14535
rect 22787 14501 22796 14535
rect 22744 14492 22796 14501
rect 23480 14560 23532 14612
rect 21916 14467 21968 14476
rect 21916 14433 21925 14467
rect 21925 14433 21959 14467
rect 21959 14433 21968 14467
rect 21916 14424 21968 14433
rect 22100 14424 22152 14476
rect 22284 14424 22336 14476
rect 22468 14467 22520 14476
rect 22468 14433 22477 14467
rect 22477 14433 22511 14467
rect 22511 14433 22520 14467
rect 22468 14424 22520 14433
rect 22652 14467 22704 14476
rect 22652 14433 22661 14467
rect 22661 14433 22695 14467
rect 22695 14433 22704 14467
rect 22652 14424 22704 14433
rect 24032 14560 24084 14612
rect 26700 14560 26752 14612
rect 27528 14560 27580 14612
rect 28908 14560 28960 14612
rect 29552 14603 29604 14612
rect 29552 14569 29561 14603
rect 29561 14569 29595 14603
rect 29595 14569 29604 14603
rect 29552 14560 29604 14569
rect 25320 14492 25372 14544
rect 23296 14424 23348 14476
rect 23388 14467 23440 14476
rect 23388 14433 23397 14467
rect 23397 14433 23431 14467
rect 23431 14433 23440 14467
rect 23388 14424 23440 14433
rect 24124 14424 24176 14476
rect 24308 14424 24360 14476
rect 24768 14424 24820 14476
rect 24860 14467 24912 14476
rect 24860 14433 24869 14467
rect 24869 14433 24903 14467
rect 24903 14433 24912 14467
rect 24860 14424 24912 14433
rect 29644 14492 29696 14544
rect 17408 14288 17460 14340
rect 26148 14356 26200 14408
rect 27436 14356 27488 14408
rect 27988 14467 28040 14476
rect 27988 14433 27997 14467
rect 27997 14433 28031 14467
rect 28031 14433 28040 14467
rect 27988 14424 28040 14433
rect 21916 14288 21968 14340
rect 26792 14288 26844 14340
rect 28448 14467 28500 14476
rect 28448 14433 28457 14467
rect 28457 14433 28491 14467
rect 28491 14433 28500 14467
rect 28448 14424 28500 14433
rect 29184 14424 29236 14476
rect 29828 14424 29880 14476
rect 30288 14467 30340 14476
rect 30288 14433 30297 14467
rect 30297 14433 30331 14467
rect 30331 14433 30340 14467
rect 30288 14424 30340 14433
rect 30472 14467 30524 14476
rect 30472 14433 30481 14467
rect 30481 14433 30515 14467
rect 30515 14433 30524 14467
rect 30472 14424 30524 14433
rect 30564 14467 30616 14476
rect 30564 14433 30573 14467
rect 30573 14433 30607 14467
rect 30607 14433 30616 14467
rect 30564 14424 30616 14433
rect 30932 14467 30984 14476
rect 30932 14433 30941 14467
rect 30941 14433 30975 14467
rect 30975 14433 30984 14467
rect 30932 14424 30984 14433
rect 29276 14399 29328 14408
rect 29276 14365 29285 14399
rect 29285 14365 29319 14399
rect 29319 14365 29328 14399
rect 29276 14356 29328 14365
rect 5080 14263 5132 14272
rect 5080 14229 5089 14263
rect 5089 14229 5123 14263
rect 5123 14229 5132 14263
rect 5080 14220 5132 14229
rect 5908 14263 5960 14272
rect 5908 14229 5917 14263
rect 5917 14229 5951 14263
rect 5951 14229 5960 14263
rect 5908 14220 5960 14229
rect 10968 14263 11020 14272
rect 10968 14229 10977 14263
rect 10977 14229 11011 14263
rect 11011 14229 11020 14263
rect 10968 14220 11020 14229
rect 17040 14220 17092 14272
rect 18604 14220 18656 14272
rect 20444 14263 20496 14272
rect 20444 14229 20453 14263
rect 20453 14229 20487 14263
rect 20487 14229 20496 14263
rect 20444 14220 20496 14229
rect 20904 14220 20956 14272
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 21732 14263 21784 14272
rect 21732 14229 21741 14263
rect 21741 14229 21775 14263
rect 21775 14229 21784 14263
rect 21732 14220 21784 14229
rect 24860 14220 24912 14272
rect 26148 14220 26200 14272
rect 26700 14220 26752 14272
rect 27988 14220 28040 14272
rect 28632 14220 28684 14272
rect 29000 14220 29052 14272
rect 29092 14220 29144 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 11436 14118 11488 14170
rect 11500 14118 11552 14170
rect 11564 14118 11616 14170
rect 11628 14118 11680 14170
rect 11692 14118 11744 14170
rect 19210 14118 19262 14170
rect 19274 14118 19326 14170
rect 19338 14118 19390 14170
rect 19402 14118 19454 14170
rect 19466 14118 19518 14170
rect 26984 14118 27036 14170
rect 27048 14118 27100 14170
rect 27112 14118 27164 14170
rect 27176 14118 27228 14170
rect 27240 14118 27292 14170
rect 3056 13948 3108 14000
rect 4068 13880 4120 13932
rect 1308 13812 1360 13864
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 3884 13855 3936 13864
rect 3884 13821 3893 13855
rect 3893 13821 3927 13855
rect 3927 13821 3936 13855
rect 3884 13812 3936 13821
rect 6276 14016 6328 14068
rect 6368 14016 6420 14068
rect 5540 13948 5592 14000
rect 9496 14016 9548 14068
rect 10600 14016 10652 14068
rect 12532 14016 12584 14068
rect 13728 14016 13780 14068
rect 15016 14059 15068 14068
rect 15016 14025 15025 14059
rect 15025 14025 15059 14059
rect 15059 14025 15068 14059
rect 15016 14016 15068 14025
rect 11244 13948 11296 14000
rect 14924 13948 14976 14000
rect 16304 14016 16356 14068
rect 16488 13948 16540 14000
rect 17500 13991 17552 14000
rect 17500 13957 17509 13991
rect 17509 13957 17543 13991
rect 17543 13957 17552 13991
rect 17500 13948 17552 13957
rect 17868 13948 17920 14000
rect 18144 14059 18196 14068
rect 18144 14025 18153 14059
rect 18153 14025 18187 14059
rect 18187 14025 18196 14059
rect 18144 14016 18196 14025
rect 21272 14016 21324 14068
rect 7104 13880 7156 13932
rect 5080 13812 5132 13864
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 5908 13855 5960 13864
rect 5908 13821 5942 13855
rect 5942 13821 5960 13855
rect 5908 13812 5960 13821
rect 6276 13812 6328 13864
rect 9496 13880 9548 13932
rect 8944 13812 8996 13864
rect 9312 13812 9364 13864
rect 9956 13812 10008 13864
rect 10968 13880 11020 13932
rect 14648 13880 14700 13932
rect 10600 13812 10652 13864
rect 5448 13744 5500 13796
rect 6736 13744 6788 13796
rect 9496 13787 9548 13796
rect 9496 13753 9505 13787
rect 9505 13753 9539 13787
rect 9539 13753 9548 13787
rect 9496 13744 9548 13753
rect 10048 13744 10100 13796
rect 11152 13812 11204 13864
rect 11980 13812 12032 13864
rect 14740 13812 14792 13864
rect 17776 13880 17828 13932
rect 16304 13855 16356 13864
rect 16304 13821 16313 13855
rect 16313 13821 16347 13855
rect 16347 13821 16356 13855
rect 16304 13812 16356 13821
rect 16488 13855 16540 13864
rect 16488 13821 16497 13855
rect 16497 13821 16531 13855
rect 16531 13821 16540 13855
rect 16488 13812 16540 13821
rect 11888 13744 11940 13796
rect 15476 13787 15528 13796
rect 15476 13753 15485 13787
rect 15485 13753 15519 13787
rect 15519 13753 15528 13787
rect 15476 13744 15528 13753
rect 17040 13744 17092 13796
rect 17592 13812 17644 13864
rect 19432 13880 19484 13932
rect 19892 13948 19944 14000
rect 20536 13991 20588 14000
rect 20536 13957 20545 13991
rect 20545 13957 20579 13991
rect 20579 13957 20588 13991
rect 20536 13948 20588 13957
rect 21088 13948 21140 14000
rect 22468 14016 22520 14068
rect 23756 14016 23808 14068
rect 25228 14059 25280 14068
rect 25228 14025 25237 14059
rect 25237 14025 25271 14059
rect 25271 14025 25280 14059
rect 25228 14016 25280 14025
rect 25688 14016 25740 14068
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 17868 13744 17920 13796
rect 20260 13812 20312 13864
rect 22376 13855 22428 13864
rect 22376 13821 22385 13855
rect 22385 13821 22419 13855
rect 22419 13821 22428 13855
rect 22376 13812 22428 13821
rect 2320 13676 2372 13728
rect 2964 13719 3016 13728
rect 2964 13685 2973 13719
rect 2973 13685 3007 13719
rect 3007 13685 3016 13719
rect 2964 13676 3016 13685
rect 5172 13676 5224 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7656 13719 7708 13728
rect 7656 13685 7665 13719
rect 7665 13685 7699 13719
rect 7699 13685 7708 13719
rect 7656 13676 7708 13685
rect 10324 13676 10376 13728
rect 11060 13676 11112 13728
rect 16764 13676 16816 13728
rect 17316 13676 17368 13728
rect 19616 13744 19668 13796
rect 19984 13744 20036 13796
rect 20996 13744 21048 13796
rect 23388 13855 23440 13864
rect 23388 13821 23397 13855
rect 23397 13821 23431 13855
rect 23431 13821 23440 13855
rect 23388 13812 23440 13821
rect 23572 13812 23624 13864
rect 23756 13812 23808 13864
rect 23848 13855 23900 13864
rect 23848 13821 23857 13855
rect 23857 13821 23891 13855
rect 23891 13821 23900 13855
rect 23848 13812 23900 13821
rect 25412 13880 25464 13932
rect 25688 13855 25740 13864
rect 25688 13821 25697 13855
rect 25697 13821 25731 13855
rect 25731 13821 25740 13855
rect 25688 13812 25740 13821
rect 26148 13880 26200 13932
rect 26792 13948 26844 14000
rect 24308 13744 24360 13796
rect 18328 13719 18380 13728
rect 18328 13685 18337 13719
rect 18337 13685 18371 13719
rect 18371 13685 18380 13719
rect 18328 13676 18380 13685
rect 20260 13719 20312 13728
rect 20260 13685 20269 13719
rect 20269 13685 20303 13719
rect 20303 13685 20312 13719
rect 20260 13676 20312 13685
rect 20812 13676 20864 13728
rect 26516 13744 26568 13796
rect 26884 13855 26936 13864
rect 26884 13821 26893 13855
rect 26893 13821 26927 13855
rect 26927 13821 26936 13855
rect 26884 13812 26936 13821
rect 26976 13855 27028 13864
rect 26976 13821 26985 13855
rect 26985 13821 27019 13855
rect 27019 13821 27028 13855
rect 26976 13812 27028 13821
rect 28172 14016 28224 14068
rect 27620 13880 27672 13932
rect 27436 13744 27488 13796
rect 29368 13948 29420 14000
rect 29828 14059 29880 14068
rect 29828 14025 29837 14059
rect 29837 14025 29871 14059
rect 29871 14025 29880 14059
rect 29828 14016 29880 14025
rect 30472 14016 30524 14068
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 30104 13855 30156 13864
rect 30104 13821 30113 13855
rect 30113 13821 30147 13855
rect 30147 13821 30156 13855
rect 30104 13812 30156 13821
rect 25320 13719 25372 13728
rect 25320 13685 25329 13719
rect 25329 13685 25363 13719
rect 25363 13685 25372 13719
rect 25320 13676 25372 13685
rect 25872 13676 25924 13728
rect 28724 13676 28776 13728
rect 29368 13719 29420 13728
rect 29368 13685 29377 13719
rect 29377 13685 29411 13719
rect 29411 13685 29420 13719
rect 29368 13676 29420 13685
rect 30748 13676 30800 13728
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 12096 13574 12148 13626
rect 12160 13574 12212 13626
rect 12224 13574 12276 13626
rect 12288 13574 12340 13626
rect 12352 13574 12404 13626
rect 19870 13574 19922 13626
rect 19934 13574 19986 13626
rect 19998 13574 20050 13626
rect 20062 13574 20114 13626
rect 20126 13574 20178 13626
rect 27644 13574 27696 13626
rect 27708 13574 27760 13626
rect 27772 13574 27824 13626
rect 27836 13574 27888 13626
rect 27900 13574 27952 13626
rect 2872 13472 2924 13524
rect 3516 13472 3568 13524
rect 4896 13472 4948 13524
rect 7656 13472 7708 13524
rect 2964 13404 3016 13456
rect 3608 13404 3660 13456
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 3424 13336 3476 13388
rect 8208 13404 8260 13456
rect 11888 13472 11940 13524
rect 12900 13515 12952 13524
rect 12900 13481 12909 13515
rect 12909 13481 12943 13515
rect 12943 13481 12952 13515
rect 12900 13472 12952 13481
rect 13636 13472 13688 13524
rect 3424 13132 3476 13184
rect 3884 13268 3936 13320
rect 5448 13379 5500 13388
rect 5448 13345 5457 13379
rect 5457 13345 5491 13379
rect 5491 13345 5500 13379
rect 5448 13336 5500 13345
rect 7196 13336 7248 13388
rect 9312 13379 9364 13388
rect 9312 13345 9321 13379
rect 9321 13345 9355 13379
rect 9355 13345 9364 13379
rect 9312 13336 9364 13345
rect 9404 13268 9456 13320
rect 7104 13200 7156 13252
rect 9680 13336 9732 13388
rect 10048 13336 10100 13388
rect 13728 13404 13780 13456
rect 16672 13472 16724 13524
rect 20444 13472 20496 13524
rect 23848 13472 23900 13524
rect 28724 13515 28776 13524
rect 28724 13481 28733 13515
rect 28733 13481 28767 13515
rect 28767 13481 28776 13515
rect 28724 13472 28776 13481
rect 29184 13472 29236 13524
rect 8300 13132 8352 13184
rect 8852 13132 8904 13184
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 11060 13336 11112 13388
rect 11796 13336 11848 13388
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 13452 13336 13504 13388
rect 14740 13404 14792 13456
rect 24308 13447 24360 13456
rect 24308 13413 24317 13447
rect 24317 13413 24351 13447
rect 24351 13413 24360 13447
rect 24308 13404 24360 13413
rect 25044 13447 25096 13456
rect 25044 13413 25053 13447
rect 25053 13413 25087 13447
rect 25087 13413 25096 13447
rect 25044 13404 25096 13413
rect 25412 13404 25464 13456
rect 25872 13447 25924 13456
rect 25872 13413 25881 13447
rect 25881 13413 25915 13447
rect 25915 13413 25924 13447
rect 25872 13404 25924 13413
rect 26056 13447 26108 13456
rect 26056 13413 26065 13447
rect 26065 13413 26099 13447
rect 26099 13413 26108 13447
rect 26056 13404 26108 13413
rect 26700 13404 26752 13456
rect 12532 13268 12584 13320
rect 13176 13200 13228 13252
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 13360 13132 13412 13184
rect 15384 13379 15436 13388
rect 15384 13345 15393 13379
rect 15393 13345 15427 13379
rect 15427 13345 15436 13379
rect 15384 13336 15436 13345
rect 17132 13336 17184 13388
rect 17960 13336 18012 13388
rect 19616 13336 19668 13388
rect 21916 13336 21968 13388
rect 22192 13336 22244 13388
rect 24584 13336 24636 13388
rect 25136 13336 25188 13388
rect 25228 13379 25280 13388
rect 25228 13345 25237 13379
rect 25237 13345 25271 13379
rect 25271 13345 25280 13379
rect 25228 13336 25280 13345
rect 16488 13268 16540 13320
rect 18236 13268 18288 13320
rect 19064 13268 19116 13320
rect 19708 13268 19760 13320
rect 20536 13268 20588 13320
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22560 13268 22612 13320
rect 25504 13379 25556 13388
rect 25504 13345 25513 13379
rect 25513 13345 25547 13379
rect 25547 13345 25556 13379
rect 25504 13336 25556 13345
rect 25596 13379 25648 13388
rect 25596 13345 25605 13379
rect 25605 13345 25639 13379
rect 25639 13345 25648 13379
rect 25596 13336 25648 13345
rect 26424 13336 26476 13388
rect 26608 13379 26660 13388
rect 26608 13345 26617 13379
rect 26617 13345 26651 13379
rect 26651 13345 26660 13379
rect 26608 13336 26660 13345
rect 26976 13404 27028 13456
rect 27988 13404 28040 13456
rect 28172 13404 28224 13456
rect 27620 13379 27672 13388
rect 27620 13345 27654 13379
rect 27654 13345 27672 13379
rect 27620 13336 27672 13345
rect 28632 13336 28684 13388
rect 29092 13379 29144 13388
rect 29092 13345 29101 13379
rect 29101 13345 29135 13379
rect 29135 13345 29144 13379
rect 29092 13336 29144 13345
rect 30748 13268 30800 13320
rect 31024 13311 31076 13320
rect 31024 13277 31033 13311
rect 31033 13277 31067 13311
rect 31067 13277 31076 13311
rect 31024 13268 31076 13277
rect 22376 13200 22428 13252
rect 22652 13200 22704 13252
rect 24216 13200 24268 13252
rect 14372 13132 14424 13184
rect 15568 13132 15620 13184
rect 16580 13175 16632 13184
rect 16580 13141 16589 13175
rect 16589 13141 16623 13175
rect 16623 13141 16632 13175
rect 16580 13132 16632 13141
rect 17132 13175 17184 13184
rect 17132 13141 17141 13175
rect 17141 13141 17175 13175
rect 17175 13141 17184 13175
rect 17132 13132 17184 13141
rect 17592 13132 17644 13184
rect 17776 13132 17828 13184
rect 18420 13175 18472 13184
rect 18420 13141 18429 13175
rect 18429 13141 18463 13175
rect 18463 13141 18472 13175
rect 18420 13132 18472 13141
rect 18604 13132 18656 13184
rect 22836 13132 22888 13184
rect 29552 13175 29604 13184
rect 29552 13141 29561 13175
rect 29561 13141 29595 13175
rect 29595 13141 29604 13175
rect 29552 13132 29604 13141
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 11436 13030 11488 13082
rect 11500 13030 11552 13082
rect 11564 13030 11616 13082
rect 11628 13030 11680 13082
rect 11692 13030 11744 13082
rect 19210 13030 19262 13082
rect 19274 13030 19326 13082
rect 19338 13030 19390 13082
rect 19402 13030 19454 13082
rect 19466 13030 19518 13082
rect 26984 13030 27036 13082
rect 27048 13030 27100 13082
rect 27112 13030 27164 13082
rect 27176 13030 27228 13082
rect 27240 13030 27292 13082
rect 9312 12928 9364 12980
rect 15108 12928 15160 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 16028 12928 16080 12980
rect 18236 12928 18288 12980
rect 18328 12928 18380 12980
rect 19064 12971 19116 12980
rect 19064 12937 19073 12971
rect 19073 12937 19107 12971
rect 19107 12937 19116 12971
rect 19064 12928 19116 12937
rect 29644 12928 29696 12980
rect 31024 12928 31076 12980
rect 2872 12860 2924 12912
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 5448 12724 5500 12776
rect 8208 12792 8260 12844
rect 7104 12767 7156 12776
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 13820 12860 13872 12912
rect 9404 12792 9456 12844
rect 1952 12699 2004 12708
rect 1952 12665 1986 12699
rect 1986 12665 2004 12699
rect 1952 12656 2004 12665
rect 2964 12656 3016 12708
rect 8852 12767 8904 12776
rect 8852 12733 8861 12767
rect 8861 12733 8895 12767
rect 8895 12733 8904 12767
rect 8852 12724 8904 12733
rect 9312 12724 9364 12776
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 11244 12792 11296 12844
rect 9128 12656 9180 12708
rect 11980 12724 12032 12776
rect 12900 12792 12952 12844
rect 12532 12767 12584 12776
rect 11704 12656 11756 12708
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 12624 12767 12676 12776
rect 12624 12733 12633 12767
rect 12633 12733 12667 12767
rect 12667 12733 12676 12767
rect 12624 12724 12676 12733
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 13268 12724 13320 12776
rect 13452 12724 13504 12776
rect 3884 12631 3936 12640
rect 3884 12597 3893 12631
rect 3893 12597 3927 12631
rect 3927 12597 3936 12631
rect 3884 12588 3936 12597
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 8024 12588 8076 12640
rect 8484 12588 8536 12640
rect 11244 12588 11296 12640
rect 13084 12656 13136 12708
rect 13728 12656 13780 12708
rect 14004 12724 14056 12776
rect 14096 12767 14148 12776
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 14372 12767 14424 12776
rect 14372 12733 14406 12767
rect 14406 12733 14424 12767
rect 14372 12724 14424 12733
rect 15476 12724 15528 12776
rect 16028 12792 16080 12844
rect 14004 12588 14056 12640
rect 16488 12860 16540 12912
rect 17500 12860 17552 12912
rect 18144 12860 18196 12912
rect 20352 12860 20404 12912
rect 26700 12860 26752 12912
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 17592 12724 17644 12776
rect 17868 12724 17920 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 15476 12588 15528 12640
rect 16672 12588 16724 12640
rect 18512 12699 18564 12708
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 25964 12767 26016 12776
rect 25964 12733 25973 12767
rect 25973 12733 26007 12767
rect 26007 12733 26016 12767
rect 25964 12724 26016 12733
rect 26148 12767 26200 12776
rect 26148 12733 26157 12767
rect 26157 12733 26191 12767
rect 26191 12733 26200 12767
rect 26148 12724 26200 12733
rect 26332 12724 26384 12776
rect 24860 12656 24912 12708
rect 28080 12724 28132 12776
rect 29552 12767 29604 12776
rect 29552 12733 29586 12767
rect 29586 12733 29604 12767
rect 29552 12724 29604 12733
rect 26332 12631 26384 12640
rect 26332 12597 26341 12631
rect 26341 12597 26375 12631
rect 26375 12597 26384 12631
rect 26332 12588 26384 12597
rect 26424 12588 26476 12640
rect 29092 12631 29144 12640
rect 29092 12597 29101 12631
rect 29101 12597 29135 12631
rect 29135 12597 29144 12631
rect 29092 12588 29144 12597
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 12096 12486 12148 12538
rect 12160 12486 12212 12538
rect 12224 12486 12276 12538
rect 12288 12486 12340 12538
rect 12352 12486 12404 12538
rect 19870 12486 19922 12538
rect 19934 12486 19986 12538
rect 19998 12486 20050 12538
rect 20062 12486 20114 12538
rect 20126 12486 20178 12538
rect 27644 12486 27696 12538
rect 27708 12486 27760 12538
rect 27772 12486 27824 12538
rect 27836 12486 27888 12538
rect 27900 12486 27952 12538
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 3884 12384 3936 12436
rect 2964 12248 3016 12300
rect 3516 12316 3568 12368
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3424 12180 3476 12232
rect 4068 12180 4120 12232
rect 5264 12291 5316 12300
rect 5264 12257 5277 12291
rect 5277 12257 5316 12291
rect 4988 12180 5040 12232
rect 5264 12248 5316 12257
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 6920 12384 6972 12436
rect 8116 12427 8168 12436
rect 8116 12393 8125 12427
rect 8125 12393 8159 12427
rect 8159 12393 8168 12427
rect 8116 12384 8168 12393
rect 9496 12384 9548 12436
rect 11152 12384 11204 12436
rect 8484 12359 8536 12368
rect 8484 12325 8518 12359
rect 8518 12325 8536 12359
rect 8484 12316 8536 12325
rect 7564 12248 7616 12300
rect 8300 12248 8352 12300
rect 5448 12112 5500 12164
rect 2688 12087 2740 12096
rect 2688 12053 2697 12087
rect 2697 12053 2731 12087
rect 2731 12053 2740 12087
rect 2688 12044 2740 12053
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 3424 12044 3476 12096
rect 5540 12044 5592 12096
rect 6184 12044 6236 12096
rect 10048 12316 10100 12368
rect 11060 12316 11112 12368
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 14096 12384 14148 12436
rect 14372 12384 14424 12436
rect 15568 12384 15620 12436
rect 17224 12384 17276 12436
rect 17408 12384 17460 12436
rect 17960 12384 18012 12436
rect 11244 12248 11296 12300
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 11796 12248 11848 12300
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 12164 12248 12216 12300
rect 12900 12291 12952 12300
rect 12900 12257 12909 12291
rect 12909 12257 12943 12291
rect 12943 12257 12952 12291
rect 12900 12248 12952 12257
rect 13268 12248 13320 12300
rect 14556 12248 14608 12300
rect 15752 12316 15804 12368
rect 15292 12248 15344 12300
rect 15660 12248 15712 12300
rect 9864 12044 9916 12096
rect 11244 12044 11296 12096
rect 12532 12112 12584 12164
rect 15384 12112 15436 12164
rect 15752 12155 15804 12164
rect 15752 12121 15761 12155
rect 15761 12121 15795 12155
rect 15795 12121 15804 12155
rect 15752 12112 15804 12121
rect 13820 12044 13872 12096
rect 15844 12044 15896 12096
rect 16580 12316 16632 12368
rect 18420 12316 18472 12368
rect 19616 12384 19668 12436
rect 16212 12248 16264 12300
rect 17132 12248 17184 12300
rect 19064 12248 19116 12300
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 20536 12316 20588 12368
rect 22192 12359 22244 12368
rect 22192 12325 22201 12359
rect 22201 12325 22235 12359
rect 22235 12325 22244 12359
rect 22192 12316 22244 12325
rect 22468 12316 22520 12368
rect 22560 12316 22612 12368
rect 25964 12384 26016 12436
rect 25688 12316 25740 12368
rect 18880 12180 18932 12232
rect 19892 12180 19944 12232
rect 20536 12180 20588 12232
rect 18972 12112 19024 12164
rect 20260 12112 20312 12164
rect 20444 12112 20496 12164
rect 22192 12180 22244 12232
rect 22744 12180 22796 12232
rect 22836 12180 22888 12232
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 24032 12248 24084 12300
rect 25320 12248 25372 12300
rect 25504 12248 25556 12300
rect 25872 12291 25924 12300
rect 25872 12257 25881 12291
rect 25881 12257 25915 12291
rect 25915 12257 25924 12291
rect 25872 12248 25924 12257
rect 25964 12291 26016 12300
rect 25964 12257 25973 12291
rect 25973 12257 26007 12291
rect 26007 12257 26016 12291
rect 25964 12248 26016 12257
rect 26332 12248 26384 12300
rect 28632 12384 28684 12436
rect 30748 12427 30800 12436
rect 30748 12393 30757 12427
rect 30757 12393 30791 12427
rect 30791 12393 30800 12427
rect 30748 12384 30800 12393
rect 26516 12316 26568 12368
rect 26148 12180 26200 12232
rect 26608 12291 26660 12300
rect 26608 12257 26617 12291
rect 26617 12257 26651 12291
rect 26651 12257 26660 12291
rect 26608 12248 26660 12257
rect 29000 12316 29052 12368
rect 26884 12248 26936 12300
rect 27436 12248 27488 12300
rect 29092 12248 29144 12300
rect 16120 12044 16172 12096
rect 25872 12112 25924 12164
rect 26792 12112 26844 12164
rect 21456 12044 21508 12096
rect 23388 12044 23440 12096
rect 25044 12087 25096 12096
rect 25044 12053 25053 12087
rect 25053 12053 25087 12087
rect 25087 12053 25096 12087
rect 25044 12044 25096 12053
rect 25780 12044 25832 12096
rect 25964 12044 26016 12096
rect 27712 12112 27764 12164
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 11436 11942 11488 11994
rect 11500 11942 11552 11994
rect 11564 11942 11616 11994
rect 11628 11942 11680 11994
rect 11692 11942 11744 11994
rect 19210 11942 19262 11994
rect 19274 11942 19326 11994
rect 19338 11942 19390 11994
rect 19402 11942 19454 11994
rect 19466 11942 19518 11994
rect 26984 11942 27036 11994
rect 27048 11942 27100 11994
rect 27112 11942 27164 11994
rect 27176 11942 27228 11994
rect 27240 11942 27292 11994
rect 3240 11840 3292 11892
rect 4252 11840 4304 11892
rect 5356 11840 5408 11892
rect 7564 11883 7616 11892
rect 7564 11849 7573 11883
rect 7573 11849 7607 11883
rect 7607 11849 7616 11883
rect 7564 11840 7616 11849
rect 12440 11840 12492 11892
rect 19800 11840 19852 11892
rect 21272 11840 21324 11892
rect 22652 11840 22704 11892
rect 26884 11840 26936 11892
rect 4988 11815 5040 11824
rect 4988 11781 4997 11815
rect 4997 11781 5031 11815
rect 5031 11781 5040 11815
rect 4988 11772 5040 11781
rect 2872 11704 2924 11756
rect 5264 11772 5316 11824
rect 16212 11772 16264 11824
rect 17132 11772 17184 11824
rect 18144 11772 18196 11824
rect 20536 11815 20588 11824
rect 20536 11781 20545 11815
rect 20545 11781 20579 11815
rect 20579 11781 20588 11815
rect 20536 11772 20588 11781
rect 26056 11772 26108 11824
rect 27988 11840 28040 11892
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 2688 11636 2740 11688
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 4068 11636 4120 11688
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 1216 11543 1268 11552
rect 1216 11509 1225 11543
rect 1225 11509 1259 11543
rect 1259 11509 1268 11543
rect 1216 11500 1268 11509
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 5448 11679 5500 11688
rect 5448 11645 5455 11679
rect 5455 11645 5500 11679
rect 5448 11636 5500 11645
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 5724 11679 5776 11688
rect 8852 11704 8904 11756
rect 5724 11645 5738 11679
rect 5738 11645 5772 11679
rect 5772 11645 5776 11679
rect 5724 11636 5776 11645
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 9128 11636 9180 11688
rect 11152 11636 11204 11688
rect 12072 11704 12124 11756
rect 11336 11636 11388 11688
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 16672 11704 16724 11756
rect 17684 11704 17736 11756
rect 17868 11704 17920 11756
rect 19892 11704 19944 11756
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 8760 11568 8812 11620
rect 13084 11679 13136 11688
rect 13084 11645 13093 11679
rect 13093 11645 13127 11679
rect 13127 11645 13136 11679
rect 13084 11636 13136 11645
rect 18144 11636 18196 11688
rect 6092 11500 6144 11552
rect 9312 11500 9364 11552
rect 11796 11500 11848 11552
rect 17868 11611 17920 11620
rect 17868 11577 17877 11611
rect 17877 11577 17911 11611
rect 17911 11577 17920 11611
rect 17868 11568 17920 11577
rect 18972 11636 19024 11688
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 21456 11679 21508 11688
rect 21456 11645 21465 11679
rect 21465 11645 21499 11679
rect 21499 11645 21508 11679
rect 21456 11636 21508 11645
rect 21732 11679 21784 11688
rect 21732 11645 21741 11679
rect 21741 11645 21775 11679
rect 21775 11645 21784 11679
rect 21732 11636 21784 11645
rect 23296 11704 23348 11756
rect 18788 11568 18840 11620
rect 20168 11568 20220 11620
rect 20996 11568 21048 11620
rect 12624 11500 12676 11552
rect 15200 11500 15252 11552
rect 15844 11500 15896 11552
rect 16028 11500 16080 11552
rect 19708 11500 19760 11552
rect 22468 11636 22520 11688
rect 23020 11636 23072 11688
rect 23388 11679 23440 11688
rect 23388 11645 23397 11679
rect 23397 11645 23431 11679
rect 23431 11645 23440 11679
rect 23388 11636 23440 11645
rect 23664 11636 23716 11688
rect 24860 11704 24912 11756
rect 25044 11636 25096 11688
rect 27712 11679 27764 11688
rect 27712 11645 27730 11679
rect 27730 11645 27764 11679
rect 27712 11636 27764 11645
rect 29000 11636 29052 11688
rect 30288 11636 30340 11688
rect 30840 11636 30892 11688
rect 22192 11568 22244 11620
rect 23112 11500 23164 11552
rect 23204 11543 23256 11552
rect 23204 11509 23213 11543
rect 23213 11509 23247 11543
rect 23247 11509 23256 11543
rect 23204 11500 23256 11509
rect 23480 11500 23532 11552
rect 25596 11500 25648 11552
rect 29368 11500 29420 11552
rect 29920 11543 29972 11552
rect 29920 11509 29929 11543
rect 29929 11509 29963 11543
rect 29963 11509 29972 11543
rect 29920 11500 29972 11509
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 12096 11398 12148 11450
rect 12160 11398 12212 11450
rect 12224 11398 12276 11450
rect 12288 11398 12340 11450
rect 12352 11398 12404 11450
rect 19870 11398 19922 11450
rect 19934 11398 19986 11450
rect 19998 11398 20050 11450
rect 20062 11398 20114 11450
rect 20126 11398 20178 11450
rect 27644 11398 27696 11450
rect 27708 11398 27760 11450
rect 27772 11398 27824 11450
rect 27836 11398 27888 11450
rect 27900 11398 27952 11450
rect 4252 11296 4304 11348
rect 2688 11228 2740 11280
rect 1216 11160 1268 11212
rect 2412 11160 2464 11212
rect 5908 11296 5960 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 5540 11160 5592 11212
rect 2872 11024 2924 11076
rect 4160 11092 4212 11144
rect 5724 11092 5776 11144
rect 6092 11203 6144 11212
rect 6092 11169 6101 11203
rect 6101 11169 6135 11203
rect 6135 11169 6144 11203
rect 6092 11160 6144 11169
rect 6368 11203 6420 11212
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 10048 11296 10100 11348
rect 14924 11296 14976 11348
rect 15568 11339 15620 11348
rect 15568 11305 15577 11339
rect 15577 11305 15611 11339
rect 15611 11305 15620 11339
rect 15568 11296 15620 11305
rect 19064 11296 19116 11348
rect 9312 11228 9364 11280
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 9128 11160 9180 11169
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 9404 11203 9456 11212
rect 9404 11169 9413 11203
rect 9413 11169 9447 11203
rect 9447 11169 9456 11203
rect 9404 11160 9456 11169
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 4896 11024 4948 11076
rect 5264 11024 5316 11076
rect 15844 11203 15896 11212
rect 15844 11169 15853 11203
rect 15853 11169 15887 11203
rect 15887 11169 15896 11203
rect 15844 11160 15896 11169
rect 16396 11203 16448 11212
rect 16396 11169 16405 11203
rect 16405 11169 16439 11203
rect 16439 11169 16448 11203
rect 16396 11160 16448 11169
rect 4068 10999 4120 11008
rect 4068 10965 4077 10999
rect 4077 10965 4111 10999
rect 4111 10965 4120 10999
rect 4068 10956 4120 10965
rect 4804 10956 4856 11008
rect 9956 10956 10008 11008
rect 14280 10956 14332 11008
rect 15752 11092 15804 11144
rect 19524 11296 19576 11348
rect 20536 11296 20588 11348
rect 21732 11296 21784 11348
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 25872 11296 25924 11348
rect 26608 11296 26660 11348
rect 27344 11296 27396 11348
rect 23204 11271 23256 11280
rect 23204 11237 23222 11271
rect 23222 11237 23256 11271
rect 23204 11228 23256 11237
rect 26700 11271 26752 11280
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 19984 11160 20036 11212
rect 20076 11203 20128 11212
rect 20076 11169 20085 11203
rect 20085 11169 20119 11203
rect 20119 11169 20128 11203
rect 20076 11160 20128 11169
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 20260 11203 20312 11212
rect 20260 11169 20269 11203
rect 20269 11169 20303 11203
rect 20303 11169 20312 11203
rect 20260 11160 20312 11169
rect 20352 11203 20404 11212
rect 20352 11169 20387 11203
rect 20387 11169 20404 11203
rect 20352 11160 20404 11169
rect 21180 11160 21232 11212
rect 23480 11203 23532 11212
rect 23480 11169 23489 11203
rect 23489 11169 23523 11203
rect 23523 11169 23532 11203
rect 23480 11160 23532 11169
rect 24032 11160 24084 11212
rect 25504 11203 25556 11212
rect 25504 11169 25513 11203
rect 25513 11169 25547 11203
rect 25547 11169 25556 11203
rect 25504 11160 25556 11169
rect 25596 11203 25648 11212
rect 25596 11169 25605 11203
rect 25605 11169 25639 11203
rect 25639 11169 25648 11203
rect 25596 11160 25648 11169
rect 25780 11203 25832 11212
rect 25780 11169 25815 11203
rect 25815 11169 25832 11203
rect 25780 11160 25832 11169
rect 25964 11203 26016 11212
rect 25964 11169 25973 11203
rect 25973 11169 26007 11203
rect 26007 11169 26016 11203
rect 25964 11160 26016 11169
rect 26056 11203 26108 11212
rect 26056 11169 26065 11203
rect 26065 11169 26099 11203
rect 26099 11169 26108 11203
rect 26056 11160 26108 11169
rect 26240 11203 26292 11212
rect 26240 11169 26249 11203
rect 26249 11169 26283 11203
rect 26283 11169 26292 11203
rect 26240 11160 26292 11169
rect 26424 11203 26476 11212
rect 26424 11169 26433 11203
rect 26433 11169 26467 11203
rect 26467 11169 26476 11203
rect 26424 11160 26476 11169
rect 26700 11237 26734 11271
rect 26734 11237 26752 11271
rect 26700 11228 26752 11237
rect 20536 11135 20588 11144
rect 20536 11101 20545 11135
rect 20545 11101 20579 11135
rect 20579 11101 20588 11135
rect 20536 11092 20588 11101
rect 28632 11203 28684 11212
rect 28632 11169 28641 11203
rect 28641 11169 28675 11203
rect 28675 11169 28684 11203
rect 28632 11160 28684 11169
rect 28816 11203 28868 11212
rect 28816 11169 28825 11203
rect 28825 11169 28859 11203
rect 28859 11169 28868 11203
rect 28816 11160 28868 11169
rect 29920 11296 29972 11348
rect 29368 11203 29420 11212
rect 29368 11169 29377 11203
rect 29377 11169 29411 11203
rect 29411 11169 29420 11203
rect 29368 11160 29420 11169
rect 29092 11092 29144 11144
rect 19340 11024 19392 11076
rect 20168 11024 20220 11076
rect 20904 11024 20956 11076
rect 22468 11024 22520 11076
rect 16580 10999 16632 11008
rect 16580 10965 16589 10999
rect 16589 10965 16623 10999
rect 16623 10965 16632 10999
rect 16580 10956 16632 10965
rect 16856 10956 16908 11008
rect 17592 10956 17644 11008
rect 19616 10956 19668 11008
rect 19984 10956 20036 11008
rect 29184 11024 29236 11076
rect 30840 11024 30892 11076
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 11436 10854 11488 10906
rect 11500 10854 11552 10906
rect 11564 10854 11616 10906
rect 11628 10854 11680 10906
rect 11692 10854 11744 10906
rect 19210 10854 19262 10906
rect 19274 10854 19326 10906
rect 19338 10854 19390 10906
rect 19402 10854 19454 10906
rect 19466 10854 19518 10906
rect 26984 10854 27036 10906
rect 27048 10854 27100 10906
rect 27112 10854 27164 10906
rect 27176 10854 27228 10906
rect 27240 10854 27292 10906
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 5540 10752 5592 10804
rect 2780 10684 2832 10736
rect 3332 10684 3384 10736
rect 4068 10684 4120 10736
rect 9864 10752 9916 10804
rect 9956 10752 10008 10804
rect 8760 10684 8812 10736
rect 9128 10684 9180 10736
rect 15844 10752 15896 10804
rect 16488 10752 16540 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 22376 10752 22428 10804
rect 26516 10684 26568 10736
rect 26792 10752 26844 10804
rect 28816 10752 28868 10804
rect 27160 10684 27212 10736
rect 28080 10684 28132 10736
rect 2596 10591 2648 10600
rect 2596 10557 2605 10591
rect 2605 10557 2639 10591
rect 2639 10557 2648 10591
rect 2596 10548 2648 10557
rect 2872 10548 2924 10600
rect 3148 10548 3200 10600
rect 4160 10548 4212 10600
rect 6276 10616 6328 10668
rect 7104 10616 7156 10668
rect 7840 10616 7892 10668
rect 6368 10548 6420 10600
rect 2136 10412 2188 10464
rect 6092 10480 6144 10532
rect 6000 10412 6052 10464
rect 7840 10523 7892 10532
rect 7840 10489 7849 10523
rect 7849 10489 7883 10523
rect 7883 10489 7892 10523
rect 7840 10480 7892 10489
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8760 10548 8812 10557
rect 9036 10591 9088 10600
rect 9036 10557 9045 10591
rect 9045 10557 9079 10591
rect 9079 10557 9088 10591
rect 9036 10548 9088 10557
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 9864 10548 9916 10600
rect 9496 10480 9548 10532
rect 10416 10523 10468 10532
rect 10416 10489 10425 10523
rect 10425 10489 10459 10523
rect 10459 10489 10468 10523
rect 10416 10480 10468 10489
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 8760 10412 8812 10464
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 11980 10480 12032 10532
rect 13084 10480 13136 10532
rect 13452 10480 13504 10532
rect 14648 10591 14700 10600
rect 14648 10557 14657 10591
rect 14657 10557 14691 10591
rect 14691 10557 14700 10591
rect 14648 10548 14700 10557
rect 15200 10548 15252 10600
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 24216 10616 24268 10668
rect 24860 10616 24912 10668
rect 17684 10548 17736 10600
rect 13176 10412 13228 10464
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 16580 10480 16632 10532
rect 16764 10480 16816 10532
rect 18788 10591 18840 10600
rect 18788 10557 18797 10591
rect 18797 10557 18831 10591
rect 18831 10557 18840 10591
rect 18788 10548 18840 10557
rect 18972 10548 19024 10600
rect 19616 10548 19668 10600
rect 21180 10591 21232 10600
rect 21180 10557 21189 10591
rect 21189 10557 21223 10591
rect 21223 10557 21232 10591
rect 21180 10548 21232 10557
rect 24032 10591 24084 10600
rect 24032 10557 24041 10591
rect 24041 10557 24075 10591
rect 24075 10557 24084 10591
rect 24032 10548 24084 10557
rect 25136 10548 25188 10600
rect 26332 10548 26384 10600
rect 27344 10548 27396 10600
rect 30840 10684 30892 10736
rect 29184 10616 29236 10668
rect 18328 10480 18380 10532
rect 17224 10412 17276 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 19892 10412 19944 10464
rect 21088 10455 21140 10464
rect 21088 10421 21097 10455
rect 21097 10421 21131 10455
rect 21131 10421 21140 10455
rect 21088 10412 21140 10421
rect 23940 10412 23992 10464
rect 24032 10412 24084 10464
rect 25780 10480 25832 10532
rect 26240 10480 26292 10532
rect 29092 10591 29144 10600
rect 29092 10557 29101 10591
rect 29101 10557 29135 10591
rect 29135 10557 29144 10591
rect 29092 10548 29144 10557
rect 29276 10591 29328 10600
rect 29276 10557 29285 10591
rect 29285 10557 29319 10591
rect 29319 10557 29328 10591
rect 29276 10548 29328 10557
rect 30104 10591 30156 10600
rect 30104 10557 30113 10591
rect 30113 10557 30147 10591
rect 30147 10557 30156 10591
rect 30104 10548 30156 10557
rect 30288 10548 30340 10600
rect 25504 10455 25556 10464
rect 25504 10421 25513 10455
rect 25513 10421 25547 10455
rect 25547 10421 25556 10455
rect 25504 10412 25556 10421
rect 26700 10412 26752 10464
rect 27988 10412 28040 10464
rect 28632 10412 28684 10464
rect 30012 10455 30064 10464
rect 30012 10421 30021 10455
rect 30021 10421 30055 10455
rect 30055 10421 30064 10455
rect 30012 10412 30064 10421
rect 30748 10412 30800 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 12096 10310 12148 10362
rect 12160 10310 12212 10362
rect 12224 10310 12276 10362
rect 12288 10310 12340 10362
rect 12352 10310 12404 10362
rect 19870 10310 19922 10362
rect 19934 10310 19986 10362
rect 19998 10310 20050 10362
rect 20062 10310 20114 10362
rect 20126 10310 20178 10362
rect 27644 10310 27696 10362
rect 27708 10310 27760 10362
rect 27772 10310 27824 10362
rect 27836 10310 27888 10362
rect 27900 10310 27952 10362
rect 2780 10208 2832 10260
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 5080 10251 5132 10260
rect 5080 10217 5089 10251
rect 5089 10217 5123 10251
rect 5123 10217 5132 10251
rect 5080 10208 5132 10217
rect 6368 10208 6420 10260
rect 7932 10208 7984 10260
rect 8208 10208 8260 10260
rect 9036 10208 9088 10260
rect 9128 10208 9180 10260
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 3516 10140 3568 10192
rect 2780 10072 2832 10124
rect 6828 10140 6880 10192
rect 8392 10140 8444 10192
rect 4988 10072 5040 10124
rect 4252 10004 4304 10056
rect 5080 10004 5132 10056
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 5908 10072 5960 10124
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 8760 10115 8812 10124
rect 8760 10081 8769 10115
rect 8769 10081 8803 10115
rect 8803 10081 8812 10115
rect 8760 10072 8812 10081
rect 8944 10072 8996 10124
rect 5724 10004 5776 10056
rect 9404 10072 9456 10124
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9680 10004 9732 10056
rect 11888 10208 11940 10260
rect 11980 10251 12032 10260
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 14648 10208 14700 10260
rect 15936 10208 15988 10260
rect 16120 10208 16172 10260
rect 16396 10208 16448 10260
rect 17224 10251 17276 10260
rect 17224 10217 17233 10251
rect 17233 10217 17267 10251
rect 17267 10217 17276 10251
rect 17224 10208 17276 10217
rect 11152 10140 11204 10192
rect 11244 10140 11296 10192
rect 10600 10115 10652 10124
rect 10600 10081 10609 10115
rect 10609 10081 10643 10115
rect 10643 10081 10652 10115
rect 10600 10072 10652 10081
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 13636 10140 13688 10192
rect 11428 10004 11480 10056
rect 13084 10072 13136 10124
rect 13176 10115 13228 10124
rect 13176 10081 13185 10115
rect 13185 10081 13219 10115
rect 13219 10081 13228 10115
rect 13176 10072 13228 10081
rect 13452 10115 13504 10124
rect 13452 10081 13486 10115
rect 13486 10081 13504 10115
rect 13452 10072 13504 10081
rect 13728 10072 13780 10124
rect 15016 10115 15068 10124
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15016 10072 15068 10081
rect 15200 10115 15252 10124
rect 15200 10081 15209 10115
rect 15209 10081 15243 10115
rect 15243 10081 15252 10115
rect 15200 10072 15252 10081
rect 15752 10072 15804 10124
rect 16764 10183 16816 10192
rect 16764 10149 16773 10183
rect 16773 10149 16807 10183
rect 16807 10149 16816 10183
rect 16764 10140 16816 10149
rect 16856 10183 16908 10192
rect 16856 10149 16865 10183
rect 16865 10149 16899 10183
rect 16899 10149 16908 10183
rect 16856 10140 16908 10149
rect 16948 10183 17000 10192
rect 16948 10149 16983 10183
rect 16983 10149 17000 10183
rect 16948 10140 17000 10149
rect 16396 10072 16448 10124
rect 16672 10115 16724 10124
rect 16672 10081 16681 10115
rect 16681 10081 16715 10115
rect 16715 10081 16724 10115
rect 16672 10072 16724 10081
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 17316 10140 17368 10192
rect 17592 10183 17644 10192
rect 17592 10149 17601 10183
rect 17601 10149 17635 10183
rect 17635 10149 17644 10183
rect 17592 10140 17644 10149
rect 20352 10208 20404 10260
rect 20720 10208 20772 10260
rect 21088 10140 21140 10192
rect 19984 10115 20036 10124
rect 19984 10081 20018 10115
rect 20018 10081 20036 10115
rect 19984 10072 20036 10081
rect 22376 10115 22428 10124
rect 22376 10081 22385 10115
rect 22385 10081 22419 10115
rect 22419 10081 22428 10115
rect 22376 10072 22428 10081
rect 25504 10140 25556 10192
rect 27436 10208 27488 10260
rect 27988 10208 28040 10260
rect 30104 10208 30156 10260
rect 26240 10140 26292 10192
rect 23940 10115 23992 10124
rect 23940 10081 23974 10115
rect 23974 10081 23992 10115
rect 23940 10072 23992 10081
rect 25412 10072 25464 10124
rect 18052 10004 18104 10056
rect 8760 9936 8812 9988
rect 9036 9936 9088 9988
rect 12808 9936 12860 9988
rect 1952 9868 2004 9920
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 4068 9868 4120 9920
rect 5632 9868 5684 9920
rect 6000 9868 6052 9920
rect 8852 9911 8904 9920
rect 8852 9877 8861 9911
rect 8861 9877 8895 9911
rect 8895 9877 8904 9911
rect 8852 9868 8904 9877
rect 10140 9911 10192 9920
rect 10140 9877 10149 9911
rect 10149 9877 10183 9911
rect 10183 9877 10192 9911
rect 10140 9868 10192 9877
rect 11336 9868 11388 9920
rect 12072 9868 12124 9920
rect 14280 9868 14332 9920
rect 15108 9868 15160 9920
rect 16672 9868 16724 9920
rect 20812 9936 20864 9988
rect 23296 10004 23348 10056
rect 26700 10115 26752 10124
rect 26700 10081 26709 10115
rect 26709 10081 26743 10115
rect 26743 10081 26752 10115
rect 26700 10072 26752 10081
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 27436 10115 27488 10124
rect 27436 10081 27445 10115
rect 27445 10081 27479 10115
rect 27479 10081 27488 10115
rect 27436 10072 27488 10081
rect 27528 10115 27580 10124
rect 27528 10081 27537 10115
rect 27537 10081 27571 10115
rect 27571 10081 27580 10115
rect 27528 10072 27580 10081
rect 28632 10140 28684 10192
rect 28908 10183 28960 10192
rect 28908 10149 28917 10183
rect 28917 10149 28951 10183
rect 28951 10149 28960 10183
rect 28908 10140 28960 10149
rect 29920 10140 29972 10192
rect 30012 10140 30064 10192
rect 21456 9868 21508 9920
rect 22560 9911 22612 9920
rect 22560 9877 22569 9911
rect 22569 9877 22603 9911
rect 22603 9877 22612 9911
rect 22560 9868 22612 9877
rect 23388 9868 23440 9920
rect 25136 9868 25188 9920
rect 25780 9936 25832 9988
rect 26884 9936 26936 9988
rect 27160 10047 27212 10056
rect 27160 10013 27169 10047
rect 27169 10013 27203 10047
rect 27203 10013 27212 10047
rect 27160 10004 27212 10013
rect 28448 10072 28500 10124
rect 29460 10072 29512 10124
rect 30748 10115 30800 10124
rect 30748 10081 30757 10115
rect 30757 10081 30791 10115
rect 30791 10081 30800 10115
rect 30748 10072 30800 10081
rect 29276 10004 29328 10056
rect 28080 9936 28132 9988
rect 26056 9911 26108 9920
rect 26056 9877 26065 9911
rect 26065 9877 26099 9911
rect 26099 9877 26108 9911
rect 26056 9868 26108 9877
rect 27896 9911 27948 9920
rect 27896 9877 27905 9911
rect 27905 9877 27939 9911
rect 27939 9877 27948 9911
rect 27896 9868 27948 9877
rect 29184 9868 29236 9920
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 11436 9766 11488 9818
rect 11500 9766 11552 9818
rect 11564 9766 11616 9818
rect 11628 9766 11680 9818
rect 11692 9766 11744 9818
rect 19210 9766 19262 9818
rect 19274 9766 19326 9818
rect 19338 9766 19390 9818
rect 19402 9766 19454 9818
rect 19466 9766 19518 9818
rect 26984 9766 27036 9818
rect 27048 9766 27100 9818
rect 27112 9766 27164 9818
rect 27176 9766 27228 9818
rect 27240 9766 27292 9818
rect 2780 9664 2832 9716
rect 3424 9596 3476 9648
rect 2872 9528 2924 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 1952 9503 2004 9512
rect 1952 9469 1986 9503
rect 1986 9469 2004 9503
rect 1952 9460 2004 9469
rect 5356 9664 5408 9716
rect 5724 9664 5776 9716
rect 5908 9664 5960 9716
rect 7104 9664 7156 9716
rect 8760 9664 8812 9716
rect 4712 9596 4764 9648
rect 4988 9596 5040 9648
rect 6000 9596 6052 9648
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 4620 9460 4672 9512
rect 2596 9392 2648 9444
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 5632 9528 5684 9580
rect 5724 9528 5776 9580
rect 6828 9596 6880 9648
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 6368 9460 6420 9512
rect 6460 9503 6512 9512
rect 6460 9469 6469 9503
rect 6469 9469 6503 9503
rect 6503 9469 6512 9503
rect 6460 9460 6512 9469
rect 1216 9367 1268 9376
rect 1216 9333 1225 9367
rect 1225 9333 1259 9367
rect 1259 9333 1268 9367
rect 1216 9324 1268 9333
rect 5724 9392 5776 9444
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7656 9460 7708 9512
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 8300 9460 8352 9512
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 10416 9664 10468 9716
rect 13452 9664 13504 9716
rect 19984 9664 20036 9716
rect 20536 9664 20588 9716
rect 25780 9664 25832 9716
rect 26240 9664 26292 9716
rect 26792 9664 26844 9716
rect 26884 9664 26936 9716
rect 28816 9664 28868 9716
rect 29000 9664 29052 9716
rect 29920 9664 29972 9716
rect 10692 9460 10744 9512
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 12532 9460 12584 9512
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 8852 9392 8904 9444
rect 10140 9392 10192 9444
rect 11060 9392 11112 9444
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 17316 9596 17368 9648
rect 17592 9596 17644 9648
rect 14556 9528 14608 9580
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 14556 9392 14608 9444
rect 15200 9392 15252 9444
rect 15936 9528 15988 9580
rect 18144 9528 18196 9580
rect 19064 9528 19116 9580
rect 15844 9460 15896 9512
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 16396 9503 16448 9512
rect 16396 9469 16405 9503
rect 16405 9469 16439 9503
rect 16439 9469 16448 9503
rect 16396 9460 16448 9469
rect 18328 9460 18380 9512
rect 20352 9503 20404 9512
rect 20352 9469 20361 9503
rect 20361 9469 20395 9503
rect 20395 9469 20404 9503
rect 20352 9460 20404 9469
rect 20812 9528 20864 9580
rect 20720 9503 20772 9512
rect 20720 9469 20729 9503
rect 20729 9469 20763 9503
rect 20763 9469 20772 9503
rect 20720 9460 20772 9469
rect 19340 9392 19392 9444
rect 20536 9435 20588 9444
rect 20536 9401 20571 9435
rect 20571 9401 20588 9435
rect 21180 9528 21232 9580
rect 22192 9528 22244 9580
rect 22560 9503 22612 9512
rect 22560 9469 22594 9503
rect 22594 9469 22612 9503
rect 22560 9460 22612 9469
rect 24492 9460 24544 9512
rect 20536 9392 20588 9401
rect 23572 9392 23624 9444
rect 24308 9392 24360 9444
rect 27896 9460 27948 9512
rect 28172 9460 28224 9512
rect 26056 9392 26108 9444
rect 9128 9324 9180 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 11612 9324 11664 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 14740 9324 14792 9376
rect 19616 9324 19668 9376
rect 21640 9324 21692 9376
rect 23756 9324 23808 9376
rect 25228 9367 25280 9376
rect 25228 9333 25237 9367
rect 25237 9333 25271 9367
rect 25271 9333 25280 9367
rect 25228 9324 25280 9333
rect 25320 9367 25372 9376
rect 25320 9333 25329 9367
rect 25329 9333 25363 9367
rect 25363 9333 25372 9367
rect 25320 9324 25372 9333
rect 27988 9324 28040 9376
rect 28540 9503 28592 9512
rect 28540 9469 28549 9503
rect 28549 9469 28583 9503
rect 28583 9469 28592 9503
rect 28540 9460 28592 9469
rect 29184 9528 29236 9580
rect 28724 9367 28776 9376
rect 28724 9333 28733 9367
rect 28733 9333 28767 9367
rect 28767 9333 28776 9367
rect 28724 9324 28776 9333
rect 29276 9324 29328 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 12096 9222 12148 9274
rect 12160 9222 12212 9274
rect 12224 9222 12276 9274
rect 12288 9222 12340 9274
rect 12352 9222 12404 9274
rect 19870 9222 19922 9274
rect 19934 9222 19986 9274
rect 19998 9222 20050 9274
rect 20062 9222 20114 9274
rect 20126 9222 20178 9274
rect 27644 9222 27696 9274
rect 27708 9222 27760 9274
rect 27772 9222 27824 9274
rect 27836 9222 27888 9274
rect 27900 9222 27952 9274
rect 1216 8984 1268 9036
rect 2504 8984 2556 9036
rect 5816 9120 5868 9172
rect 6460 9120 6512 9172
rect 7288 9120 7340 9172
rect 9404 9120 9456 9172
rect 11704 9120 11756 9172
rect 6000 9027 6052 9036
rect 6000 8993 6009 9027
rect 6009 8993 6043 9027
rect 6043 8993 6052 9027
rect 6000 8984 6052 8993
rect 8300 9052 8352 9104
rect 8760 9052 8812 9104
rect 3240 8916 3292 8968
rect 3516 8959 3568 8968
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 4344 8916 4396 8968
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 8208 8984 8260 9036
rect 8484 8984 8536 9036
rect 10324 9052 10376 9104
rect 9772 8984 9824 9036
rect 11612 8984 11664 9036
rect 11888 9052 11940 9104
rect 12532 9120 12584 9172
rect 14740 9120 14792 9172
rect 16120 9120 16172 9172
rect 22376 9120 22428 9172
rect 22560 9120 22612 9172
rect 22744 9120 22796 9172
rect 22836 9120 22888 9172
rect 14556 9052 14608 9104
rect 18788 9052 18840 9104
rect 12716 8984 12768 9036
rect 14464 8984 14516 9036
rect 15292 8984 15344 9036
rect 15660 8984 15712 9036
rect 4068 8848 4120 8900
rect 3516 8780 3568 8832
rect 4252 8780 4304 8832
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 5816 8780 5868 8832
rect 6368 8780 6420 8832
rect 17408 8984 17460 9036
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 14280 8848 14332 8900
rect 18144 8916 18196 8968
rect 17960 8848 18012 8900
rect 18420 8916 18472 8968
rect 18972 8848 19024 8900
rect 20352 8984 20404 9036
rect 22192 9052 22244 9104
rect 27436 9120 27488 9172
rect 21180 8984 21232 9036
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 22376 8984 22428 9036
rect 25320 9052 25372 9104
rect 26516 9052 26568 9104
rect 27528 9052 27580 9104
rect 27988 9052 28040 9104
rect 22284 8916 22336 8968
rect 22836 8984 22888 9036
rect 23572 8984 23624 9036
rect 24032 9027 24084 9036
rect 24032 8993 24041 9027
rect 24041 8993 24075 9027
rect 24075 8993 24084 9027
rect 24032 8984 24084 8993
rect 24124 9027 24176 9036
rect 24124 8993 24133 9027
rect 24133 8993 24167 9027
rect 24167 8993 24176 9027
rect 24124 8984 24176 8993
rect 13544 8780 13596 8832
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 18880 8780 18932 8832
rect 19708 8848 19760 8900
rect 21824 8848 21876 8900
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 24216 8916 24268 8968
rect 24308 8959 24360 8968
rect 24308 8925 24317 8959
rect 24317 8925 24351 8959
rect 24351 8925 24360 8959
rect 24308 8916 24360 8925
rect 24860 8984 24912 9036
rect 28724 8984 28776 9036
rect 29000 9027 29052 9036
rect 29000 8993 29009 9027
rect 29009 8993 29043 9027
rect 29043 8993 29052 9027
rect 29000 8984 29052 8993
rect 29276 9027 29328 9036
rect 29276 8993 29285 9027
rect 29285 8993 29319 9027
rect 29319 8993 29328 9027
rect 29276 8984 29328 8993
rect 23756 8848 23808 8900
rect 24584 8848 24636 8900
rect 26516 8891 26568 8900
rect 26516 8857 26525 8891
rect 26525 8857 26559 8891
rect 26559 8857 26568 8891
rect 26516 8848 26568 8857
rect 20904 8780 20956 8832
rect 24492 8823 24544 8832
rect 24492 8789 24501 8823
rect 24501 8789 24535 8823
rect 24535 8789 24544 8823
rect 24492 8780 24544 8789
rect 25780 8780 25832 8832
rect 26332 8780 26384 8832
rect 28632 8916 28684 8968
rect 29460 8780 29512 8832
rect 30656 8823 30708 8832
rect 30656 8789 30665 8823
rect 30665 8789 30699 8823
rect 30699 8789 30708 8823
rect 30656 8780 30708 8789
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 11436 8678 11488 8730
rect 11500 8678 11552 8730
rect 11564 8678 11616 8730
rect 11628 8678 11680 8730
rect 11692 8678 11744 8730
rect 19210 8678 19262 8730
rect 19274 8678 19326 8730
rect 19338 8678 19390 8730
rect 19402 8678 19454 8730
rect 19466 8678 19518 8730
rect 26984 8678 27036 8730
rect 27048 8678 27100 8730
rect 27112 8678 27164 8730
rect 27176 8678 27228 8730
rect 27240 8678 27292 8730
rect 2504 8576 2556 8628
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 1400 8440 1452 8492
rect 2596 8415 2648 8424
rect 2596 8381 2605 8415
rect 2605 8381 2639 8415
rect 2639 8381 2648 8415
rect 2596 8372 2648 8381
rect 6000 8576 6052 8628
rect 8392 8576 8444 8628
rect 17408 8576 17460 8628
rect 18972 8576 19024 8628
rect 21272 8576 21324 8628
rect 4344 8551 4396 8560
rect 4344 8517 4353 8551
rect 4353 8517 4387 8551
rect 4387 8517 4396 8551
rect 4344 8508 4396 8517
rect 18696 8508 18748 8560
rect 21640 8576 21692 8628
rect 22376 8576 22428 8628
rect 22744 8576 22796 8628
rect 22928 8576 22980 8628
rect 25688 8576 25740 8628
rect 25964 8619 26016 8628
rect 25964 8585 25973 8619
rect 25973 8585 26007 8619
rect 26007 8585 26016 8619
rect 25964 8576 26016 8585
rect 4160 8440 4212 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 3240 8304 3292 8356
rect 3424 8347 3476 8356
rect 3424 8313 3451 8347
rect 3451 8313 3476 8347
rect 3424 8304 3476 8313
rect 3516 8304 3568 8356
rect 4804 8372 4856 8424
rect 5724 8372 5776 8424
rect 8300 8372 8352 8424
rect 9312 8372 9364 8424
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 13728 8372 13780 8424
rect 14832 8372 14884 8424
rect 16580 8372 16632 8424
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 17960 8372 18012 8424
rect 22008 8440 22060 8492
rect 20904 8415 20956 8424
rect 20904 8381 20938 8415
rect 20938 8381 20956 8415
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 4712 8236 4764 8288
rect 5724 8236 5776 8288
rect 11060 8236 11112 8288
rect 11336 8236 11388 8288
rect 11704 8236 11756 8288
rect 12992 8236 13044 8288
rect 15844 8236 15896 8288
rect 16212 8236 16264 8288
rect 17224 8236 17276 8288
rect 18788 8304 18840 8356
rect 19064 8304 19116 8356
rect 20904 8372 20956 8381
rect 22100 8372 22152 8424
rect 22560 8415 22612 8424
rect 22560 8381 22569 8415
rect 22569 8381 22603 8415
rect 22603 8381 22612 8415
rect 22560 8372 22612 8381
rect 24308 8440 24360 8492
rect 24860 8440 24912 8492
rect 22744 8415 22796 8424
rect 22744 8381 22753 8415
rect 22753 8381 22787 8415
rect 22787 8381 22796 8415
rect 22744 8372 22796 8381
rect 23388 8415 23440 8424
rect 23388 8381 23397 8415
rect 23397 8381 23431 8415
rect 23431 8381 23440 8415
rect 23388 8372 23440 8381
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 25780 8415 25832 8424
rect 25780 8381 25789 8415
rect 25789 8381 25823 8415
rect 25823 8381 25832 8415
rect 25780 8372 25832 8381
rect 26240 8372 26292 8424
rect 17960 8236 18012 8288
rect 20720 8304 20772 8356
rect 21916 8236 21968 8288
rect 24124 8304 24176 8356
rect 25136 8304 25188 8356
rect 26424 8372 26476 8424
rect 28540 8576 28592 8628
rect 29000 8576 29052 8628
rect 28264 8508 28316 8560
rect 28908 8508 28960 8560
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 28632 8440 28684 8492
rect 29092 8440 29144 8492
rect 28540 8415 28592 8424
rect 28540 8381 28549 8415
rect 28549 8381 28583 8415
rect 28583 8381 28592 8415
rect 28540 8372 28592 8381
rect 28816 8372 28868 8424
rect 29460 8415 29512 8424
rect 29460 8381 29469 8415
rect 29469 8381 29503 8415
rect 29503 8381 29512 8415
rect 29460 8372 29512 8381
rect 28448 8304 28500 8356
rect 22836 8236 22888 8288
rect 23020 8279 23072 8288
rect 23020 8245 23029 8279
rect 23029 8245 23063 8279
rect 23063 8245 23072 8279
rect 23020 8236 23072 8245
rect 23572 8279 23624 8288
rect 23572 8245 23581 8279
rect 23581 8245 23615 8279
rect 23615 8245 23624 8279
rect 23572 8236 23624 8245
rect 28632 8236 28684 8288
rect 29276 8347 29328 8356
rect 29276 8313 29285 8347
rect 29285 8313 29319 8347
rect 29319 8313 29328 8347
rect 29276 8304 29328 8313
rect 30656 8304 30708 8356
rect 30748 8236 30800 8288
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 12096 8134 12148 8186
rect 12160 8134 12212 8186
rect 12224 8134 12276 8186
rect 12288 8134 12340 8186
rect 12352 8134 12404 8186
rect 19870 8134 19922 8186
rect 19934 8134 19986 8186
rect 19998 8134 20050 8186
rect 20062 8134 20114 8186
rect 20126 8134 20178 8186
rect 27644 8134 27696 8186
rect 27708 8134 27760 8186
rect 27772 8134 27824 8186
rect 27836 8134 27888 8186
rect 27900 8134 27952 8186
rect 4988 8075 5040 8084
rect 4988 8041 4997 8075
rect 4997 8041 5031 8075
rect 5031 8041 5040 8075
rect 4988 8032 5040 8041
rect 4068 7964 4120 8016
rect 2964 7896 3016 7948
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 6828 7828 6880 7880
rect 8208 7896 8260 7948
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 12624 8032 12676 8084
rect 14556 8032 14608 8084
rect 10140 7896 10192 7948
rect 10692 7896 10744 7948
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 10232 7828 10284 7880
rect 11704 7896 11756 7948
rect 12072 7964 12124 8016
rect 12532 7964 12584 8016
rect 14648 8007 14700 8016
rect 14648 7973 14657 8007
rect 14657 7973 14691 8007
rect 14691 7973 14700 8007
rect 14648 7964 14700 7973
rect 15016 8032 15068 8084
rect 15292 8032 15344 8084
rect 15384 8032 15436 8084
rect 16304 8032 16356 8084
rect 16764 8032 16816 8084
rect 18512 8032 18564 8084
rect 16212 7964 16264 8016
rect 16488 8007 16540 8016
rect 16488 7973 16497 8007
rect 16497 7973 16531 8007
rect 16531 7973 16540 8007
rect 16488 7964 16540 7973
rect 16856 7964 16908 8016
rect 17592 8007 17644 8016
rect 17592 7973 17627 8007
rect 17627 7973 17644 8007
rect 17592 7964 17644 7973
rect 18144 8007 18196 8016
rect 18144 7973 18153 8007
rect 18153 7973 18187 8007
rect 18187 7973 18196 8007
rect 18144 7964 18196 7973
rect 18420 7964 18472 8016
rect 13176 7896 13228 7948
rect 13728 7896 13780 7948
rect 8576 7760 8628 7812
rect 11888 7828 11940 7880
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12992 7828 13044 7880
rect 13084 7828 13136 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 15292 7896 15344 7948
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 15660 7939 15712 7948
rect 15660 7905 15695 7939
rect 15695 7905 15712 7939
rect 15660 7896 15712 7905
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 16120 7896 16172 7948
rect 17224 7896 17276 7948
rect 16580 7828 16632 7880
rect 15384 7760 15436 7812
rect 17776 7939 17828 7948
rect 17776 7905 17785 7939
rect 17785 7905 17819 7939
rect 17819 7905 17828 7939
rect 17776 7896 17828 7905
rect 19616 8032 19668 8084
rect 20352 8075 20404 8084
rect 20352 8041 20361 8075
rect 20361 8041 20395 8075
rect 20395 8041 20404 8075
rect 20352 8032 20404 8041
rect 18972 8007 19024 8016
rect 18972 7973 18981 8007
rect 18981 7973 19015 8007
rect 19015 7973 19024 8007
rect 18972 7964 19024 7973
rect 22560 8032 22612 8084
rect 24308 8075 24360 8084
rect 24308 8041 24317 8075
rect 24317 8041 24351 8075
rect 24351 8041 24360 8075
rect 24308 8032 24360 8041
rect 20812 8007 20864 8016
rect 20812 7973 20847 8007
rect 20847 7973 20864 8007
rect 20812 7964 20864 7973
rect 19156 7939 19208 7948
rect 19156 7905 19191 7939
rect 19191 7905 19208 7939
rect 19156 7896 19208 7905
rect 20444 7896 20496 7948
rect 20628 7939 20680 7948
rect 20628 7905 20637 7939
rect 20637 7905 20671 7939
rect 20671 7905 20680 7939
rect 20628 7896 20680 7905
rect 21088 7964 21140 8016
rect 22284 7964 22336 8016
rect 17960 7828 18012 7880
rect 18052 7828 18104 7880
rect 18328 7828 18380 7880
rect 21456 7939 21508 7948
rect 21456 7905 21465 7939
rect 21465 7905 21499 7939
rect 21499 7905 21508 7939
rect 21456 7896 21508 7905
rect 21640 7896 21692 7948
rect 21824 7896 21876 7948
rect 22560 7939 22612 7948
rect 22560 7905 22569 7939
rect 22569 7905 22603 7939
rect 22603 7905 22612 7939
rect 22560 7896 22612 7905
rect 22652 7939 22704 7948
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 23572 7964 23624 8016
rect 26424 8007 26476 8016
rect 26424 7973 26433 8007
rect 26433 7973 26467 8007
rect 26467 7973 26476 8007
rect 26424 7964 26476 7973
rect 27436 7964 27488 8016
rect 28448 8032 28500 8084
rect 28540 8032 28592 8084
rect 28816 8032 28868 8084
rect 28264 8007 28316 8016
rect 28264 7973 28273 8007
rect 28273 7973 28307 8007
rect 28307 7973 28316 8007
rect 28264 7964 28316 7973
rect 29276 7964 29328 8016
rect 30748 7964 30800 8016
rect 23020 7896 23072 7948
rect 27896 7896 27948 7948
rect 21088 7828 21140 7880
rect 28080 7828 28132 7880
rect 28540 7896 28592 7948
rect 28632 7896 28684 7948
rect 29460 7896 29512 7948
rect 30840 7939 30892 7948
rect 30840 7905 30849 7939
rect 30849 7905 30883 7939
rect 30883 7905 30892 7939
rect 30840 7896 30892 7905
rect 20444 7760 20496 7812
rect 22100 7803 22152 7812
rect 22100 7769 22109 7803
rect 22109 7769 22143 7803
rect 22143 7769 22152 7803
rect 22100 7760 22152 7769
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 8668 7692 8720 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 10876 7692 10928 7744
rect 12256 7735 12308 7744
rect 12256 7701 12265 7735
rect 12265 7701 12299 7735
rect 12299 7701 12308 7735
rect 12256 7692 12308 7701
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 14004 7692 14056 7744
rect 18052 7692 18104 7744
rect 20628 7692 20680 7744
rect 21640 7735 21692 7744
rect 21640 7701 21649 7735
rect 21649 7701 21683 7735
rect 21683 7701 21692 7735
rect 21640 7692 21692 7701
rect 22284 7692 22336 7744
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 22468 7692 22520 7744
rect 23296 7692 23348 7744
rect 28632 7692 28684 7744
rect 30104 7735 30156 7744
rect 30104 7701 30113 7735
rect 30113 7701 30147 7735
rect 30147 7701 30156 7735
rect 30104 7692 30156 7701
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 11436 7590 11488 7642
rect 11500 7590 11552 7642
rect 11564 7590 11616 7642
rect 11628 7590 11680 7642
rect 11692 7590 11744 7642
rect 19210 7590 19262 7642
rect 19274 7590 19326 7642
rect 19338 7590 19390 7642
rect 19402 7590 19454 7642
rect 19466 7590 19518 7642
rect 26984 7590 27036 7642
rect 27048 7590 27100 7642
rect 27112 7590 27164 7642
rect 27176 7590 27228 7642
rect 27240 7590 27292 7642
rect 7748 7488 7800 7540
rect 11520 7488 11572 7540
rect 12532 7488 12584 7540
rect 12256 7420 12308 7472
rect 14464 7488 14516 7540
rect 14740 7488 14792 7540
rect 17592 7488 17644 7540
rect 17960 7488 18012 7540
rect 18788 7488 18840 7540
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 22560 7488 22612 7540
rect 25872 7488 25924 7540
rect 28816 7531 28868 7540
rect 28816 7497 28825 7531
rect 28825 7497 28859 7531
rect 28859 7497 28868 7531
rect 28816 7488 28868 7497
rect 16396 7420 16448 7472
rect 7564 7284 7616 7336
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 8852 7352 8904 7404
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 11888 7352 11940 7404
rect 13084 7352 13136 7404
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 17500 7395 17552 7404
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 22376 7420 22428 7472
rect 26332 7420 26384 7472
rect 30104 7488 30156 7540
rect 9772 7284 9824 7336
rect 10140 7284 10192 7336
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 10876 7327 10928 7336
rect 10876 7293 10910 7327
rect 10910 7293 10928 7327
rect 8760 7259 8812 7268
rect 8760 7225 8769 7259
rect 8769 7225 8803 7259
rect 8803 7225 8812 7259
rect 8760 7216 8812 7225
rect 10876 7284 10928 7293
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 14004 7327 14056 7336
rect 14004 7293 14038 7327
rect 14038 7293 14056 7327
rect 14004 7284 14056 7293
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 15568 7327 15620 7336
rect 15568 7293 15577 7327
rect 15577 7293 15611 7327
rect 15611 7293 15620 7327
rect 15568 7284 15620 7293
rect 15660 7284 15712 7336
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 15844 7284 15896 7293
rect 16028 7284 16080 7336
rect 16212 7284 16264 7336
rect 6828 7148 6880 7200
rect 11152 7216 11204 7268
rect 9220 7148 9272 7200
rect 11060 7148 11112 7200
rect 13820 7216 13872 7268
rect 15292 7216 15344 7268
rect 14556 7148 14608 7200
rect 18696 7284 18748 7336
rect 19340 7284 19392 7336
rect 20352 7327 20404 7336
rect 20352 7293 20361 7327
rect 20361 7293 20395 7327
rect 20395 7293 20404 7327
rect 20352 7284 20404 7293
rect 22468 7352 22520 7404
rect 24032 7352 24084 7404
rect 25228 7352 25280 7404
rect 20812 7327 20864 7336
rect 20812 7293 20821 7327
rect 20821 7293 20855 7327
rect 20855 7293 20864 7327
rect 20812 7284 20864 7293
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 20996 7216 21048 7268
rect 22836 7216 22888 7268
rect 27896 7284 27948 7336
rect 28080 7284 28132 7336
rect 28356 7284 28408 7336
rect 28632 7327 28684 7336
rect 28632 7293 28641 7327
rect 28641 7293 28675 7327
rect 28675 7293 28684 7327
rect 28632 7284 28684 7293
rect 29092 7284 29144 7336
rect 26608 7216 26660 7268
rect 17960 7148 18012 7200
rect 21548 7148 21600 7200
rect 22100 7148 22152 7200
rect 23848 7148 23900 7200
rect 24400 7148 24452 7200
rect 25228 7148 25280 7200
rect 26700 7191 26752 7200
rect 26700 7157 26709 7191
rect 26709 7157 26743 7191
rect 26743 7157 26752 7191
rect 26700 7148 26752 7157
rect 26792 7191 26844 7200
rect 26792 7157 26801 7191
rect 26801 7157 26835 7191
rect 26835 7157 26844 7191
rect 26792 7148 26844 7157
rect 28540 7148 28592 7200
rect 29920 7148 29972 7200
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 12096 7046 12148 7098
rect 12160 7046 12212 7098
rect 12224 7046 12276 7098
rect 12288 7046 12340 7098
rect 12352 7046 12404 7098
rect 19870 7046 19922 7098
rect 19934 7046 19986 7098
rect 19998 7046 20050 7098
rect 20062 7046 20114 7098
rect 20126 7046 20178 7098
rect 27644 7046 27696 7098
rect 27708 7046 27760 7098
rect 27772 7046 27824 7098
rect 27836 7046 27888 7098
rect 27900 7046 27952 7098
rect 8760 6944 8812 6996
rect 3148 6808 3200 6860
rect 4252 6876 4304 6928
rect 6828 6876 6880 6928
rect 2964 6740 3016 6792
rect 5172 6808 5224 6860
rect 7104 6808 7156 6860
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 8392 6851 8444 6860
rect 8392 6817 8410 6851
rect 8410 6817 8444 6851
rect 8392 6808 8444 6817
rect 8576 6876 8628 6928
rect 12532 6944 12584 6996
rect 15936 6944 15988 6996
rect 16120 6944 16172 6996
rect 18144 6944 18196 6996
rect 22468 6944 22520 6996
rect 22652 6944 22704 6996
rect 23020 6944 23072 6996
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 9220 6851 9272 6860
rect 9220 6817 9255 6851
rect 9255 6817 9272 6851
rect 9220 6808 9272 6817
rect 9680 6808 9732 6860
rect 11336 6876 11388 6928
rect 12348 6876 12400 6928
rect 10692 6808 10744 6860
rect 11060 6808 11112 6860
rect 11520 6808 11572 6860
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 13820 6876 13872 6928
rect 18236 6876 18288 6928
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 15568 6851 15620 6860
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 18696 6808 18748 6860
rect 8944 6672 8996 6724
rect 14464 6740 14516 6792
rect 17132 6740 17184 6792
rect 17960 6740 18012 6792
rect 9588 6672 9640 6724
rect 15292 6672 15344 6724
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 18972 6876 19024 6928
rect 19248 6851 19300 6860
rect 19248 6817 19257 6851
rect 19257 6817 19291 6851
rect 19291 6817 19300 6851
rect 19248 6808 19300 6817
rect 19340 6851 19392 6860
rect 19340 6817 19349 6851
rect 19349 6817 19383 6851
rect 19383 6817 19392 6851
rect 19340 6808 19392 6817
rect 20720 6876 20772 6928
rect 25872 6944 25924 6996
rect 26516 6944 26568 6996
rect 19616 6808 19668 6860
rect 21180 6808 21232 6860
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 21364 6808 21416 6860
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 24308 6919 24360 6928
rect 24308 6885 24317 6919
rect 24317 6885 24351 6919
rect 24351 6885 24360 6919
rect 24308 6876 24360 6885
rect 26332 6876 26384 6928
rect 23296 6851 23348 6860
rect 23296 6817 23305 6851
rect 23305 6817 23339 6851
rect 23339 6817 23348 6851
rect 23296 6808 23348 6817
rect 23480 6851 23532 6860
rect 23480 6817 23489 6851
rect 23489 6817 23523 6851
rect 23523 6817 23532 6851
rect 23480 6808 23532 6817
rect 23940 6851 23992 6860
rect 23940 6817 23949 6851
rect 23949 6817 23983 6851
rect 23983 6817 23992 6851
rect 23940 6808 23992 6817
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 19156 6740 19208 6792
rect 18696 6672 18748 6724
rect 22560 6740 22612 6792
rect 3516 6604 3568 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 8024 6604 8076 6656
rect 11336 6604 11388 6656
rect 12164 6604 12216 6656
rect 15936 6647 15988 6656
rect 15936 6613 15945 6647
rect 15945 6613 15979 6647
rect 15979 6613 15988 6647
rect 15936 6604 15988 6613
rect 18972 6647 19024 6656
rect 18972 6613 18981 6647
rect 18981 6613 19015 6647
rect 19015 6613 19024 6647
rect 18972 6604 19024 6613
rect 19340 6604 19392 6656
rect 21732 6672 21784 6724
rect 22284 6604 22336 6656
rect 23296 6672 23348 6724
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 23664 6672 23716 6724
rect 24584 6808 24636 6860
rect 22560 6604 22612 6656
rect 23480 6647 23532 6656
rect 23480 6613 23489 6647
rect 23489 6613 23523 6647
rect 23523 6613 23532 6647
rect 23480 6604 23532 6613
rect 24492 6672 24544 6724
rect 25044 6851 25096 6860
rect 25044 6817 25053 6851
rect 25053 6817 25087 6851
rect 25087 6817 25096 6851
rect 25044 6808 25096 6817
rect 25228 6851 25280 6860
rect 25228 6817 25237 6851
rect 25237 6817 25271 6851
rect 25271 6817 25280 6851
rect 25228 6808 25280 6817
rect 26792 6808 26844 6860
rect 29000 6808 29052 6860
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 25504 6647 25556 6656
rect 25504 6613 25513 6647
rect 25513 6613 25547 6647
rect 25547 6613 25556 6647
rect 25504 6604 25556 6613
rect 26240 6740 26292 6792
rect 29184 6783 29236 6792
rect 29184 6749 29193 6783
rect 29193 6749 29227 6783
rect 29227 6749 29236 6783
rect 29184 6740 29236 6749
rect 29644 6851 29696 6860
rect 29644 6817 29654 6851
rect 29654 6817 29688 6851
rect 29688 6817 29696 6851
rect 29644 6808 29696 6817
rect 29828 6851 29880 6860
rect 29828 6817 29837 6851
rect 29837 6817 29871 6851
rect 29871 6817 29880 6851
rect 29828 6808 29880 6817
rect 30104 6808 30156 6860
rect 30380 6808 30432 6860
rect 30656 6851 30708 6860
rect 30656 6817 30665 6851
rect 30665 6817 30699 6851
rect 30699 6817 30708 6851
rect 30656 6808 30708 6817
rect 26332 6604 26384 6656
rect 26424 6647 26476 6656
rect 26424 6613 26433 6647
rect 26433 6613 26467 6647
rect 26467 6613 26476 6647
rect 26424 6604 26476 6613
rect 26608 6715 26660 6724
rect 26608 6681 26617 6715
rect 26617 6681 26651 6715
rect 26651 6681 26660 6715
rect 26608 6672 26660 6681
rect 27436 6647 27488 6656
rect 27436 6613 27445 6647
rect 27445 6613 27479 6647
rect 27479 6613 27488 6647
rect 27436 6604 27488 6613
rect 30196 6715 30248 6724
rect 30196 6681 30205 6715
rect 30205 6681 30239 6715
rect 30239 6681 30248 6715
rect 30196 6672 30248 6681
rect 30380 6604 30432 6656
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 11436 6502 11488 6554
rect 11500 6502 11552 6554
rect 11564 6502 11616 6554
rect 11628 6502 11680 6554
rect 11692 6502 11744 6554
rect 19210 6502 19262 6554
rect 19274 6502 19326 6554
rect 19338 6502 19390 6554
rect 19402 6502 19454 6554
rect 19466 6502 19518 6554
rect 26984 6502 27036 6554
rect 27048 6502 27100 6554
rect 27112 6502 27164 6554
rect 27176 6502 27228 6554
rect 27240 6502 27292 6554
rect 8392 6400 8444 6452
rect 9588 6400 9640 6452
rect 3516 6332 3568 6384
rect 11152 6400 11204 6452
rect 12164 6400 12216 6452
rect 12348 6332 12400 6384
rect 2044 6128 2096 6180
rect 6828 6196 6880 6248
rect 7932 6239 7984 6248
rect 7932 6205 7941 6239
rect 7941 6205 7975 6239
rect 7975 6205 7984 6239
rect 7932 6196 7984 6205
rect 8024 6239 8076 6248
rect 8024 6205 8033 6239
rect 8033 6205 8067 6239
rect 8067 6205 8076 6239
rect 8024 6196 8076 6205
rect 2872 6060 2924 6112
rect 4252 6060 4304 6112
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 5172 6060 5224 6112
rect 7104 6171 7156 6180
rect 7104 6137 7113 6171
rect 7113 6137 7147 6171
rect 7147 6137 7156 6171
rect 7104 6128 7156 6137
rect 8116 6060 8168 6112
rect 8392 6060 8444 6112
rect 8668 6128 8720 6180
rect 12440 6264 12492 6316
rect 12164 6239 12216 6248
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 11796 6128 11848 6180
rect 12532 6196 12584 6248
rect 12808 6196 12860 6248
rect 18788 6400 18840 6452
rect 19524 6400 19576 6452
rect 15016 6264 15068 6316
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 17408 6264 17460 6316
rect 13176 6128 13228 6180
rect 13268 6128 13320 6180
rect 15568 6196 15620 6248
rect 18880 6264 18932 6316
rect 19524 6264 19576 6316
rect 19156 6239 19208 6248
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 17224 6128 17276 6180
rect 17316 6128 17368 6180
rect 17500 6128 17552 6180
rect 18144 6171 18196 6180
rect 18144 6137 18153 6171
rect 18153 6137 18187 6171
rect 18187 6137 18196 6171
rect 18144 6128 18196 6137
rect 18696 6060 18748 6112
rect 19156 6205 19170 6239
rect 19170 6205 19204 6239
rect 19204 6205 19208 6239
rect 19156 6196 19208 6205
rect 19616 6239 19668 6248
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 19708 6239 19760 6248
rect 19708 6205 19717 6239
rect 19717 6205 19751 6239
rect 19751 6205 19760 6239
rect 19708 6196 19760 6205
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 22008 6400 22060 6452
rect 22560 6443 22612 6452
rect 22560 6409 22569 6443
rect 22569 6409 22603 6443
rect 22603 6409 22612 6443
rect 22560 6400 22612 6409
rect 23572 6400 23624 6452
rect 26700 6400 26752 6452
rect 29644 6443 29696 6452
rect 29644 6409 29653 6443
rect 29653 6409 29687 6443
rect 29687 6409 29696 6443
rect 29644 6400 29696 6409
rect 29828 6443 29880 6452
rect 29828 6409 29837 6443
rect 29837 6409 29871 6443
rect 29871 6409 29880 6443
rect 29828 6400 29880 6409
rect 30104 6443 30156 6452
rect 30104 6409 30113 6443
rect 30113 6409 30147 6443
rect 30147 6409 30156 6443
rect 30104 6400 30156 6409
rect 22284 6332 22336 6384
rect 23020 6375 23072 6384
rect 23020 6341 23029 6375
rect 23029 6341 23063 6375
rect 23063 6341 23072 6375
rect 23020 6332 23072 6341
rect 23112 6332 23164 6384
rect 23756 6332 23808 6384
rect 20352 6239 20404 6248
rect 20352 6205 20361 6239
rect 20361 6205 20395 6239
rect 20395 6205 20404 6239
rect 20352 6196 20404 6205
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22192 6196 22244 6248
rect 22468 6196 22520 6248
rect 18972 6171 19024 6180
rect 18972 6137 18981 6171
rect 18981 6137 19015 6171
rect 19015 6137 19024 6171
rect 18972 6128 19024 6137
rect 19064 6171 19116 6180
rect 19064 6137 19073 6171
rect 19073 6137 19107 6171
rect 19107 6137 19116 6171
rect 19064 6128 19116 6137
rect 19248 6128 19300 6180
rect 19156 6060 19208 6112
rect 21732 6128 21784 6180
rect 21824 6171 21876 6180
rect 21824 6137 21833 6171
rect 21833 6137 21867 6171
rect 21867 6137 21876 6171
rect 21824 6128 21876 6137
rect 22376 6128 22428 6180
rect 25136 6128 25188 6180
rect 26148 6264 26200 6316
rect 26332 6239 26384 6248
rect 26332 6205 26341 6239
rect 26341 6205 26375 6239
rect 26375 6205 26384 6239
rect 26332 6196 26384 6205
rect 27436 6196 27488 6248
rect 26424 6128 26476 6180
rect 29920 6239 29972 6248
rect 29920 6205 29929 6239
rect 29929 6205 29963 6239
rect 29963 6205 29972 6239
rect 29920 6196 29972 6205
rect 30656 6196 30708 6248
rect 30380 6128 30432 6180
rect 19616 6060 19668 6112
rect 23112 6060 23164 6112
rect 23204 6060 23256 6112
rect 23848 6060 23900 6112
rect 26700 6103 26752 6112
rect 26700 6069 26709 6103
rect 26709 6069 26743 6103
rect 26743 6069 26752 6103
rect 26700 6060 26752 6069
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 12096 5958 12148 6010
rect 12160 5958 12212 6010
rect 12224 5958 12276 6010
rect 12288 5958 12340 6010
rect 12352 5958 12404 6010
rect 19870 5958 19922 6010
rect 19934 5958 19986 6010
rect 19998 5958 20050 6010
rect 20062 5958 20114 6010
rect 20126 5958 20178 6010
rect 27644 5958 27696 6010
rect 27708 5958 27760 6010
rect 27772 5958 27824 6010
rect 27836 5958 27888 6010
rect 27900 5958 27952 6010
rect 3148 5856 3200 5908
rect 2872 5763 2924 5772
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 4896 5856 4948 5908
rect 4068 5788 4120 5840
rect 4160 5788 4212 5840
rect 4252 5788 4304 5840
rect 8668 5856 8720 5908
rect 8760 5856 8812 5908
rect 8392 5788 8444 5840
rect 9588 5856 9640 5908
rect 2320 5652 2372 5704
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 3516 5652 3568 5704
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 8576 5720 8628 5772
rect 6276 5652 6328 5704
rect 3332 5516 3384 5568
rect 4712 5584 4764 5636
rect 5908 5584 5960 5636
rect 8760 5763 8812 5772
rect 8760 5729 8769 5763
rect 8769 5729 8803 5763
rect 8803 5729 8812 5763
rect 8760 5720 8812 5729
rect 12992 5788 13044 5840
rect 13636 5788 13688 5840
rect 9404 5763 9456 5772
rect 9404 5729 9413 5763
rect 9413 5729 9447 5763
rect 9447 5729 9456 5763
rect 9404 5720 9456 5729
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 9588 5763 9640 5772
rect 9588 5729 9597 5763
rect 9597 5729 9631 5763
rect 9631 5729 9640 5763
rect 9588 5720 9640 5729
rect 9220 5652 9272 5704
rect 10048 5720 10100 5772
rect 11244 5720 11296 5772
rect 13268 5763 13320 5772
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 13176 5652 13228 5704
rect 15844 5856 15896 5908
rect 19708 5856 19760 5908
rect 19800 5856 19852 5908
rect 20352 5856 20404 5908
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 19616 5788 19668 5840
rect 22928 5856 22980 5908
rect 23480 5856 23532 5908
rect 18972 5652 19024 5704
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 9404 5584 9456 5636
rect 12900 5584 12952 5636
rect 16488 5584 16540 5636
rect 19156 5695 19208 5704
rect 19156 5661 19165 5695
rect 19165 5661 19199 5695
rect 19199 5661 19208 5695
rect 22008 5720 22060 5772
rect 22100 5763 22152 5772
rect 22100 5729 22109 5763
rect 22109 5729 22143 5763
rect 22143 5729 22152 5763
rect 22100 5720 22152 5729
rect 19156 5652 19208 5661
rect 5540 5516 5592 5525
rect 9128 5516 9180 5568
rect 12164 5516 12216 5568
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 18696 5559 18748 5568
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 19248 5584 19300 5636
rect 19340 5584 19392 5636
rect 21824 5652 21876 5704
rect 22284 5788 22336 5840
rect 22376 5831 22428 5840
rect 22376 5797 22385 5831
rect 22385 5797 22419 5831
rect 22419 5797 22428 5831
rect 22376 5788 22428 5797
rect 23020 5788 23072 5840
rect 22376 5652 22428 5704
rect 22652 5763 22704 5772
rect 22652 5729 22661 5763
rect 22661 5729 22695 5763
rect 22695 5729 22704 5763
rect 22652 5720 22704 5729
rect 23204 5720 23256 5772
rect 22928 5695 22980 5704
rect 22928 5661 22937 5695
rect 22937 5661 22971 5695
rect 22971 5661 22980 5695
rect 22928 5652 22980 5661
rect 23664 5788 23716 5840
rect 23940 5788 23992 5840
rect 23572 5763 23624 5772
rect 23572 5729 23581 5763
rect 23581 5729 23615 5763
rect 23615 5729 23624 5763
rect 23572 5720 23624 5729
rect 24032 5763 24084 5772
rect 24032 5729 24041 5763
rect 24041 5729 24075 5763
rect 24075 5729 24084 5763
rect 24032 5720 24084 5729
rect 24952 5788 25004 5840
rect 26608 5788 26660 5840
rect 24400 5763 24452 5772
rect 24400 5729 24409 5763
rect 24409 5729 24443 5763
rect 24443 5729 24452 5763
rect 24400 5720 24452 5729
rect 24676 5720 24728 5772
rect 25412 5763 25464 5772
rect 25412 5729 25421 5763
rect 25421 5729 25455 5763
rect 25455 5729 25464 5763
rect 25412 5720 25464 5729
rect 26056 5720 26108 5772
rect 28172 5720 28224 5772
rect 28632 5788 28684 5840
rect 29000 5788 29052 5840
rect 28448 5720 28500 5772
rect 28724 5720 28776 5772
rect 21364 5516 21416 5568
rect 23480 5584 23532 5636
rect 23940 5584 23992 5636
rect 21732 5516 21784 5568
rect 22192 5516 22244 5568
rect 22744 5559 22796 5568
rect 22744 5525 22753 5559
rect 22753 5525 22787 5559
rect 22787 5525 22796 5559
rect 22744 5516 22796 5525
rect 22928 5516 22980 5568
rect 23204 5559 23256 5568
rect 23204 5525 23213 5559
rect 23213 5525 23247 5559
rect 23247 5525 23256 5559
rect 23204 5516 23256 5525
rect 23296 5559 23348 5568
rect 23296 5525 23305 5559
rect 23305 5525 23339 5559
rect 23339 5525 23348 5559
rect 23296 5516 23348 5525
rect 23756 5559 23808 5568
rect 23756 5525 23765 5559
rect 23765 5525 23799 5559
rect 23799 5525 23808 5559
rect 23756 5516 23808 5525
rect 24216 5695 24268 5704
rect 24216 5661 24225 5695
rect 24225 5661 24259 5695
rect 24259 5661 24268 5695
rect 24216 5652 24268 5661
rect 28540 5627 28592 5636
rect 28540 5593 28549 5627
rect 28549 5593 28583 5627
rect 28583 5593 28592 5627
rect 28540 5584 28592 5593
rect 24308 5516 24360 5568
rect 29092 5559 29144 5568
rect 29092 5525 29101 5559
rect 29101 5525 29135 5559
rect 29135 5525 29144 5559
rect 29092 5516 29144 5525
rect 29552 5559 29604 5568
rect 29552 5525 29561 5559
rect 29561 5525 29595 5559
rect 29595 5525 29604 5559
rect 29552 5516 29604 5525
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 11436 5414 11488 5466
rect 11500 5414 11552 5466
rect 11564 5414 11616 5466
rect 11628 5414 11680 5466
rect 11692 5414 11744 5466
rect 19210 5414 19262 5466
rect 19274 5414 19326 5466
rect 19338 5414 19390 5466
rect 19402 5414 19454 5466
rect 19466 5414 19518 5466
rect 26984 5414 27036 5466
rect 27048 5414 27100 5466
rect 27112 5414 27164 5466
rect 27176 5414 27228 5466
rect 27240 5414 27292 5466
rect 3424 5312 3476 5364
rect 3608 5312 3660 5364
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 5632 5312 5684 5364
rect 11336 5312 11388 5364
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 12532 5355 12584 5364
rect 12532 5321 12550 5355
rect 12550 5321 12584 5355
rect 12532 5312 12584 5321
rect 13084 5312 13136 5364
rect 13912 5355 13964 5364
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 14464 5312 14516 5364
rect 21732 5312 21784 5364
rect 22284 5312 22336 5364
rect 23756 5312 23808 5364
rect 24216 5312 24268 5364
rect 24768 5312 24820 5364
rect 28172 5355 28224 5364
rect 28172 5321 28181 5355
rect 28181 5321 28215 5355
rect 28215 5321 28224 5355
rect 28172 5312 28224 5321
rect 7932 5244 7984 5296
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 6276 5176 6328 5228
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 4712 5108 4764 5160
rect 1952 5083 2004 5092
rect 1952 5049 1986 5083
rect 1986 5049 2004 5083
rect 1952 5040 2004 5049
rect 2044 4972 2096 5024
rect 3240 5040 3292 5092
rect 3792 5040 3844 5092
rect 5908 5151 5960 5160
rect 5908 5117 5942 5151
rect 5942 5117 5960 5151
rect 5908 5108 5960 5117
rect 6092 5151 6144 5160
rect 6092 5117 6101 5151
rect 6101 5117 6135 5151
rect 6135 5117 6144 5151
rect 6092 5108 6144 5117
rect 8116 5151 8168 5160
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 9128 5151 9180 5160
rect 9128 5117 9137 5151
rect 9137 5117 9171 5151
rect 9171 5117 9180 5151
rect 9128 5108 9180 5117
rect 11152 5151 11204 5160
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 12992 5176 13044 5228
rect 9496 5040 9548 5092
rect 12440 5108 12492 5160
rect 15200 5176 15252 5228
rect 13636 5108 13688 5160
rect 14372 5108 14424 5160
rect 18328 5244 18380 5296
rect 21548 5244 21600 5296
rect 21456 5176 21508 5228
rect 22008 5287 22060 5296
rect 22008 5253 22017 5287
rect 22017 5253 22051 5287
rect 22051 5253 22060 5287
rect 22008 5244 22060 5253
rect 23112 5244 23164 5296
rect 23664 5287 23716 5296
rect 23664 5253 23673 5287
rect 23673 5253 23707 5287
rect 23707 5253 23716 5287
rect 23664 5244 23716 5253
rect 24676 5244 24728 5296
rect 23204 5176 23256 5228
rect 24216 5219 24268 5228
rect 18604 5108 18656 5160
rect 22100 5108 22152 5160
rect 22744 5151 22796 5160
rect 22744 5117 22753 5151
rect 22753 5117 22787 5151
rect 22787 5117 22796 5151
rect 22744 5108 22796 5117
rect 12808 5040 12860 5092
rect 14740 5040 14792 5092
rect 21548 5083 21600 5092
rect 21548 5049 21557 5083
rect 21557 5049 21591 5083
rect 21591 5049 21600 5083
rect 21548 5040 21600 5049
rect 21640 5040 21692 5092
rect 22376 5040 22428 5092
rect 22928 5108 22980 5160
rect 24216 5185 24225 5219
rect 24225 5185 24259 5219
rect 24259 5185 24268 5219
rect 24216 5176 24268 5185
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 25872 5287 25924 5296
rect 25872 5253 25881 5287
rect 25881 5253 25915 5287
rect 25915 5253 25924 5287
rect 25872 5244 25924 5253
rect 29552 5312 29604 5364
rect 26148 5219 26200 5228
rect 26148 5185 26157 5219
rect 26157 5185 26191 5219
rect 26191 5185 26200 5219
rect 26148 5176 26200 5185
rect 23848 5151 23900 5160
rect 23848 5117 23857 5151
rect 23857 5117 23891 5151
rect 23891 5117 23900 5151
rect 23848 5108 23900 5117
rect 23940 5108 23992 5160
rect 24124 5108 24176 5160
rect 25044 5151 25096 5160
rect 25044 5117 25053 5151
rect 25053 5117 25087 5151
rect 25087 5117 25096 5151
rect 25044 5108 25096 5117
rect 25228 5108 25280 5160
rect 3332 4972 3384 5024
rect 3976 4972 4028 5024
rect 5816 4972 5868 5024
rect 7840 4972 7892 5024
rect 8668 4972 8720 5024
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 10968 4972 11020 5024
rect 11244 5015 11296 5024
rect 11244 4981 11253 5015
rect 11253 4981 11287 5015
rect 11287 4981 11296 5015
rect 11244 4972 11296 4981
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 11888 4972 11940 5024
rect 12992 4972 13044 5024
rect 13820 4972 13872 5024
rect 14280 5015 14332 5024
rect 14280 4981 14307 5015
rect 14307 4981 14332 5015
rect 14280 4972 14332 4981
rect 17316 4972 17368 5024
rect 23204 5083 23256 5092
rect 23204 5049 23213 5083
rect 23213 5049 23247 5083
rect 23247 5049 23256 5083
rect 23204 5040 23256 5049
rect 23388 5040 23440 5092
rect 27160 5108 27212 5160
rect 25872 5040 25924 5092
rect 23480 4972 23532 5024
rect 23572 4972 23624 5024
rect 27988 5151 28040 5160
rect 27988 5117 27997 5151
rect 27997 5117 28031 5151
rect 28031 5117 28040 5151
rect 27988 5108 28040 5117
rect 28264 5108 28316 5160
rect 28724 5108 28776 5160
rect 29000 5244 29052 5296
rect 28080 5040 28132 5092
rect 28172 4972 28224 5024
rect 28632 5015 28684 5024
rect 28632 4981 28641 5015
rect 28641 4981 28675 5015
rect 28675 4981 28684 5015
rect 28632 4972 28684 4981
rect 30932 5015 30984 5024
rect 30932 4981 30941 5015
rect 30941 4981 30975 5015
rect 30975 4981 30984 5015
rect 30932 4972 30984 4981
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 12096 4870 12148 4922
rect 12160 4870 12212 4922
rect 12224 4870 12276 4922
rect 12288 4870 12340 4922
rect 12352 4870 12404 4922
rect 19870 4870 19922 4922
rect 19934 4870 19986 4922
rect 19998 4870 20050 4922
rect 20062 4870 20114 4922
rect 20126 4870 20178 4922
rect 27644 4870 27696 4922
rect 27708 4870 27760 4922
rect 27772 4870 27824 4922
rect 27836 4870 27888 4922
rect 27900 4870 27952 4922
rect 1952 4768 2004 4820
rect 3424 4768 3476 4820
rect 3516 4768 3568 4820
rect 3976 4768 4028 4820
rect 9496 4768 9548 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 2044 4675 2096 4684
rect 2044 4641 2053 4675
rect 2053 4641 2087 4675
rect 2087 4641 2096 4675
rect 2044 4632 2096 4641
rect 4252 4700 4304 4752
rect 4896 4743 4948 4752
rect 4896 4709 4905 4743
rect 4905 4709 4939 4743
rect 4939 4709 4948 4743
rect 4896 4700 4948 4709
rect 8944 4700 8996 4752
rect 11244 4743 11296 4752
rect 11244 4709 11278 4743
rect 11278 4709 11296 4743
rect 11244 4700 11296 4709
rect 11888 4700 11940 4752
rect 12808 4743 12860 4752
rect 12808 4709 12817 4743
rect 12817 4709 12851 4743
rect 12851 4709 12860 4743
rect 12808 4700 12860 4709
rect 14372 4811 14424 4820
rect 14372 4777 14381 4811
rect 14381 4777 14415 4811
rect 14415 4777 14424 4811
rect 14372 4768 14424 4777
rect 16120 4768 16172 4820
rect 16488 4768 16540 4820
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 18696 4768 18748 4820
rect 14280 4700 14332 4752
rect 14740 4743 14792 4752
rect 14740 4709 14749 4743
rect 14749 4709 14783 4743
rect 14783 4709 14792 4743
rect 14740 4700 14792 4709
rect 3792 4675 3844 4684
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 3792 4641 3801 4675
rect 3801 4641 3835 4675
rect 3835 4641 3844 4675
rect 3792 4632 3844 4641
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 12900 4675 12952 4684
rect 12900 4641 12909 4675
rect 12909 4641 12943 4675
rect 12943 4641 12952 4675
rect 12900 4632 12952 4641
rect 12992 4632 13044 4684
rect 13636 4632 13688 4684
rect 5540 4564 5592 4616
rect 14372 4632 14424 4684
rect 17408 4700 17460 4752
rect 19616 4768 19668 4820
rect 22928 4768 22980 4820
rect 23020 4768 23072 4820
rect 23388 4811 23440 4820
rect 23388 4777 23397 4811
rect 23397 4777 23431 4811
rect 23431 4777 23440 4811
rect 23388 4768 23440 4777
rect 15476 4632 15528 4684
rect 16120 4675 16172 4684
rect 16120 4641 16129 4675
rect 16129 4641 16163 4675
rect 16163 4641 16172 4675
rect 16120 4632 16172 4641
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 15016 4564 15068 4616
rect 16580 4632 16632 4684
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 17500 4675 17552 4684
rect 17500 4641 17509 4675
rect 17509 4641 17543 4675
rect 17543 4641 17552 4675
rect 17500 4632 17552 4641
rect 23756 4700 23808 4752
rect 27160 4811 27212 4820
rect 27160 4777 27187 4811
rect 27187 4777 27212 4811
rect 24032 4743 24084 4752
rect 24032 4709 24041 4743
rect 24041 4709 24075 4743
rect 24075 4709 24084 4743
rect 24032 4700 24084 4709
rect 17960 4632 18012 4684
rect 18144 4632 18196 4684
rect 17224 4564 17276 4616
rect 18512 4564 18564 4616
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 20628 4632 20680 4684
rect 22652 4675 22704 4684
rect 22652 4641 22661 4675
rect 22661 4641 22695 4675
rect 22695 4641 22704 4675
rect 22652 4632 22704 4641
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 3608 4496 3660 4548
rect 12532 4496 12584 4548
rect 14464 4496 14516 4548
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 23296 4632 23348 4684
rect 23480 4564 23532 4616
rect 23664 4632 23716 4684
rect 24492 4700 24544 4752
rect 25044 4700 25096 4752
rect 27160 4768 27212 4777
rect 28540 4768 28592 4820
rect 28264 4743 28316 4752
rect 28264 4709 28291 4743
rect 28291 4709 28316 4743
rect 24216 4632 24268 4684
rect 25228 4675 25280 4684
rect 25228 4641 25237 4675
rect 25237 4641 25271 4675
rect 25271 4641 25280 4675
rect 25228 4632 25280 4641
rect 25964 4632 26016 4684
rect 28264 4700 28316 4709
rect 28448 4743 28500 4752
rect 28448 4709 28457 4743
rect 28457 4709 28491 4743
rect 28491 4709 28500 4743
rect 28448 4700 28500 4709
rect 29092 4700 29144 4752
rect 22376 4539 22428 4548
rect 22376 4505 22385 4539
rect 22385 4505 22419 4539
rect 22419 4505 22428 4539
rect 22376 4496 22428 4505
rect 24308 4564 24360 4616
rect 2688 4471 2740 4480
rect 2688 4437 2697 4471
rect 2697 4437 2731 4471
rect 2731 4437 2740 4471
rect 2688 4428 2740 4437
rect 4068 4471 4120 4480
rect 4068 4437 4077 4471
rect 4077 4437 4111 4471
rect 4111 4437 4120 4471
rect 4068 4428 4120 4437
rect 4528 4471 4580 4480
rect 4528 4437 4537 4471
rect 4537 4437 4571 4471
rect 4571 4437 4580 4471
rect 4528 4428 4580 4437
rect 4712 4471 4764 4480
rect 4712 4437 4721 4471
rect 4721 4437 4755 4471
rect 4755 4437 4764 4471
rect 4712 4428 4764 4437
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 12624 4471 12676 4480
rect 12624 4437 12633 4471
rect 12633 4437 12667 4471
rect 12667 4437 12676 4471
rect 12624 4428 12676 4437
rect 14372 4428 14424 4480
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 14556 4428 14608 4437
rect 14924 4428 14976 4480
rect 16304 4428 16356 4480
rect 16948 4428 17000 4480
rect 17868 4428 17920 4480
rect 19432 4428 19484 4480
rect 22008 4428 22060 4480
rect 24032 4496 24084 4548
rect 24952 4496 25004 4548
rect 26056 4607 26108 4616
rect 26056 4573 26065 4607
rect 26065 4573 26099 4607
rect 26099 4573 26108 4607
rect 26056 4564 26108 4573
rect 28908 4632 28960 4684
rect 30932 4632 30984 4684
rect 24676 4471 24728 4480
rect 24676 4437 24685 4471
rect 24685 4437 24719 4471
rect 24719 4437 24728 4471
rect 24676 4428 24728 4437
rect 24768 4428 24820 4480
rect 26884 4428 26936 4480
rect 28448 4496 28500 4548
rect 27620 4471 27672 4480
rect 27620 4437 27629 4471
rect 27629 4437 27663 4471
rect 27663 4437 27672 4471
rect 27620 4428 27672 4437
rect 28172 4428 28224 4480
rect 29000 4428 29052 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 11436 4326 11488 4378
rect 11500 4326 11552 4378
rect 11564 4326 11616 4378
rect 11628 4326 11680 4378
rect 11692 4326 11744 4378
rect 19210 4326 19262 4378
rect 19274 4326 19326 4378
rect 19338 4326 19390 4378
rect 19402 4326 19454 4378
rect 19466 4326 19518 4378
rect 26984 4326 27036 4378
rect 27048 4326 27100 4378
rect 27112 4326 27164 4378
rect 27176 4326 27228 4378
rect 27240 4326 27292 4378
rect 2044 4063 2096 4072
rect 2044 4029 2053 4063
rect 2053 4029 2087 4063
rect 2087 4029 2096 4063
rect 2044 4020 2096 4029
rect 2688 4199 2740 4208
rect 2688 4165 2697 4199
rect 2697 4165 2731 4199
rect 2731 4165 2740 4199
rect 2688 4156 2740 4165
rect 4068 4224 4120 4276
rect 3424 4156 3476 4208
rect 4252 4156 4304 4208
rect 4528 4199 4580 4208
rect 4528 4165 4537 4199
rect 4537 4165 4571 4199
rect 4571 4165 4580 4199
rect 4528 4156 4580 4165
rect 4712 4156 4764 4208
rect 2504 4088 2556 4140
rect 4068 4088 4120 4140
rect 5540 4088 5592 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 8852 4224 8904 4276
rect 14556 4224 14608 4276
rect 16212 4224 16264 4276
rect 6184 4088 6236 4097
rect 2872 4020 2924 4072
rect 1768 3884 1820 3936
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 3332 4020 3384 4072
rect 4896 4020 4948 4072
rect 4988 4063 5040 4072
rect 4988 4029 4997 4063
rect 4997 4029 5031 4063
rect 5031 4029 5040 4063
rect 4988 4020 5040 4029
rect 6000 4063 6052 4072
rect 6000 4029 6034 4063
rect 6034 4029 6052 4063
rect 6000 4020 6052 4029
rect 9128 4156 9180 4208
rect 18144 4267 18196 4276
rect 18144 4233 18153 4267
rect 18153 4233 18187 4267
rect 18187 4233 18196 4267
rect 18144 4224 18196 4233
rect 9496 4088 9548 4140
rect 18604 4156 18656 4208
rect 17408 4088 17460 4140
rect 18512 4088 18564 4140
rect 19616 4224 19668 4276
rect 23480 4224 23532 4276
rect 24492 4224 24544 4276
rect 27620 4224 27672 4276
rect 22192 4156 22244 4208
rect 3976 3927 4028 3936
rect 3976 3893 3985 3927
rect 3985 3893 4019 3927
rect 4019 3893 4028 3927
rect 3976 3884 4028 3893
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 4896 3884 4948 3936
rect 6000 3884 6052 3936
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 8668 3927 8720 3936
rect 8668 3893 8677 3927
rect 8677 3893 8711 3927
rect 8711 3893 8720 3927
rect 8668 3884 8720 3893
rect 9588 4020 9640 4072
rect 11152 4020 11204 4072
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 13820 4063 13872 4072
rect 13820 4029 13854 4063
rect 13854 4029 13872 4063
rect 13820 4020 13872 4029
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 17868 4063 17920 4072
rect 17868 4029 17876 4063
rect 17876 4029 17910 4063
rect 17910 4029 17920 4063
rect 17868 4020 17920 4029
rect 18236 4063 18288 4072
rect 18236 4029 18245 4063
rect 18245 4029 18279 4063
rect 18279 4029 18288 4063
rect 18236 4020 18288 4029
rect 18420 4063 18472 4072
rect 18420 4029 18429 4063
rect 18429 4029 18463 4063
rect 18463 4029 18472 4063
rect 18420 4020 18472 4029
rect 18604 4020 18656 4072
rect 18972 4088 19024 4140
rect 11796 3952 11848 4004
rect 16120 3952 16172 4004
rect 9312 3884 9364 3936
rect 12624 3884 12676 3936
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 16764 3884 16816 3893
rect 18972 3995 19024 4004
rect 18972 3961 18981 3995
rect 18981 3961 19015 3995
rect 19015 3961 19024 3995
rect 18972 3952 19024 3961
rect 19064 3995 19116 4004
rect 19064 3961 19073 3995
rect 19073 3961 19107 3995
rect 19107 3961 19116 3995
rect 19064 3952 19116 3961
rect 17960 3884 18012 3936
rect 22744 4088 22796 4140
rect 22836 4088 22888 4140
rect 24768 4088 24820 4140
rect 26884 4088 26936 4140
rect 22100 4020 22152 4072
rect 23756 4020 23808 4072
rect 25228 4020 25280 4072
rect 27252 4063 27304 4072
rect 27252 4029 27261 4063
rect 27261 4029 27295 4063
rect 27295 4029 27304 4063
rect 27252 4020 27304 4029
rect 27988 4020 28040 4072
rect 29000 4063 29052 4072
rect 29000 4029 29009 4063
rect 29009 4029 29043 4063
rect 29043 4029 29052 4063
rect 29000 4020 29052 4029
rect 27896 3952 27948 4004
rect 28632 3995 28684 4004
rect 28632 3961 28641 3995
rect 28641 3961 28675 3995
rect 28675 3961 28684 3995
rect 28632 3952 28684 3961
rect 28908 3884 28960 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 12096 3782 12148 3834
rect 12160 3782 12212 3834
rect 12224 3782 12276 3834
rect 12288 3782 12340 3834
rect 12352 3782 12404 3834
rect 19870 3782 19922 3834
rect 19934 3782 19986 3834
rect 19998 3782 20050 3834
rect 20062 3782 20114 3834
rect 20126 3782 20178 3834
rect 27644 3782 27696 3834
rect 27708 3782 27760 3834
rect 27772 3782 27824 3834
rect 27836 3782 27888 3834
rect 27900 3782 27952 3834
rect 3332 3680 3384 3732
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 2688 3612 2740 3664
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 3424 3544 3476 3596
rect 5080 3612 5132 3664
rect 10968 3612 11020 3664
rect 3976 3476 4028 3528
rect 8484 3544 8536 3596
rect 17132 3612 17184 3664
rect 18236 3680 18288 3732
rect 18972 3680 19024 3732
rect 21548 3680 21600 3732
rect 22376 3680 22428 3732
rect 18420 3612 18472 3664
rect 14924 3544 14976 3596
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 16488 3587 16540 3596
rect 16488 3553 16497 3587
rect 16497 3553 16531 3587
rect 16531 3553 16540 3587
rect 16488 3544 16540 3553
rect 16764 3544 16816 3596
rect 5632 3476 5684 3528
rect 7932 3476 7984 3528
rect 8760 3476 8812 3528
rect 10508 3476 10560 3528
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 18880 3544 18932 3596
rect 22100 3655 22152 3664
rect 22100 3621 22109 3655
rect 22109 3621 22143 3655
rect 22143 3621 22152 3655
rect 22100 3612 22152 3621
rect 21548 3476 21600 3528
rect 8944 3408 8996 3460
rect 4988 3340 5040 3392
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 8484 3340 8536 3392
rect 11796 3408 11848 3460
rect 11060 3340 11112 3392
rect 14372 3340 14424 3392
rect 20904 3340 20956 3392
rect 22192 3587 22244 3596
rect 22192 3553 22201 3587
rect 22201 3553 22235 3587
rect 22235 3553 22244 3587
rect 22192 3544 22244 3553
rect 22652 3680 22704 3732
rect 24676 3680 24728 3732
rect 25136 3723 25188 3732
rect 25136 3689 25145 3723
rect 25145 3689 25179 3723
rect 25179 3689 25188 3723
rect 25136 3680 25188 3689
rect 25228 3723 25280 3732
rect 25228 3689 25237 3723
rect 25237 3689 25271 3723
rect 25271 3689 25280 3723
rect 25228 3680 25280 3689
rect 26884 3612 26936 3664
rect 29000 3680 29052 3732
rect 22836 3544 22888 3596
rect 22376 3408 22428 3460
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 22836 3383 22888 3392
rect 22836 3349 22845 3383
rect 22845 3349 22879 3383
rect 22879 3349 22888 3383
rect 22836 3340 22888 3349
rect 24584 3476 24636 3528
rect 26148 3587 26200 3596
rect 26148 3553 26157 3587
rect 26157 3553 26191 3587
rect 26191 3553 26200 3587
rect 26148 3544 26200 3553
rect 27988 3655 28040 3664
rect 27988 3621 27997 3655
rect 27997 3621 28031 3655
rect 28031 3621 28040 3655
rect 27988 3612 28040 3621
rect 30380 3612 30432 3664
rect 26516 3476 26568 3528
rect 28080 3476 28132 3528
rect 24952 3451 25004 3460
rect 24952 3417 24961 3451
rect 24961 3417 24995 3451
rect 24995 3417 25004 3451
rect 24952 3408 25004 3417
rect 26608 3383 26660 3392
rect 26608 3349 26617 3383
rect 26617 3349 26651 3383
rect 26651 3349 26660 3383
rect 26608 3340 26660 3349
rect 27252 3408 27304 3460
rect 28356 3383 28408 3392
rect 28356 3349 28365 3383
rect 28365 3349 28399 3383
rect 28399 3349 28408 3383
rect 28356 3340 28408 3349
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 11436 3238 11488 3290
rect 11500 3238 11552 3290
rect 11564 3238 11616 3290
rect 11628 3238 11680 3290
rect 11692 3238 11744 3290
rect 19210 3238 19262 3290
rect 19274 3238 19326 3290
rect 19338 3238 19390 3290
rect 19402 3238 19454 3290
rect 19466 3238 19518 3290
rect 26984 3238 27036 3290
rect 27048 3238 27100 3290
rect 27112 3238 27164 3290
rect 27176 3238 27228 3290
rect 27240 3238 27292 3290
rect 4160 3136 4212 3188
rect 5540 3136 5592 3188
rect 6368 3136 6420 3188
rect 9312 3179 9364 3188
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 2228 2932 2280 2984
rect 4988 3068 5040 3120
rect 6184 3068 6236 3120
rect 9220 3111 9272 3120
rect 9220 3077 9229 3111
rect 9229 3077 9263 3111
rect 9263 3077 9272 3111
rect 9220 3068 9272 3077
rect 2044 2864 2096 2916
rect 3424 2864 3476 2916
rect 4712 3000 4764 3052
rect 5448 3000 5500 3052
rect 4896 2932 4948 2984
rect 3516 2796 3568 2848
rect 5172 2796 5224 2848
rect 6092 2864 6144 2916
rect 6460 2975 6512 2984
rect 6460 2941 6469 2975
rect 6469 2941 6503 2975
rect 6503 2941 6512 2975
rect 6460 2932 6512 2941
rect 6736 2975 6788 2984
rect 6736 2941 6745 2975
rect 6745 2941 6779 2975
rect 6779 2941 6788 2975
rect 6736 2932 6788 2941
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 7012 2864 7064 2916
rect 8116 3000 8168 3052
rect 9036 3000 9088 3052
rect 10416 3136 10468 3188
rect 19064 3136 19116 3188
rect 22100 3136 22152 3188
rect 22284 3179 22336 3188
rect 22284 3145 22293 3179
rect 22293 3145 22327 3179
rect 22327 3145 22336 3179
rect 22284 3136 22336 3145
rect 26516 3179 26568 3188
rect 26516 3145 26525 3179
rect 26525 3145 26559 3179
rect 26559 3145 26568 3179
rect 26516 3136 26568 3145
rect 27068 3136 27120 3188
rect 28356 3179 28408 3188
rect 28356 3145 28365 3179
rect 28365 3145 28399 3179
rect 28399 3145 28408 3179
rect 28356 3136 28408 3145
rect 30380 3179 30432 3188
rect 30380 3145 30389 3179
rect 30389 3145 30423 3179
rect 30423 3145 30432 3179
rect 30380 3136 30432 3145
rect 10508 3111 10560 3120
rect 10508 3077 10517 3111
rect 10517 3077 10551 3111
rect 10551 3077 10560 3111
rect 10508 3068 10560 3077
rect 11796 3068 11848 3120
rect 14096 3068 14148 3120
rect 26700 3111 26752 3120
rect 26700 3077 26709 3111
rect 26709 3077 26743 3111
rect 26743 3077 26752 3111
rect 26700 3068 26752 3077
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9588 3000 9640 3052
rect 12532 3000 12584 3052
rect 13176 3000 13228 3052
rect 10140 2975 10192 2984
rect 10140 2941 10158 2975
rect 10158 2941 10192 2975
rect 10140 2932 10192 2941
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 8484 2907 8536 2916
rect 8484 2873 8493 2907
rect 8493 2873 8527 2907
rect 8527 2873 8536 2907
rect 8484 2864 8536 2873
rect 6000 2839 6052 2848
rect 6000 2805 6027 2839
rect 6027 2805 6052 2839
rect 6000 2796 6052 2805
rect 7104 2796 7156 2848
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 10048 2796 10100 2848
rect 10324 2796 10376 2848
rect 11244 2932 11296 2984
rect 11336 2932 11388 2984
rect 12624 2932 12676 2984
rect 15016 3000 15068 3052
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 18604 2932 18656 2984
rect 20352 2932 20404 2984
rect 20720 3000 20772 3052
rect 24400 3000 24452 3052
rect 23664 2975 23716 2984
rect 23664 2941 23673 2975
rect 23673 2941 23707 2975
rect 23707 2941 23716 2975
rect 23664 2932 23716 2941
rect 13728 2864 13780 2916
rect 14832 2864 14884 2916
rect 21272 2864 21324 2916
rect 11336 2796 11388 2848
rect 12440 2796 12492 2848
rect 12992 2796 13044 2848
rect 16948 2796 17000 2848
rect 23296 2864 23348 2916
rect 26148 2864 26200 2916
rect 26608 2932 26660 2984
rect 27436 3000 27488 3052
rect 27068 2975 27120 2984
rect 27068 2941 27077 2975
rect 27077 2941 27111 2975
rect 27111 2941 27120 2975
rect 27068 2932 27120 2941
rect 28080 2932 28132 2984
rect 24032 2839 24084 2848
rect 24032 2805 24041 2839
rect 24041 2805 24075 2839
rect 24075 2805 24084 2839
rect 24032 2796 24084 2805
rect 24124 2796 24176 2848
rect 25136 2796 25188 2848
rect 26792 2907 26844 2916
rect 26792 2873 26801 2907
rect 26801 2873 26835 2907
rect 26835 2873 26844 2907
rect 26792 2864 26844 2873
rect 28264 2864 28316 2916
rect 28448 2864 28500 2916
rect 27988 2796 28040 2848
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 12096 2694 12148 2746
rect 12160 2694 12212 2746
rect 12224 2694 12276 2746
rect 12288 2694 12340 2746
rect 12352 2694 12404 2746
rect 19870 2694 19922 2746
rect 19934 2694 19986 2746
rect 19998 2694 20050 2746
rect 20062 2694 20114 2746
rect 20126 2694 20178 2746
rect 27644 2694 27696 2746
rect 27708 2694 27760 2746
rect 27772 2694 27824 2746
rect 27836 2694 27888 2746
rect 27900 2694 27952 2746
rect 2964 2592 3016 2644
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 3516 2499 3568 2508
rect 3516 2465 3525 2499
rect 3525 2465 3559 2499
rect 3559 2465 3568 2499
rect 3516 2456 3568 2465
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 6460 2592 6512 2644
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 9588 2592 9640 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 10968 2635 11020 2644
rect 10968 2601 10977 2635
rect 10977 2601 11011 2635
rect 11011 2601 11020 2635
rect 10968 2592 11020 2601
rect 6000 2456 6052 2508
rect 6736 2524 6788 2576
rect 9864 2524 9916 2576
rect 10232 2524 10284 2576
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 11244 2499 11296 2508
rect 4068 2388 4120 2440
rect 5816 2388 5868 2440
rect 6092 2320 6144 2372
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 6828 2320 6880 2372
rect 8300 2431 8352 2440
rect 8300 2397 8334 2431
rect 8334 2397 8352 2431
rect 8300 2388 8352 2397
rect 9128 2388 9180 2440
rect 9496 2388 9548 2440
rect 4712 2252 4764 2304
rect 8944 2252 8996 2304
rect 9404 2295 9456 2304
rect 9404 2261 9413 2295
rect 9413 2261 9447 2295
rect 9447 2261 9456 2295
rect 9404 2252 9456 2261
rect 11244 2465 11253 2499
rect 11253 2465 11287 2499
rect 11287 2465 11296 2499
rect 11244 2456 11296 2465
rect 11336 2499 11388 2508
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 12440 2567 12492 2576
rect 12440 2533 12449 2567
rect 12449 2533 12483 2567
rect 12483 2533 12492 2567
rect 12440 2524 12492 2533
rect 13728 2592 13780 2644
rect 15016 2592 15068 2644
rect 12808 2456 12860 2508
rect 12992 2456 13044 2508
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 17224 2592 17276 2644
rect 18880 2592 18932 2644
rect 19708 2592 19760 2644
rect 21272 2635 21324 2644
rect 21272 2601 21281 2635
rect 21281 2601 21315 2635
rect 21315 2601 21324 2635
rect 21272 2592 21324 2601
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 10140 2320 10192 2372
rect 11888 2388 11940 2440
rect 17040 2456 17092 2508
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 18788 2524 18840 2576
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 18972 2456 19024 2508
rect 20904 2499 20956 2508
rect 20904 2465 20913 2499
rect 20913 2465 20947 2499
rect 20947 2465 20956 2499
rect 20904 2456 20956 2465
rect 21640 2499 21692 2508
rect 21640 2465 21649 2499
rect 21649 2465 21683 2499
rect 21683 2465 21692 2499
rect 21640 2456 21692 2465
rect 18328 2388 18380 2440
rect 20352 2388 20404 2440
rect 10232 2252 10284 2304
rect 11796 2252 11848 2304
rect 14096 2320 14148 2372
rect 17132 2320 17184 2372
rect 18604 2363 18656 2372
rect 18604 2329 18613 2363
rect 18613 2329 18647 2363
rect 18647 2329 18656 2363
rect 18604 2320 18656 2329
rect 22192 2456 22244 2508
rect 22652 2456 22704 2508
rect 23756 2456 23808 2508
rect 23940 2499 23992 2508
rect 23940 2465 23949 2499
rect 23949 2465 23983 2499
rect 23983 2465 23992 2499
rect 23940 2456 23992 2465
rect 24124 2499 24176 2508
rect 24124 2465 24133 2499
rect 24133 2465 24167 2499
rect 24167 2465 24176 2499
rect 24124 2456 24176 2465
rect 23112 2388 23164 2440
rect 24492 2524 24544 2576
rect 26700 2592 26752 2644
rect 26884 2592 26936 2644
rect 28264 2592 28316 2644
rect 24400 2499 24452 2508
rect 24400 2465 24409 2499
rect 24409 2465 24443 2499
rect 24443 2465 24452 2499
rect 24400 2456 24452 2465
rect 26516 2524 26568 2576
rect 27436 2524 27488 2576
rect 24676 2499 24728 2508
rect 24676 2465 24685 2499
rect 24685 2465 24719 2499
rect 24719 2465 24728 2499
rect 24676 2456 24728 2465
rect 24860 2499 24912 2508
rect 24860 2465 24869 2499
rect 24869 2465 24903 2499
rect 24903 2465 24912 2499
rect 24860 2456 24912 2465
rect 24584 2388 24636 2440
rect 25320 2456 25372 2508
rect 25780 2456 25832 2508
rect 27068 2456 27120 2508
rect 27620 2499 27672 2508
rect 27620 2465 27629 2499
rect 27629 2465 27663 2499
rect 27663 2465 27672 2499
rect 27620 2456 27672 2465
rect 28080 2388 28132 2440
rect 13636 2252 13688 2304
rect 15292 2252 15344 2304
rect 15752 2252 15804 2304
rect 16304 2295 16356 2304
rect 16304 2261 16313 2295
rect 16313 2261 16347 2295
rect 16347 2261 16356 2295
rect 16304 2252 16356 2261
rect 16488 2295 16540 2304
rect 16488 2261 16497 2295
rect 16497 2261 16531 2295
rect 16531 2261 16540 2295
rect 16488 2252 16540 2261
rect 17868 2295 17920 2304
rect 17868 2261 17877 2295
rect 17877 2261 17911 2295
rect 17911 2261 17920 2295
rect 17868 2252 17920 2261
rect 19064 2252 19116 2304
rect 20076 2252 20128 2304
rect 23296 2363 23348 2372
rect 23296 2329 23305 2363
rect 23305 2329 23339 2363
rect 23339 2329 23348 2363
rect 23296 2320 23348 2329
rect 23664 2320 23716 2372
rect 23020 2252 23072 2304
rect 25136 2320 25188 2372
rect 26240 2320 26292 2372
rect 26700 2320 26752 2372
rect 25228 2252 25280 2304
rect 25688 2295 25740 2304
rect 25688 2261 25697 2295
rect 25697 2261 25731 2295
rect 25731 2261 25740 2295
rect 25688 2252 25740 2261
rect 26424 2252 26476 2304
rect 27988 2320 28040 2372
rect 27344 2295 27396 2304
rect 27344 2261 27353 2295
rect 27353 2261 27387 2295
rect 27387 2261 27396 2295
rect 27344 2252 27396 2261
rect 27436 2295 27488 2304
rect 27436 2261 27445 2295
rect 27445 2261 27479 2295
rect 27479 2261 27488 2295
rect 27436 2252 27488 2261
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 11436 2150 11488 2202
rect 11500 2150 11552 2202
rect 11564 2150 11616 2202
rect 11628 2150 11680 2202
rect 11692 2150 11744 2202
rect 19210 2150 19262 2202
rect 19274 2150 19326 2202
rect 19338 2150 19390 2202
rect 19402 2150 19454 2202
rect 19466 2150 19518 2202
rect 26984 2150 27036 2202
rect 27048 2150 27100 2202
rect 27112 2150 27164 2202
rect 27176 2150 27228 2202
rect 27240 2150 27292 2202
rect 6368 2048 6420 2100
rect 7288 2048 7340 2100
rect 8024 2048 8076 2100
rect 10232 2048 10284 2100
rect 10416 2048 10468 2100
rect 11888 2048 11940 2100
rect 12348 2048 12400 2100
rect 6828 1912 6880 1964
rect 8300 1912 8352 1964
rect 5172 1887 5224 1896
rect 5172 1853 5206 1887
rect 5206 1853 5224 1887
rect 5172 1844 5224 1853
rect 9772 1887 9824 1896
rect 9772 1853 9781 1887
rect 9781 1853 9815 1887
rect 9815 1853 9824 1887
rect 9772 1844 9824 1853
rect 11060 1887 11112 1896
rect 11796 1912 11848 1964
rect 12532 1912 12584 1964
rect 12900 2048 12952 2100
rect 13636 2048 13688 2100
rect 15568 2048 15620 2100
rect 18604 2048 18656 2100
rect 11060 1853 11078 1887
rect 11078 1853 11112 1887
rect 11060 1844 11112 1853
rect 5080 1776 5132 1828
rect 6092 1776 6144 1828
rect 8852 1776 8904 1828
rect 10600 1776 10652 1828
rect 4252 1708 4304 1760
rect 7104 1708 7156 1760
rect 9404 1708 9456 1760
rect 12348 1887 12400 1896
rect 12348 1853 12357 1887
rect 12357 1853 12391 1887
rect 12391 1853 12400 1887
rect 12348 1844 12400 1853
rect 13636 1844 13688 1896
rect 13728 1887 13780 1896
rect 13728 1853 13737 1887
rect 13737 1853 13771 1887
rect 13771 1853 13780 1887
rect 13728 1844 13780 1853
rect 14004 1887 14056 1896
rect 14004 1853 14013 1887
rect 14013 1853 14047 1887
rect 14047 1853 14056 1887
rect 14004 1844 14056 1853
rect 14832 1955 14884 1964
rect 14832 1921 14841 1955
rect 14841 1921 14875 1955
rect 14875 1921 14884 1955
rect 14832 1912 14884 1921
rect 15292 1955 15344 1964
rect 15292 1921 15301 1955
rect 15301 1921 15335 1955
rect 15335 1921 15344 1955
rect 15292 1912 15344 1921
rect 16580 1912 16632 1964
rect 17040 1912 17092 1964
rect 17132 1955 17184 1964
rect 17132 1921 17141 1955
rect 17141 1921 17175 1955
rect 17175 1921 17184 1955
rect 17132 1912 17184 1921
rect 11980 1708 12032 1760
rect 13360 1751 13412 1760
rect 13360 1717 13369 1751
rect 13369 1717 13403 1751
rect 13403 1717 13412 1751
rect 13360 1708 13412 1717
rect 13728 1708 13780 1760
rect 16948 1887 17000 1896
rect 16948 1853 16957 1887
rect 16957 1853 16991 1887
rect 16991 1853 17000 1887
rect 16948 1844 17000 1853
rect 19156 1844 19208 1896
rect 20076 1980 20128 2032
rect 20444 1980 20496 2032
rect 19708 1887 19760 1896
rect 19708 1853 19717 1887
rect 19717 1853 19751 1887
rect 19751 1853 19760 1887
rect 19708 1844 19760 1853
rect 15568 1819 15620 1828
rect 15568 1785 15602 1819
rect 15602 1785 15620 1819
rect 15568 1776 15620 1785
rect 17684 1776 17736 1828
rect 17960 1776 18012 1828
rect 18788 1776 18840 1828
rect 20076 1887 20128 1896
rect 20076 1853 20085 1887
rect 20085 1853 20119 1887
rect 20119 1853 20128 1887
rect 20076 1844 20128 1853
rect 20352 1887 20404 1896
rect 20352 1853 20361 1887
rect 20361 1853 20395 1887
rect 20395 1853 20404 1887
rect 20352 1844 20404 1853
rect 20444 1887 20496 1896
rect 20444 1853 20453 1887
rect 20453 1853 20487 1887
rect 20487 1853 20496 1887
rect 20444 1844 20496 1853
rect 24216 2048 24268 2100
rect 22836 1887 22888 1896
rect 22836 1853 22845 1887
rect 22845 1853 22879 1887
rect 22879 1853 22888 1887
rect 22836 1844 22888 1853
rect 24032 1980 24084 2032
rect 24492 2048 24544 2100
rect 25688 2091 25740 2100
rect 25688 2057 25697 2091
rect 25697 2057 25731 2091
rect 25731 2057 25740 2091
rect 25688 2048 25740 2057
rect 26148 2091 26200 2100
rect 26148 2057 26157 2091
rect 26157 2057 26191 2091
rect 26191 2057 26200 2091
rect 26148 2048 26200 2057
rect 23756 1912 23808 1964
rect 27620 2048 27672 2100
rect 28908 1980 28960 2032
rect 25228 1955 25280 1964
rect 25228 1921 25237 1955
rect 25237 1921 25271 1955
rect 25271 1921 25280 1955
rect 25228 1912 25280 1921
rect 26424 1955 26476 1964
rect 26424 1921 26433 1955
rect 26433 1921 26467 1955
rect 26467 1921 26476 1955
rect 26424 1912 26476 1921
rect 23112 1887 23164 1896
rect 23112 1853 23121 1887
rect 23121 1853 23155 1887
rect 23155 1853 23164 1887
rect 23112 1844 23164 1853
rect 23204 1887 23256 1896
rect 23204 1853 23213 1887
rect 23213 1853 23247 1887
rect 23247 1853 23256 1887
rect 23204 1844 23256 1853
rect 22376 1776 22428 1828
rect 24676 1844 24728 1896
rect 25136 1844 25188 1896
rect 26516 1844 26568 1896
rect 28080 1887 28132 1896
rect 28080 1853 28089 1887
rect 28089 1853 28123 1887
rect 28123 1853 28132 1887
rect 28080 1844 28132 1853
rect 15476 1708 15528 1760
rect 19432 1751 19484 1760
rect 19432 1717 19441 1751
rect 19441 1717 19475 1751
rect 19475 1717 19484 1751
rect 19432 1708 19484 1717
rect 19616 1708 19668 1760
rect 20628 1708 20680 1760
rect 22652 1751 22704 1760
rect 22652 1717 22661 1751
rect 22661 1717 22695 1751
rect 22695 1717 22704 1751
rect 22652 1708 22704 1717
rect 25780 1776 25832 1828
rect 26976 1776 27028 1828
rect 23204 1708 23256 1760
rect 24860 1708 24912 1760
rect 25872 1751 25924 1760
rect 25872 1717 25881 1751
rect 25881 1717 25915 1751
rect 25915 1717 25924 1751
rect 25872 1708 25924 1717
rect 26424 1708 26476 1760
rect 26792 1708 26844 1760
rect 27988 1751 28040 1760
rect 27988 1717 27997 1751
rect 27997 1717 28031 1751
rect 28031 1717 28040 1751
rect 27988 1708 28040 1717
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 12096 1606 12148 1658
rect 12160 1606 12212 1658
rect 12224 1606 12276 1658
rect 12288 1606 12340 1658
rect 12352 1606 12404 1658
rect 19870 1606 19922 1658
rect 19934 1606 19986 1658
rect 19998 1606 20050 1658
rect 20062 1606 20114 1658
rect 20126 1606 20178 1658
rect 27644 1606 27696 1658
rect 27708 1606 27760 1658
rect 27772 1606 27824 1658
rect 27836 1606 27888 1658
rect 27900 1606 27952 1658
rect 6828 1504 6880 1556
rect 8300 1504 8352 1556
rect 8852 1547 8904 1556
rect 8852 1513 8861 1547
rect 8861 1513 8895 1547
rect 8895 1513 8904 1547
rect 8852 1504 8904 1513
rect 4712 1436 4764 1488
rect 7012 1436 7064 1488
rect 8024 1479 8076 1488
rect 8024 1445 8033 1479
rect 8033 1445 8067 1479
rect 8067 1445 8076 1479
rect 8024 1436 8076 1445
rect 8668 1479 8720 1488
rect 8668 1445 8677 1479
rect 8677 1445 8711 1479
rect 8711 1445 8720 1479
rect 8668 1436 8720 1445
rect 4252 1411 4304 1420
rect 4252 1377 4261 1411
rect 4261 1377 4295 1411
rect 4295 1377 4304 1411
rect 4252 1368 4304 1377
rect 6092 1411 6144 1420
rect 6092 1377 6101 1411
rect 6101 1377 6135 1411
rect 6135 1377 6144 1411
rect 6092 1368 6144 1377
rect 8392 1368 8444 1420
rect 8852 1368 8904 1420
rect 5816 1343 5868 1352
rect 5816 1309 5825 1343
rect 5825 1309 5859 1343
rect 5859 1309 5868 1343
rect 5816 1300 5868 1309
rect 6184 1343 6236 1352
rect 6184 1309 6193 1343
rect 6193 1309 6227 1343
rect 6227 1309 6236 1343
rect 6184 1300 6236 1309
rect 7196 1300 7248 1352
rect 5448 1232 5500 1284
rect 7472 1232 7524 1284
rect 10600 1504 10652 1556
rect 9220 1436 9272 1488
rect 12624 1436 12676 1488
rect 13360 1436 13412 1488
rect 14004 1547 14056 1556
rect 14004 1513 14013 1547
rect 14013 1513 14047 1547
rect 14047 1513 14056 1547
rect 14004 1504 14056 1513
rect 15476 1547 15528 1556
rect 15476 1513 15485 1547
rect 15485 1513 15519 1547
rect 15519 1513 15528 1547
rect 15476 1504 15528 1513
rect 15568 1547 15620 1556
rect 15568 1513 15577 1547
rect 15577 1513 15611 1547
rect 15611 1513 15620 1547
rect 15568 1504 15620 1513
rect 17224 1504 17276 1556
rect 17684 1547 17736 1556
rect 17684 1513 17693 1547
rect 17693 1513 17727 1547
rect 17727 1513 17736 1547
rect 17684 1504 17736 1513
rect 19064 1504 19116 1556
rect 19708 1504 19760 1556
rect 20628 1504 20680 1556
rect 23020 1547 23072 1556
rect 23020 1513 23029 1547
rect 23029 1513 23063 1547
rect 23063 1513 23072 1547
rect 23020 1504 23072 1513
rect 16488 1479 16540 1488
rect 16488 1445 16522 1479
rect 16522 1445 16540 1479
rect 16488 1436 16540 1445
rect 17868 1436 17920 1488
rect 9036 1411 9088 1420
rect 9036 1377 9045 1411
rect 9045 1377 9079 1411
rect 9079 1377 9088 1411
rect 9036 1368 9088 1377
rect 11980 1368 12032 1420
rect 13728 1368 13780 1420
rect 14096 1411 14148 1420
rect 14096 1377 14105 1411
rect 14105 1377 14139 1411
rect 14139 1377 14148 1411
rect 14096 1368 14148 1377
rect 15752 1411 15804 1420
rect 15752 1377 15761 1411
rect 15761 1377 15795 1411
rect 15795 1377 15804 1411
rect 15752 1368 15804 1377
rect 16304 1368 16356 1420
rect 17960 1411 18012 1420
rect 17960 1377 17969 1411
rect 17969 1377 18003 1411
rect 18003 1377 18012 1411
rect 17960 1368 18012 1377
rect 19432 1436 19484 1488
rect 24124 1504 24176 1556
rect 25780 1504 25832 1556
rect 25872 1436 25924 1488
rect 19156 1368 19208 1420
rect 19616 1411 19668 1420
rect 19616 1377 19625 1411
rect 19625 1377 19659 1411
rect 19659 1377 19668 1411
rect 19616 1368 19668 1377
rect 22652 1368 22704 1420
rect 24032 1368 24084 1420
rect 26884 1504 26936 1556
rect 26976 1547 27028 1556
rect 26976 1513 26985 1547
rect 26985 1513 27019 1547
rect 27019 1513 27028 1547
rect 26976 1504 27028 1513
rect 27344 1504 27396 1556
rect 27988 1436 28040 1488
rect 11796 1232 11848 1284
rect 6000 1207 6052 1216
rect 6000 1173 6009 1207
rect 6009 1173 6043 1207
rect 6043 1173 6052 1207
rect 6000 1164 6052 1173
rect 8576 1164 8628 1216
rect 18696 1300 18748 1352
rect 26240 1343 26292 1352
rect 26240 1309 26249 1343
rect 26249 1309 26283 1343
rect 26283 1309 26292 1343
rect 26240 1300 26292 1309
rect 26424 1343 26476 1352
rect 26424 1309 26433 1343
rect 26433 1309 26467 1343
rect 26467 1309 26476 1343
rect 26424 1300 26476 1309
rect 28908 1547 28960 1556
rect 28908 1513 28917 1547
rect 28917 1513 28951 1547
rect 28951 1513 28960 1547
rect 28908 1504 28960 1513
rect 23112 1232 23164 1284
rect 16580 1164 16632 1216
rect 19156 1207 19208 1216
rect 19156 1173 19165 1207
rect 19165 1173 19199 1207
rect 19199 1173 19208 1207
rect 19156 1164 19208 1173
rect 19616 1164 19668 1216
rect 23940 1164 23992 1216
rect 27436 1164 27488 1216
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 11436 1062 11488 1114
rect 11500 1062 11552 1114
rect 11564 1062 11616 1114
rect 11628 1062 11680 1114
rect 11692 1062 11744 1114
rect 19210 1062 19262 1114
rect 19274 1062 19326 1114
rect 19338 1062 19390 1114
rect 19402 1062 19454 1114
rect 19466 1062 19518 1114
rect 26984 1062 27036 1114
rect 27048 1062 27100 1114
rect 27112 1062 27164 1114
rect 27176 1062 27228 1114
rect 27240 1062 27292 1114
rect 6920 1003 6972 1012
rect 6920 969 6929 1003
rect 6929 969 6963 1003
rect 6963 969 6972 1003
rect 6920 960 6972 969
rect 7196 1003 7248 1012
rect 7196 969 7205 1003
rect 7205 969 7239 1003
rect 7239 969 7248 1003
rect 7196 960 7248 969
rect 8024 960 8076 1012
rect 8668 960 8720 1012
rect 9772 960 9824 1012
rect 18696 1003 18748 1012
rect 18696 969 18705 1003
rect 18705 969 18739 1003
rect 18739 969 18748 1003
rect 18696 960 18748 969
rect 18880 1003 18932 1012
rect 18880 969 18889 1003
rect 18889 969 18923 1003
rect 18923 969 18932 1003
rect 18880 960 18932 969
rect 5816 824 5868 876
rect 8576 824 8628 876
rect 7104 799 7156 808
rect 7104 765 7113 799
rect 7113 765 7147 799
rect 7147 765 7156 799
rect 7104 756 7156 765
rect 8392 799 8444 808
rect 8392 765 8401 799
rect 8401 765 8435 799
rect 8435 765 8444 799
rect 8392 756 8444 765
rect 9036 756 9088 808
rect 18328 799 18380 808
rect 18328 765 18337 799
rect 18337 765 18371 799
rect 18371 765 18380 799
rect 18328 756 18380 765
rect 19616 799 19668 808
rect 19616 765 19650 799
rect 19650 765 19668 799
rect 19616 756 19668 765
rect 7472 688 7524 740
rect 18880 731 18932 740
rect 18880 697 18907 731
rect 18907 697 18932 731
rect 18880 688 18932 697
rect 18972 688 19024 740
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 12096 518 12148 570
rect 12160 518 12212 570
rect 12224 518 12276 570
rect 12288 518 12340 570
rect 12352 518 12404 570
rect 19870 518 19922 570
rect 19934 518 19986 570
rect 19998 518 20050 570
rect 20062 518 20114 570
rect 20126 518 20178 570
rect 27644 518 27696 570
rect 27708 518 27760 570
rect 27772 518 27824 570
rect 27836 518 27888 570
rect 27900 518 27952 570
<< metal2 >>
rect 11794 21992 11850 22001
rect 11794 21927 11850 21936
rect 12254 21992 12310 22001
rect 12254 21927 12310 21936
rect 24398 21992 24454 22001
rect 24398 21927 24454 21936
rect 27342 21992 27398 22001
rect 27342 21927 27398 21936
rect 27710 21992 27766 22001
rect 27710 21927 27766 21936
rect 8666 21856 8722 21865
rect 3662 21788 3970 21797
rect 8666 21791 8722 21800
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 6090 21720 6146 21729
rect 6090 21655 6092 21664
rect 6144 21655 6146 21664
rect 8022 21720 8078 21729
rect 8022 21655 8024 21664
rect 6092 21626 6144 21632
rect 8076 21655 8078 21664
rect 8390 21720 8446 21729
rect 8680 21690 8708 21791
rect 11436 21788 11744 21797
rect 11436 21786 11442 21788
rect 11498 21786 11522 21788
rect 11578 21786 11602 21788
rect 11658 21786 11682 21788
rect 11738 21786 11744 21788
rect 11498 21734 11500 21786
rect 11680 21734 11682 21786
rect 11436 21732 11442 21734
rect 11498 21732 11522 21734
rect 11578 21732 11602 21734
rect 11658 21732 11682 21734
rect 11738 21732 11744 21734
rect 11436 21723 11744 21732
rect 11808 21690 11836 21927
rect 12268 21690 12296 21927
rect 22190 21856 22246 21865
rect 19210 21788 19518 21797
rect 22190 21791 22246 21800
rect 23846 21856 23902 21865
rect 23846 21791 23902 21800
rect 19210 21786 19216 21788
rect 19272 21786 19296 21788
rect 19352 21786 19376 21788
rect 19432 21786 19456 21788
rect 19512 21786 19518 21788
rect 19272 21734 19274 21786
rect 19454 21734 19456 21786
rect 19210 21732 19216 21734
rect 19272 21732 19296 21734
rect 19352 21732 19376 21734
rect 19432 21732 19456 21734
rect 19512 21732 19518 21734
rect 12990 21720 13046 21729
rect 19210 21723 19518 21732
rect 8390 21655 8392 21664
rect 8024 21626 8076 21632
rect 8444 21655 8446 21664
rect 8668 21684 8720 21690
rect 8392 21626 8444 21632
rect 8668 21626 8720 21632
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 12256 21684 12308 21690
rect 12990 21655 12992 21664
rect 12256 21626 12308 21632
rect 13044 21655 13046 21664
rect 18788 21684 18840 21690
rect 12992 21626 13044 21632
rect 18788 21626 18840 21632
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 1412 20602 1440 21422
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 1964 21010 1992 21286
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 2504 21004 2556 21010
rect 2504 20946 2556 20952
rect 1400 20596 1452 20602
rect 1400 20538 1452 20544
rect 1308 20392 1360 20398
rect 1412 20346 1440 20538
rect 1360 20340 1440 20346
rect 1308 20334 1440 20340
rect 1320 20318 1440 20334
rect 1412 19310 1440 20318
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2332 20058 2360 20266
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2056 19446 2084 19858
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 2148 19310 2176 19654
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 1412 17066 1440 19246
rect 2516 19242 2544 20946
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2792 20058 2820 20198
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2884 19990 2912 21286
rect 2976 21146 3004 21422
rect 3148 21412 3200 21418
rect 3148 21354 3200 21360
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 2976 19310 3004 21082
rect 3056 20324 3108 20330
rect 3056 20266 3108 20272
rect 3068 20058 3096 20266
rect 3160 20058 3188 21354
rect 4172 21010 4200 21422
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 5276 21010 5304 21286
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 3240 20868 3292 20874
rect 3240 20810 3292 20816
rect 3252 20466 3280 20810
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 3160 19854 3188 19994
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3160 19718 3188 19790
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1596 18834 1624 19110
rect 3160 18986 3188 19654
rect 3252 19514 3280 19654
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3344 19378 3372 20742
rect 3528 20244 3556 20946
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3608 20256 3660 20262
rect 3528 20216 3608 20244
rect 3608 20198 3660 20204
rect 3896 19922 3924 20334
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3988 19922 4016 20198
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3528 19718 3556 19858
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 2976 18958 3188 18986
rect 3252 18970 3280 19246
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3240 18964 3292 18970
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2792 17746 2820 18090
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2424 17134 2452 17478
rect 2700 17202 2728 17682
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 1400 17060 1452 17066
rect 1400 17002 1452 17008
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 1412 16046 1440 17002
rect 2700 16658 2728 17002
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2792 16522 2820 17682
rect 2976 16658 3004 18958
rect 3240 18906 3292 18912
rect 3148 18896 3200 18902
rect 3148 18838 3200 18844
rect 3056 17740 3108 17746
rect 3160 17728 3188 18838
rect 3252 18222 3280 18906
rect 3344 18834 3372 19110
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3436 18154 3464 18770
rect 3528 18222 3556 19654
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 4080 19514 4108 20946
rect 4172 20602 4200 20946
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4172 19394 4200 19654
rect 4724 19446 4752 20946
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4816 19990 4844 20742
rect 4908 20602 4936 20946
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 5368 19922 5396 21422
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6656 21078 6684 21286
rect 6840 21146 6868 21286
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6932 21010 6960 21422
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6932 20602 6960 20946
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 5448 20392 5500 20398
rect 6920 20392 6972 20398
rect 5448 20334 5500 20340
rect 6734 20360 6790 20369
rect 5460 20058 5488 20334
rect 5908 20324 5960 20330
rect 6920 20334 6972 20340
rect 6734 20295 6736 20304
rect 5908 20266 5960 20272
rect 6788 20295 6790 20304
rect 6736 20266 6788 20272
rect 5920 20058 5948 20266
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 6104 19922 6132 20198
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 4080 19378 4200 19394
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4068 19372 4200 19378
rect 4120 19366 4200 19372
rect 4068 19314 4120 19320
rect 4080 19242 4108 19314
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 4080 18290 4108 18770
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3108 17700 3188 17728
rect 3056 17682 3108 17688
rect 3252 17610 3280 18022
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3240 17604 3292 17610
rect 3240 17546 3292 17552
rect 3252 16794 3280 17546
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16046 1992 16390
rect 2688 16176 2740 16182
rect 2688 16118 2740 16124
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1412 15638 1440 15982
rect 2700 15706 2728 16118
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 1400 15632 1452 15638
rect 1400 15574 1452 15580
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 14958 1348 15506
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1412 15026 1440 15302
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 1320 13870 1348 14894
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14482 1532 14758
rect 1596 14550 1624 15302
rect 1584 14544 1636 14550
rect 1584 14486 1636 14492
rect 2792 14482 2820 16458
rect 2976 14550 3004 16594
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 3068 14346 3096 15438
rect 3344 15026 3372 16934
rect 3436 16658 3464 17818
rect 3528 17338 3556 18158
rect 3896 17882 3924 18158
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3896 17746 3924 17818
rect 4080 17746 4108 18226
rect 4172 17814 4200 18566
rect 4264 18154 4292 18634
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4264 17864 4292 18090
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 4264 17836 4384 17864
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 3884 17740 3936 17746
rect 3884 17682 3936 17688
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4160 17672 4212 17678
rect 4158 17640 4160 17649
rect 4212 17640 4214 17649
rect 4068 17604 4120 17610
rect 4158 17575 4214 17584
rect 4068 17546 4120 17552
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 4080 17338 4108 17546
rect 4356 17542 4384 17836
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 4160 17536 4212 17542
rect 4344 17536 4396 17542
rect 4212 17496 4292 17524
rect 4160 17478 4212 17484
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3896 16998 3924 17206
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3896 16590 3924 16934
rect 4172 16794 4200 17070
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4080 16674 4108 16730
rect 4080 16658 4200 16674
rect 4264 16658 4292 17496
rect 4344 17478 4396 17484
rect 4356 16998 4384 17478
rect 4540 17134 4568 17682
rect 4724 17649 4752 18702
rect 4816 18630 4844 19110
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4816 18222 4844 18566
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4710 17640 4766 17649
rect 4710 17575 4766 17584
rect 4816 17134 4844 18022
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4724 16726 4752 17002
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4080 16652 4212 16658
rect 4080 16646 4160 16652
rect 4160 16594 4212 16600
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 4172 16046 4200 16594
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4264 16114 4292 16390
rect 4724 16182 4752 16662
rect 4908 16658 4936 19858
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 19378 5120 19654
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5000 18426 5028 18702
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4988 18216 5040 18222
rect 4988 18158 5040 18164
rect 5000 17814 5028 18158
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 4986 17640 5042 17649
rect 4986 17575 5042 17584
rect 5000 17134 5028 17575
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4816 16538 4844 16594
rect 4816 16510 4936 16538
rect 4908 16250 4936 16510
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3424 14544 3476 14550
rect 3424 14486 3476 14492
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 3068 14006 3096 14282
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 1308 13864 1360 13870
rect 2872 13864 2924 13870
rect 1360 13812 1440 13818
rect 1308 13806 1440 13812
rect 2872 13806 2924 13812
rect 1320 13790 1440 13806
rect 1412 12782 1440 13790
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13394 2360 13670
rect 2884 13530 2912 13806
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2976 13462 3004 13670
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 3436 13394 3464 14486
rect 3528 14414 3556 14894
rect 3988 14550 4016 14894
rect 4080 14550 4108 15438
rect 4816 15026 4844 15846
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4620 14952 4672 14958
rect 4172 14900 4620 14906
rect 4172 14894 4672 14900
rect 4172 14890 4660 14894
rect 4160 14884 4660 14890
rect 4212 14878 4660 14884
rect 4160 14826 4212 14832
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3528 13954 3556 14350
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 3528 13926 3648 13954
rect 4080 13938 4108 14350
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 11694 1440 12718
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1964 12238 1992 12650
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 2884 12102 2912 12854
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2976 12306 3004 12650
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 3436 12238 3464 13126
rect 3528 12374 3556 13466
rect 3620 13462 3648 13926
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3608 13456 3660 13462
rect 3608 13398 3660 13404
rect 3896 13326 3924 13806
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3896 12442 3924 12582
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 3884 12436 3936 12442
rect 4724 12434 4752 14758
rect 4816 14618 4844 14962
rect 4908 14958 4936 16186
rect 4896 14952 4948 14958
rect 5000 14929 5028 17070
rect 4896 14894 4948 14900
rect 4986 14920 5042 14929
rect 4986 14855 5042 14864
rect 5092 14770 5120 19314
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18970 5764 19246
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5828 18766 5856 19858
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5184 18426 5212 18566
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5828 18290 5856 18702
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 5356 18216 5408 18222
rect 5408 18176 5488 18204
rect 5356 18158 5408 18164
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17746 5212 18022
rect 5460 17898 5488 18176
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5644 17898 5672 18090
rect 5460 17870 5672 17898
rect 5724 17876 5776 17882
rect 5460 17746 5488 17870
rect 5828 17864 5856 18226
rect 5776 17836 5856 17864
rect 5724 17818 5776 17824
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5184 17338 5212 17682
rect 5276 17610 5304 17682
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5276 17134 5304 17546
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5368 17116 5396 17614
rect 5552 17542 5580 17750
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5448 17128 5500 17134
rect 5368 17088 5448 17116
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16250 5212 16934
rect 5368 16794 5396 17088
rect 5448 17070 5500 17076
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5644 16658 5672 17002
rect 5264 16652 5316 16658
rect 5632 16652 5684 16658
rect 5264 16594 5316 16600
rect 5552 16612 5632 16640
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 4908 14742 5120 14770
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4908 13530 4936 14742
rect 4986 14648 5042 14657
rect 4986 14583 5042 14592
rect 5000 14346 5028 14583
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 13870 5120 14214
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4724 12406 4844 12434
rect 3884 12378 3936 12384
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2700 11694 2728 12038
rect 2884 11762 2912 12038
rect 3252 11898 3280 12174
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 3436 11694 3464 12038
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 4080 11694 4108 12174
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 1216 11552 1268 11558
rect 1216 11494 1268 11500
rect 1228 11218 1256 11494
rect 2700 11286 2728 11630
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 1216 11212 1268 11218
rect 1216 11154 1268 11160
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2424 10810 2452 11154
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2596 10600 2648 10606
rect 2700 10588 2728 11222
rect 4172 11150 4200 11630
rect 4264 11354 4292 11834
rect 4620 11688 4672 11694
rect 4672 11648 4752 11676
rect 4620 11630 4672 11636
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2648 10560 2728 10588
rect 2596 10542 2648 10548
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10130 2176 10406
rect 2792 10266 2820 10678
rect 2884 10606 2912 11018
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 4080 10742 4108 10950
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 10266 3188 10542
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 9518 1992 9862
rect 2792 9722 2820 10066
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2884 9586 2912 9862
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1216 9376 1268 9382
rect 1216 9318 1268 9324
rect 1228 9042 1256 9318
rect 1216 9036 1268 9042
rect 1216 8978 1268 8984
rect 1412 8498 1440 9454
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2516 8634 2544 8978
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 2608 8430 2636 9386
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8634 3280 8910
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 3252 8362 3280 8570
rect 3240 8356 3292 8362
rect 3344 8344 3372 10678
rect 4172 10606 4200 11086
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3436 8634 3464 9590
rect 3528 8974 3556 10134
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 4080 9024 4108 9862
rect 4160 9512 4212 9518
rect 4264 9500 4292 9998
rect 4724 9654 4752 11648
rect 4816 11014 4844 12406
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5000 11830 5028 12174
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4908 9518 4936 11018
rect 5092 10266 5120 13806
rect 5184 13734 5212 14826
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5276 12434 5304 16594
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5368 16046 5396 16458
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5552 15978 5580 16612
rect 5632 16594 5684 16600
rect 5828 16182 5856 17614
rect 5920 17066 5948 18770
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6012 18222 6040 18566
rect 6288 18426 6316 19858
rect 6932 19242 6960 20334
rect 7024 20058 7052 21354
rect 7208 21146 7236 21490
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12624 21344 12676 21350
rect 8942 21312 8998 21321
rect 12624 21286 12676 21292
rect 8942 21247 8998 21256
rect 8574 21176 8630 21185
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 8116 21140 8168 21146
rect 8956 21146 8984 21247
rect 12096 21244 12404 21253
rect 12096 21242 12102 21244
rect 12158 21242 12182 21244
rect 12238 21242 12262 21244
rect 12318 21242 12342 21244
rect 12398 21242 12404 21244
rect 12158 21190 12160 21242
rect 12340 21190 12342 21242
rect 12096 21188 12102 21190
rect 12158 21188 12182 21190
rect 12238 21188 12262 21190
rect 12318 21188 12342 21190
rect 12398 21188 12404 21190
rect 9770 21176 9826 21185
rect 12096 21179 12404 21188
rect 8574 21111 8576 21120
rect 8116 21082 8168 21088
rect 8628 21111 8630 21120
rect 8944 21140 8996 21146
rect 8576 21082 8628 21088
rect 9770 21111 9772 21120
rect 8944 21082 8996 21088
rect 9824 21111 9826 21120
rect 9772 21082 9824 21088
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7024 19854 7052 19994
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 7576 19174 7604 19450
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7760 18834 7788 19178
rect 7852 18873 7880 20742
rect 8128 20398 8156 21082
rect 12636 21010 12664 21286
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9496 21004 9548 21010
rect 9496 20946 9548 20952
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 7838 18864 7894 18873
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 7748 18828 7800 18834
rect 7838 18799 7894 18808
rect 7748 18770 7800 18776
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6472 18222 6500 18770
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6000 18216 6052 18222
rect 6184 18216 6236 18222
rect 6000 18158 6052 18164
rect 6104 18176 6184 18204
rect 6012 17882 6040 18158
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6012 17338 6040 17818
rect 6104 17746 6132 18176
rect 6184 18158 6236 18164
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6472 18086 6500 18158
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6196 17746 6224 18022
rect 6460 17808 6512 17814
rect 6644 17808 6696 17814
rect 6512 17768 6644 17796
rect 6460 17750 6512 17756
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 6196 17202 6224 17682
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6288 17134 6316 17478
rect 6380 17270 6408 17682
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 6000 17128 6052 17134
rect 6092 17128 6144 17134
rect 6000 17070 6052 17076
rect 6090 17096 6092 17105
rect 6276 17128 6328 17134
rect 6144 17096 6146 17105
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5920 16726 5948 17002
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 6012 16454 6040 17070
rect 6472 17105 6500 17614
rect 6276 17070 6328 17076
rect 6458 17096 6514 17105
rect 6090 17031 6146 17040
rect 6458 17031 6514 17040
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14618 5396 14758
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 13870 5396 14282
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5184 12406 5304 12434
rect 5184 11676 5212 12406
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5276 11830 5304 12242
rect 5368 11898 5396 13806
rect 5460 13802 5488 15506
rect 5552 14958 5580 15574
rect 5644 15094 5672 15982
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5736 15638 5764 15914
rect 6012 15706 6040 16390
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5632 15088 5684 15094
rect 5632 15030 5684 15036
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5552 14006 5580 14894
rect 5644 14385 5672 15030
rect 5630 14376 5686 14385
rect 5630 14311 5686 14320
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5920 13870 5948 14214
rect 6288 14074 6316 16730
rect 6564 16726 6592 17768
rect 6644 17750 6696 17756
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6748 17066 6776 17682
rect 6840 17354 6868 18022
rect 6932 17882 6960 18702
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6932 17542 6960 17818
rect 7104 17740 7156 17746
rect 7024 17700 7104 17728
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 7024 17354 7052 17700
rect 7104 17682 7156 17688
rect 6840 17326 7052 17354
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6748 16794 6776 17002
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6368 16720 6420 16726
rect 6368 16662 6420 16668
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 6380 16590 6408 16662
rect 6736 16652 6788 16658
rect 6840 16640 6868 17326
rect 6788 16612 6868 16640
rect 6736 16594 6788 16600
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6564 14822 6592 15982
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6656 15638 6684 15914
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 14414 6592 14758
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6380 14074 6408 14350
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6288 13870 6316 14010
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6748 13802 6776 16594
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15706 7328 15846
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 14890 6868 15302
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 7116 14482 7144 15438
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7116 13938 7144 14418
rect 7944 14414 7972 19382
rect 8036 19310 8064 19722
rect 8024 19304 8076 19310
rect 8220 19281 8248 20742
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8024 19246 8076 19252
rect 8206 19272 8262 19281
rect 8036 18426 8064 19246
rect 8206 19207 8262 19216
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8312 18222 8340 20334
rect 8864 19990 8892 20878
rect 9416 20534 9444 20946
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8404 18970 8432 19246
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8588 18630 8616 19246
rect 8680 18737 8708 19246
rect 8666 18728 8722 18737
rect 8864 18698 8892 19926
rect 9140 19922 9168 20198
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 8942 19408 8998 19417
rect 8942 19343 8998 19352
rect 9140 19366 9352 19394
rect 8956 19242 8984 19343
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 9140 18970 9168 19366
rect 9324 19310 9352 19366
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 8666 18663 8722 18672
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8956 18290 8984 18838
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9048 18358 9076 18770
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9232 18290 9260 19246
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9324 18834 9352 18906
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8312 17338 8340 18158
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8680 17746 8708 18022
rect 8772 17814 8800 18022
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8312 17202 8340 17274
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8036 16046 8064 17070
rect 8588 16182 8616 17682
rect 9324 16640 9352 18294
rect 9416 17066 9444 20470
rect 9508 20330 9536 20946
rect 9692 20602 9720 20946
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20641 11100 20742
rect 11058 20632 11114 20641
rect 9680 20596 9732 20602
rect 11058 20567 11114 20576
rect 9680 20538 9732 20544
rect 9954 20496 10010 20505
rect 9588 20460 9640 20466
rect 9954 20431 9956 20440
rect 9588 20402 9640 20408
rect 10008 20431 10010 20440
rect 9956 20402 10008 20408
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9600 20262 9628 20402
rect 9956 20324 10008 20330
rect 9956 20266 10008 20272
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9600 19514 9628 20198
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9692 19310 9720 19994
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9876 19310 9904 19858
rect 9968 19514 9996 20266
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9508 18086 9536 18634
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9600 17542 9628 18702
rect 9692 17814 9720 18702
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9784 16794 9812 18770
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10060 18426 10088 18702
rect 9864 18420 9916 18426
rect 10048 18420 10100 18426
rect 9916 18380 9996 18408
rect 9864 18362 9916 18368
rect 9968 18290 9996 18380
rect 10048 18362 10100 18368
rect 10152 18290 10180 20198
rect 11256 19786 11284 20946
rect 11436 20700 11744 20709
rect 11436 20698 11442 20700
rect 11498 20698 11522 20700
rect 11578 20698 11602 20700
rect 11658 20698 11682 20700
rect 11738 20698 11744 20700
rect 11498 20646 11500 20698
rect 11680 20646 11682 20698
rect 11436 20644 11442 20646
rect 11498 20644 11522 20646
rect 11578 20644 11602 20646
rect 11658 20644 11682 20646
rect 11738 20644 11744 20646
rect 11436 20635 11744 20644
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 11992 19922 12020 20198
rect 12096 20156 12404 20165
rect 12096 20154 12102 20156
rect 12158 20154 12182 20156
rect 12238 20154 12262 20156
rect 12318 20154 12342 20156
rect 12398 20154 12404 20156
rect 12158 20102 12160 20154
rect 12340 20102 12342 20154
rect 12096 20100 12102 20102
rect 12158 20100 12182 20102
rect 12238 20100 12262 20102
rect 12318 20100 12342 20102
rect 12398 20100 12404 20102
rect 12096 20091 12404 20100
rect 12544 19922 12572 20198
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10690 19408 10746 19417
rect 10690 19343 10746 19352
rect 10704 19310 10732 19343
rect 10324 19304 10376 19310
rect 10600 19304 10652 19310
rect 10376 19264 10456 19292
rect 10324 19246 10376 19252
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10244 18630 10272 18838
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9876 17882 9904 18090
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9876 17270 9904 17682
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9968 17202 9996 18022
rect 10046 17912 10102 17921
rect 10046 17847 10102 17856
rect 10060 17678 10088 17847
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10048 17128 10100 17134
rect 10152 17116 10180 18022
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10244 17134 10272 17818
rect 10336 17134 10364 18838
rect 10428 17241 10456 19264
rect 10600 19246 10652 19252
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10520 18970 10548 19178
rect 10612 18970 10640 19246
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10520 18834 10548 18906
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10520 17610 10548 18294
rect 10704 18222 10732 18702
rect 10888 18222 10916 19654
rect 11436 19612 11744 19621
rect 11436 19610 11442 19612
rect 11498 19610 11522 19612
rect 11578 19610 11602 19612
rect 11658 19610 11682 19612
rect 11738 19610 11744 19612
rect 11498 19558 11500 19610
rect 11680 19558 11682 19610
rect 11436 19556 11442 19558
rect 11498 19556 11522 19558
rect 11578 19556 11602 19558
rect 11658 19556 11682 19558
rect 11738 19556 11744 19558
rect 11436 19547 11744 19556
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10612 17785 10640 18158
rect 10704 17882 10732 18158
rect 10796 17921 10824 18158
rect 10782 17912 10838 17921
rect 10692 17876 10744 17882
rect 10782 17847 10838 17856
rect 10692 17818 10744 17824
rect 10598 17776 10654 17785
rect 10598 17711 10654 17720
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10414 17232 10470 17241
rect 10414 17167 10470 17176
rect 10100 17088 10180 17116
rect 10232 17128 10284 17134
rect 10048 17070 10100 17076
rect 10232 17070 10284 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9588 16652 9640 16658
rect 9324 16612 9588 16640
rect 9588 16594 9640 16600
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 9508 16046 9536 16186
rect 9784 16046 9812 16526
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9324 15910 9352 15982
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 8128 15570 8156 15846
rect 9048 15570 9076 15846
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 9692 14958 9720 15982
rect 9784 15706 9812 15982
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9876 15570 9904 16526
rect 10244 16114 10272 17070
rect 10428 16794 10456 17070
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10520 16674 10548 17546
rect 10612 17134 10640 17614
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10888 16794 10916 18158
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10428 16646 10548 16674
rect 11072 16658 11100 18838
rect 11992 18834 12020 19450
rect 12096 19068 12404 19077
rect 12096 19066 12102 19068
rect 12158 19066 12182 19068
rect 12238 19066 12262 19068
rect 12318 19066 12342 19068
rect 12398 19066 12404 19068
rect 12158 19014 12160 19066
rect 12340 19014 12342 19066
rect 12096 19012 12102 19014
rect 12158 19012 12182 19014
rect 12238 19012 12262 19014
rect 12318 19012 12342 19014
rect 12398 19012 12404 19014
rect 12096 19003 12404 19012
rect 12636 18902 12664 20402
rect 12820 20330 12848 21422
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12912 20602 12940 20878
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 13004 20398 13032 21286
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13268 20800 13320 20806
rect 13268 20742 13320 20748
rect 13280 20641 13308 20742
rect 13266 20632 13322 20641
rect 13266 20567 13322 20576
rect 13452 20528 13504 20534
rect 13188 20476 13452 20482
rect 13188 20470 13504 20476
rect 13188 20466 13492 20470
rect 13176 20460 13492 20466
rect 13228 20454 13492 20460
rect 13176 20402 13228 20408
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 13648 20330 13676 20810
rect 13924 20534 13952 21490
rect 18050 21448 18106 21457
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 17868 21412 17920 21418
rect 18050 21383 18052 21392
rect 17868 21354 17920 21360
rect 18104 21383 18106 21392
rect 18052 21354 18104 21360
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12820 18834 12848 20266
rect 13832 18902 13860 20266
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 11164 17882 11192 18770
rect 11436 18524 11744 18533
rect 11436 18522 11442 18524
rect 11498 18522 11522 18524
rect 11578 18522 11602 18524
rect 11658 18522 11682 18524
rect 11738 18522 11744 18524
rect 11498 18470 11500 18522
rect 11680 18470 11682 18522
rect 11436 18468 11442 18470
rect 11498 18468 11522 18470
rect 11578 18468 11602 18470
rect 11658 18468 11682 18470
rect 11738 18468 11744 18470
rect 11436 18459 11744 18468
rect 11808 18290 11836 18770
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11624 17882 11652 18158
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11612 17876 11664 17882
rect 11664 17836 11836 17864
rect 11612 17818 11664 17824
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11348 17542 11376 17682
rect 11612 17672 11664 17678
rect 11610 17640 11612 17649
rect 11664 17640 11666 17649
rect 11610 17575 11666 17584
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 17338 11376 17478
rect 11436 17436 11744 17445
rect 11436 17434 11442 17436
rect 11498 17434 11522 17436
rect 11578 17434 11602 17436
rect 11658 17434 11682 17436
rect 11738 17434 11744 17436
rect 11498 17382 11500 17434
rect 11680 17382 11682 17434
rect 11436 17380 11442 17382
rect 11498 17380 11522 17382
rect 11578 17380 11602 17382
rect 11658 17380 11682 17382
rect 11738 17380 11744 17382
rect 11436 17371 11744 17380
rect 11808 17338 11836 17836
rect 11992 17728 12020 18566
rect 12096 17980 12404 17989
rect 12096 17978 12102 17980
rect 12158 17978 12182 17980
rect 12238 17978 12262 17980
rect 12318 17978 12342 17980
rect 12398 17978 12404 17980
rect 12158 17926 12160 17978
rect 12340 17926 12342 17978
rect 12096 17924 12102 17926
rect 12158 17924 12182 17926
rect 12238 17924 12262 17926
rect 12318 17924 12342 17926
rect 12398 17924 12404 17926
rect 12096 17915 12404 17924
rect 12452 17882 12480 18770
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12072 17740 12124 17746
rect 11992 17700 12072 17728
rect 12072 17682 12124 17688
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11164 17134 11192 17206
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11426 17096 11482 17105
rect 11426 17031 11482 17040
rect 11704 17060 11756 17066
rect 11060 16652 11112 16658
rect 10428 16590 10456 16646
rect 11060 16594 11112 16600
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9876 15162 9904 15506
rect 9968 15162 9996 16050
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9968 15026 9996 15098
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8864 14482 8892 14758
rect 9048 14550 9076 14758
rect 9036 14544 9088 14550
rect 9036 14486 9088 14492
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 9324 13870 9352 14894
rect 9508 14074 9536 14894
rect 9692 14822 9720 14894
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 9312 13864 9364 13870
rect 9508 13841 9536 13874
rect 9312 13806 9364 13812
rect 9494 13832 9550 13841
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 5460 13394 5488 13738
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7208 13394 7236 13670
rect 7668 13530 7696 13670
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 5460 12782 5488 13330
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 12782 7144 13194
rect 8220 12850 8248 13398
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12442 6960 12582
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 5460 11694 5488 12106
rect 6196 12102 6224 12242
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 5552 11694 5580 12038
rect 5448 11688 5500 11694
rect 5184 11648 5304 11676
rect 5276 11082 5304 11648
rect 5448 11630 5500 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5552 10810 5580 11154
rect 5736 11150 5764 11630
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 5920 11354 5948 11494
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 6104 11218 6132 11494
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 6288 10674 6316 11086
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6380 10606 6408 11154
rect 7116 10674 7144 12718
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7576 11898 7604 12242
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 8036 11694 8064 12582
rect 8128 12442 8156 12718
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8312 12306 8340 13126
rect 8864 12782 8892 13126
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12374 8524 12582
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 6012 10130 6040 10406
rect 6104 10130 6132 10474
rect 6380 10266 6408 10542
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 5000 9654 5028 10066
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4212 9472 4292 9500
rect 4160 9454 4212 9460
rect 4080 8996 4200 9024
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3528 8362 3556 8774
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 3424 8356 3476 8362
rect 3344 8316 3424 8344
rect 3240 8298 3292 8304
rect 3424 8298 3476 8304
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7954 3004 8230
rect 4080 8022 4108 8842
rect 4172 8498 4200 8996
rect 4264 8838 4292 9472
rect 4620 9512 4672 9518
rect 4896 9512 4948 9518
rect 4672 9472 4752 9500
rect 4620 9454 4672 9460
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4356 8566 4384 8910
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4724 8294 4752 9472
rect 4896 9454 4948 9460
rect 5000 8974 5028 9590
rect 5092 9518 5120 9998
rect 5460 9738 5488 10066
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5368 9722 5488 9738
rect 5356 9716 5488 9722
rect 5408 9710 5488 9716
rect 5356 9658 5408 9664
rect 5644 9586 5672 9862
rect 5736 9722 5764 9998
rect 5920 9722 5948 10066
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5736 9586 5764 9658
rect 6012 9654 6040 9862
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 6012 9518 6040 9590
rect 6380 9518 6408 10066
rect 6840 9654 6868 10134
rect 7116 9722 7144 10610
rect 7852 10538 7880 10610
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 8220 10266 8248 11630
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8772 11354 8800 11562
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8772 10606 8800 10678
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 7116 9518 7144 9658
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7656 9512 7708 9518
rect 7944 9466 7972 10202
rect 8404 10198 8432 10406
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8680 9976 8708 10542
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8772 10130 8800 10406
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8864 10010 8892 11698
rect 8956 10130 8984 13806
rect 9494 13767 9496 13776
rect 9548 13767 9550 13776
rect 9496 13738 9548 13744
rect 9692 13394 9720 14758
rect 9954 13968 10010 13977
rect 9954 13903 10010 13912
rect 9968 13870 9996 13903
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 13394 10088 13738
rect 10336 13734 10364 15846
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10428 15366 10456 15642
rect 10520 15502 10548 16526
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10980 16046 11008 16458
rect 11072 16182 11100 16594
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15586 11008 15982
rect 10888 15570 11008 15586
rect 11072 15570 11100 16118
rect 11164 15706 11192 16594
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 10876 15564 11008 15570
rect 10928 15558 11008 15564
rect 10876 15506 10928 15512
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10520 14346 10548 15438
rect 10980 15366 11008 15558
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11256 15434 11284 16594
rect 11440 16522 11468 17031
rect 11808 17048 11836 17274
rect 11756 17020 11836 17048
rect 11704 17002 11756 17008
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11624 16658 11652 16934
rect 12096 16892 12404 16901
rect 12096 16890 12102 16892
rect 12158 16890 12182 16892
rect 12238 16890 12262 16892
rect 12318 16890 12342 16892
rect 12398 16890 12404 16892
rect 12158 16838 12160 16890
rect 12340 16838 12342 16890
rect 12096 16836 12102 16838
rect 12158 16836 12182 16838
rect 12238 16836 12262 16838
rect 12318 16836 12342 16838
rect 12398 16836 12404 16838
rect 12096 16827 12404 16836
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11436 16348 11744 16357
rect 11436 16346 11442 16348
rect 11498 16346 11522 16348
rect 11578 16346 11602 16348
rect 11658 16346 11682 16348
rect 11738 16346 11744 16348
rect 11498 16294 11500 16346
rect 11680 16294 11682 16346
rect 11436 16292 11442 16294
rect 11498 16292 11522 16294
rect 11578 16292 11602 16294
rect 11658 16292 11682 16294
rect 11738 16292 11744 16294
rect 11436 16283 11744 16292
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 11436 15260 11744 15269
rect 11436 15258 11442 15260
rect 11498 15258 11522 15260
rect 11578 15258 11602 15260
rect 11658 15258 11682 15260
rect 11738 15258 11744 15260
rect 11498 15206 11500 15258
rect 11680 15206 11682 15258
rect 11436 15204 11442 15206
rect 11498 15204 11522 15206
rect 11578 15204 11602 15206
rect 11658 15204 11682 15206
rect 11738 15204 11744 15206
rect 11436 15195 11744 15204
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11624 14958 11652 15098
rect 11808 14958 11836 16662
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11992 16046 12020 16526
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15570 11928 15846
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11992 14958 12020 15982
rect 12096 15804 12404 15813
rect 12096 15802 12102 15804
rect 12158 15802 12182 15804
rect 12238 15802 12262 15804
rect 12318 15802 12342 15804
rect 12398 15802 12404 15804
rect 12158 15750 12160 15802
rect 12340 15750 12342 15802
rect 12096 15748 12102 15750
rect 12158 15748 12182 15750
rect 12238 15748 12262 15750
rect 12318 15748 12342 15750
rect 12398 15748 12404 15750
rect 12096 15739 12404 15748
rect 12452 15638 12480 16594
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 11060 14952 11112 14958
rect 11612 14952 11664 14958
rect 11112 14900 11192 14906
rect 11060 14894 11192 14900
rect 11612 14894 11664 14900
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11072 14878 11192 14894
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10612 13870 10640 14010
rect 10980 13938 11008 14214
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11164 13870 11192 14878
rect 11624 14550 11652 14894
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11436 14172 11744 14181
rect 11436 14170 11442 14172
rect 11498 14170 11522 14172
rect 11578 14170 11602 14172
rect 11658 14170 11682 14172
rect 11738 14170 11744 14172
rect 11498 14118 11500 14170
rect 11680 14118 11682 14170
rect 11436 14116 11442 14118
rect 11498 14116 11522 14118
rect 11578 14116 11602 14118
rect 11658 14116 11682 14118
rect 11738 14116 11744 14118
rect 11436 14107 11744 14116
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10336 13394 10364 13670
rect 11072 13394 11100 13670
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 9324 12986 9352 13330
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9416 12850 9444 13262
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9140 11694 9168 12650
rect 9324 12434 9352 12718
rect 9496 12436 9548 12442
rect 9324 12406 9496 12434
rect 9496 12378 9548 12384
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11218 9168 11630
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11286 9352 11494
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9404 11212 9456 11218
rect 9508 11200 9536 12378
rect 10060 12374 10088 12718
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9876 11218 9904 12038
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9456 11172 9536 11200
rect 9404 11154 9456 11160
rect 9140 10742 9168 11154
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9048 10266 9076 10542
rect 9140 10266 9168 10678
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8760 9988 8812 9994
rect 8680 9948 8760 9976
rect 8864 9982 8984 10010
rect 8760 9930 8812 9936
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8312 9574 8524 9602
rect 8312 9518 8340 9574
rect 7708 9460 7972 9466
rect 7656 9454 7972 9460
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8430 4844 8774
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 5000 8090 5028 8910
rect 5736 8430 5764 9386
rect 5828 9178 5856 9454
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8498 5856 8774
rect 6012 8634 6040 8978
rect 6380 8838 6408 9454
rect 6472 9178 6500 9454
rect 7288 9444 7340 9450
rect 7668 9438 7972 9454
rect 7288 9386 7340 9392
rect 7300 9178 7328 9386
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8294 5764 8366
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 6840 7206 6868 7822
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7342 7604 7686
rect 7760 7546 7788 7890
rect 7944 7886 7972 9438
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9042 8248 9318
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8312 8430 8340 9046
rect 8404 8634 8432 9454
rect 8496 9042 8524 9574
rect 8772 9110 8800 9658
rect 8864 9450 8892 9862
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 7970 8340 8366
rect 8220 7954 8340 7970
rect 8208 7948 8340 7954
rect 8260 7942 8340 7948
rect 8208 7890 8260 7896
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 6840 6934 6868 7142
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2044 6180 2096 6186
rect 2044 6122 2096 6128
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1964 4826 1992 5034
rect 2056 5030 2084 6122
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 5778 2912 6054
rect 2976 5778 3004 6734
rect 3160 5914 3188 6802
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3528 6390 3556 6598
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 4080 5846 4108 6598
rect 4264 6118 4292 6870
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6118 4936 6734
rect 5184 6118 5212 6802
rect 6840 6254 6868 6870
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 7116 6186 7144 6802
rect 7944 6254 7972 7822
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8588 7342 8616 7754
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 6934 8616 7278
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6254 8064 6598
rect 8404 6458 8432 6802
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 4264 5846 4292 6054
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4908 5914 4936 6054
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2056 4690 2084 4966
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 1780 4593 1808 4626
rect 1766 4584 1822 4593
rect 1766 4519 1822 4528
rect 2056 4078 2084 4626
rect 2332 4622 2360 5646
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2686 4584 2742 4593
rect 2332 4128 2360 4558
rect 2686 4519 2742 4528
rect 2700 4486 2728 4519
rect 2688 4480 2740 4486
rect 2884 4468 2912 5714
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3252 5098 3280 5646
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3344 5030 3372 5510
rect 3436 5370 3464 5646
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3436 4826 3464 5102
rect 3528 4826 3556 5646
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3620 4554 3648 5306
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3804 4690 3832 5034
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4826 4016 4966
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 2740 4440 2912 4468
rect 4068 4480 4120 4486
rect 2688 4422 2740 4428
rect 4172 4468 4200 5782
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4724 5166 4752 5578
rect 4908 5234 4936 5850
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4120 4440 4200 4468
rect 4068 4422 4120 4428
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 4080 4282 4108 4422
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 2504 4140 2556 4146
rect 2332 4100 2504 4128
rect 2504 4082 2556 4088
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3602 1808 3878
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 2056 2922 2084 4014
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 2990 2268 3878
rect 2700 3670 2728 4150
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2044 2916 2096 2922
rect 2044 2858 2096 2864
rect 2884 2774 2912 4014
rect 3344 3738 3372 4014
rect 3436 3738 3464 4150
rect 4080 4146 4108 4218
rect 4264 4214 4292 4694
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4540 4214 4568 4422
rect 4724 4214 4752 4422
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3436 2922 3464 3538
rect 3988 3534 4016 3878
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 2884 2746 3004 2774
rect 2976 2650 3004 2746
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3436 2514 3464 2858
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3528 2514 3556 2790
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 4080 2446 4108 4082
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4172 3194 4200 3878
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4724 3058 4752 4150
rect 4908 4078 4936 4694
rect 5184 4690 5212 6054
rect 7944 5778 7972 6190
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4908 3942 4936 4014
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4908 2990 4936 3878
rect 5000 3398 5028 4014
rect 5092 3670 5120 4422
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 3126 5028 3334
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4896 2984 4948 2990
rect 5184 2938 5212 4626
rect 5552 4622 5580 5510
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5644 4146 5672 5306
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5828 5030 5856 5170
rect 5920 5166 5948 5578
rect 6288 5234 6316 5646
rect 7944 5302 7972 5714
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 8128 5166 8156 6054
rect 8404 5846 8432 6054
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8588 5778 8616 6870
rect 8680 6866 8708 7686
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8772 7002 8800 7210
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8680 5914 8708 6122
rect 8772 5914 8800 6938
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6092 5160 6144 5166
rect 8116 5160 8168 5166
rect 6144 5120 6224 5148
rect 6092 5102 6144 5108
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 6196 4146 6224 5120
rect 8116 5102 8168 5108
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4690 7880 4966
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3058 5488 3334
rect 5552 3194 5580 4082
rect 5644 3534 5672 4082
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6012 3942 6040 4014
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 4896 2926 4948 2932
rect 5092 2910 5212 2938
rect 6092 2916 6144 2922
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4252 1760 4304 1766
rect 4252 1702 4304 1708
rect 4264 1426 4292 1702
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 4724 1494 4752 2246
rect 5092 1834 5120 2910
rect 6092 2858 6144 2864
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 5184 1902 5212 2790
rect 6012 2514 6040 2790
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 5080 1828 5132 1834
rect 5080 1770 5132 1776
rect 4712 1488 4764 1494
rect 4712 1430 4764 1436
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 5460 1290 5488 2450
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5828 1358 5856 2382
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 5448 1284 5500 1290
rect 5448 1226 5500 1232
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 5828 882 5856 1294
rect 6012 1222 6040 2450
rect 6104 2378 6132 2858
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6092 1828 6144 1834
rect 6092 1770 6144 1776
rect 6104 1426 6132 1770
rect 6092 1420 6144 1426
rect 6092 1362 6144 1368
rect 6196 1358 6224 3062
rect 6380 2514 6408 3130
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6472 2650 6500 2926
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6748 2582 6776 2926
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6380 2106 6408 2450
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6840 1970 6868 2314
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 6840 1562 6868 1906
rect 6828 1556 6880 1562
rect 6828 1498 6880 1504
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 6000 1216 6052 1222
rect 6000 1158 6052 1164
rect 6932 1018 6960 2926
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7024 2650 7052 2858
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7116 1850 7144 2790
rect 7944 2446 7972 3470
rect 8128 3058 8156 5102
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 3942 8708 4966
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8496 3602 8524 3878
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8772 3534 8800 5714
rect 8864 5166 8892 7346
rect 8956 6730 8984 9982
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 9048 7410 9076 9930
rect 9140 9382 9168 10202
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9324 8430 9352 10542
rect 9508 10538 9536 11172
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9876 10810 9904 11154
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10810 9996 10950
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9876 10606 9904 10746
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9508 10130 9536 10474
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9416 9178 9444 10066
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6866 9260 7142
rect 9692 6866 9720 9998
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 9042 9812 9318
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9862 7984 9918 7993
rect 9862 7919 9864 7928
rect 9916 7919 9918 7928
rect 9864 7890 9916 7896
rect 9772 7336 9824 7342
rect 9876 7324 9904 7890
rect 9824 7296 9904 7324
rect 9772 7278 9824 7284
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8864 4282 8892 5102
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 9048 4978 9076 6802
rect 9232 5710 9260 6802
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9600 6458 9628 6666
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9600 5778 9628 5850
rect 10060 5778 10088 11290
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 10152 9450 10180 9862
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10336 9110 10364 13330
rect 11164 12442 11192 13806
rect 11256 12850 11284 13942
rect 11808 13394 11836 14418
rect 11992 13870 12020 14894
rect 12096 14716 12404 14725
rect 12096 14714 12102 14716
rect 12158 14714 12182 14716
rect 12238 14714 12262 14716
rect 12318 14714 12342 14716
rect 12398 14714 12404 14716
rect 12158 14662 12160 14714
rect 12340 14662 12342 14714
rect 12096 14660 12102 14662
rect 12158 14660 12182 14662
rect 12238 14660 12262 14662
rect 12318 14660 12342 14662
rect 12398 14660 12404 14662
rect 12096 14651 12404 14660
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11900 13530 11928 13738
rect 12096 13628 12404 13637
rect 12096 13626 12102 13628
rect 12158 13626 12182 13628
rect 12238 13626 12262 13628
rect 12318 13626 12342 13628
rect 12398 13626 12404 13628
rect 12158 13574 12160 13626
rect 12340 13574 12342 13626
rect 12096 13572 12102 13574
rect 12158 13572 12182 13574
rect 12238 13572 12262 13574
rect 12318 13572 12342 13574
rect 12398 13572 12404 13574
rect 12096 13563 12404 13572
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11436 13084 11744 13093
rect 11436 13082 11442 13084
rect 11498 13082 11522 13084
rect 11578 13082 11602 13084
rect 11658 13082 11682 13084
rect 11738 13082 11744 13084
rect 11498 13030 11500 13082
rect 11680 13030 11682 13082
rect 11436 13028 11442 13030
rect 11498 13028 11522 13030
rect 11578 13028 11602 13030
rect 11658 13028 11682 13030
rect 11738 13028 11744 13030
rect 11436 13019 11744 13028
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10428 9722 10456 10474
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10130 10640 10406
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10704 7954 10732 9454
rect 11072 9450 11100 12310
rect 11164 11694 11192 12378
rect 11256 12306 11284 12582
rect 11716 12306 11744 12650
rect 11808 12306 11836 13330
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12424 12020 12718
rect 12096 12540 12404 12549
rect 12096 12538 12102 12540
rect 12158 12538 12182 12540
rect 12238 12538 12262 12540
rect 12318 12538 12342 12540
rect 12398 12538 12404 12540
rect 12158 12486 12160 12538
rect 12340 12486 12342 12538
rect 12096 12484 12102 12486
rect 12158 12484 12182 12486
rect 12238 12484 12262 12486
rect 12318 12484 12342 12486
rect 12398 12484 12404 12486
rect 12096 12475 12404 12484
rect 11992 12396 12204 12424
rect 12176 12306 12204 12396
rect 11244 12300 11296 12306
rect 11704 12300 11756 12306
rect 11296 12260 11376 12288
rect 11244 12242 11296 12248
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11256 10554 11284 12038
rect 11348 11694 11376 12260
rect 11704 12242 11756 12248
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 11436 11996 11744 12005
rect 11436 11994 11442 11996
rect 11498 11994 11522 11996
rect 11578 11994 11602 11996
rect 11658 11994 11682 11996
rect 11738 11994 11744 11996
rect 11498 11942 11500 11994
rect 11680 11942 11682 11994
rect 11436 11940 11442 11942
rect 11498 11940 11522 11942
rect 11578 11940 11602 11942
rect 11658 11940 11682 11942
rect 11738 11940 11744 11942
rect 11436 11931 11744 11940
rect 12084 11762 12112 12242
rect 12452 11898 12480 15574
rect 12544 15502 12572 17682
rect 12636 17134 12664 18022
rect 12728 17814 12756 18566
rect 13004 18222 13032 18702
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 13096 18222 13124 18634
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 12912 18057 12940 18158
rect 12898 18048 12954 18057
rect 12898 17983 12954 17992
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 13372 17610 13400 18158
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13648 17814 13676 18022
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13740 17134 13768 18770
rect 13924 18222 13952 19178
rect 14016 19174 14044 21286
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14200 20262 14228 20742
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14280 20528 14332 20534
rect 14278 20496 14280 20505
rect 14332 20496 14334 20505
rect 14278 20431 14334 20440
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14292 19786 14320 20334
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19378 14136 19654
rect 14292 19514 14320 19722
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14568 18766 14596 20538
rect 14660 20534 14688 21354
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16868 21010 16896 21286
rect 17880 21146 17908 21354
rect 18064 21146 18092 21354
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 17868 21140 17920 21146
rect 18052 21140 18104 21146
rect 17920 21100 18000 21128
rect 17868 21082 17920 21088
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 15198 20904 15254 20913
rect 14844 20602 14872 20878
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14660 20058 14688 20470
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14844 19689 14872 19858
rect 14830 19680 14886 19689
rect 14830 19615 14886 19624
rect 14936 19378 14964 20878
rect 15198 20839 15254 20848
rect 15212 20806 15240 20839
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 16210 20768 16266 20777
rect 15212 20466 15240 20742
rect 16210 20703 16266 20712
rect 15474 20632 15530 20641
rect 15474 20567 15530 20576
rect 15488 20534 15516 20567
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 16224 20466 16252 20703
rect 16486 20632 16542 20641
rect 17144 20602 17172 20946
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 16486 20567 16488 20576
rect 16540 20567 16542 20576
rect 17132 20596 17184 20602
rect 16488 20538 16540 20544
rect 17132 20538 17184 20544
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 15856 20369 15884 20402
rect 15842 20360 15898 20369
rect 15292 20324 15344 20330
rect 15842 20295 15898 20304
rect 15292 20266 15344 20272
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15212 19990 15240 20198
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14740 19304 14792 19310
rect 15016 19304 15068 19310
rect 14740 19246 14792 19252
rect 15014 19272 15016 19281
rect 15068 19272 15070 19281
rect 14752 18970 14780 19246
rect 15014 19207 15070 19216
rect 15212 18970 15240 19926
rect 15304 19786 15332 20266
rect 15566 20088 15622 20097
rect 15396 20046 15566 20074
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15396 19334 15424 20046
rect 15566 20023 15622 20032
rect 15580 19922 15608 20023
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15488 19718 15516 19858
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15304 19306 15424 19334
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13924 17134 13952 18158
rect 14200 17134 14228 18226
rect 14738 18048 14794 18057
rect 14738 17983 14794 17992
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14372 17536 14424 17542
rect 14278 17504 14334 17513
rect 14372 17478 14424 17484
rect 14278 17439 14334 17448
rect 14292 17202 14320 17439
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 13740 16726 13768 17070
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 14200 16046 14228 17070
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15638 13124 15846
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 14346 12572 15438
rect 13280 14958 13308 15982
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15570 13584 15846
rect 14016 15706 14044 15982
rect 14200 15706 14228 15982
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14096 15564 14148 15570
rect 14292 15552 14320 17138
rect 14384 17134 14412 17478
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14148 15524 14320 15552
rect 14096 15506 14148 15512
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13740 15162 13768 15438
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13728 15020 13780 15026
rect 13832 15008 13860 15506
rect 14016 15162 14044 15506
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 14108 15026 14136 15370
rect 13780 14980 13860 15008
rect 14096 15020 14148 15026
rect 13728 14962 13780 14968
rect 14096 14962 14148 14968
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12912 14618 12940 14894
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12544 14074 12572 14282
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12544 12782 12572 13262
rect 12636 12782 12664 14418
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12782 12756 13126
rect 12912 12850 12940 13466
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12716 12776 12768 12782
rect 13004 12753 13032 14418
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12716 12718 12768 12724
rect 12990 12744 13046 12753
rect 12636 12434 12664 12718
rect 13096 12714 13124 14350
rect 13188 13258 13216 14826
rect 13280 13376 13308 14894
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13372 14550 13400 14758
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13464 13394 13492 14962
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13648 14482 13676 14894
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13832 14482 13860 14826
rect 14200 14822 14228 15524
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 14958 14412 15302
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14476 14890 14504 17682
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 16794 14596 17614
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 13648 13841 13676 14418
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 14074 13768 14350
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13726 13968 13782 13977
rect 13726 13903 13782 13912
rect 13634 13832 13690 13841
rect 13634 13767 13690 13776
rect 13648 13530 13676 13767
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13740 13462 13768 13903
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13360 13388 13412 13394
rect 13280 13348 13360 13376
rect 13360 13330 13412 13336
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13372 13190 13400 13330
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13268 12776 13320 12782
rect 13372 12764 13400 13126
rect 13452 12776 13504 12782
rect 13372 12736 13452 12764
rect 13268 12718 13320 12724
rect 13452 12718 13504 12724
rect 12990 12679 13046 12688
rect 13084 12708 13136 12714
rect 12544 12406 12664 12434
rect 12544 12170 12572 12406
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12544 12050 12572 12106
rect 12912 12050 12940 12242
rect 12544 12022 12940 12050
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11436 10908 11744 10917
rect 11436 10906 11442 10908
rect 11498 10906 11522 10908
rect 11578 10906 11602 10908
rect 11658 10906 11682 10908
rect 11738 10906 11744 10908
rect 11498 10854 11500 10906
rect 11680 10854 11682 10906
rect 11436 10852 11442 10854
rect 11498 10852 11522 10854
rect 11578 10852 11602 10854
rect 11658 10852 11682 10854
rect 11738 10852 11744 10854
rect 11436 10843 11744 10852
rect 11164 10526 11468 10554
rect 11164 10198 11192 10526
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 10198 11284 10406
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9926 11376 10066
rect 11440 10062 11468 10526
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11436 9820 11744 9829
rect 11436 9818 11442 9820
rect 11498 9818 11522 9820
rect 11578 9818 11602 9820
rect 11658 9818 11682 9820
rect 11738 9818 11744 9820
rect 11498 9766 11500 9818
rect 11680 9766 11682 9818
rect 11436 9764 11442 9766
rect 11498 9764 11522 9766
rect 11578 9764 11602 9766
rect 11658 9764 11682 9766
rect 11738 9764 11744 9766
rect 11436 9755 11744 9764
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 8294 11100 9386
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 9042 11652 9318
rect 11704 9172 11756 9178
rect 11808 9160 11836 11494
rect 12096 11452 12404 11461
rect 12096 11450 12102 11452
rect 12158 11450 12182 11452
rect 12238 11450 12262 11452
rect 12318 11450 12342 11452
rect 12398 11450 12404 11452
rect 12158 11398 12160 11450
rect 12340 11398 12342 11450
rect 12096 11396 12102 11398
rect 12158 11396 12182 11398
rect 12238 11396 12262 11398
rect 12318 11396 12342 11398
rect 12398 11396 12404 11398
rect 12096 11387 12404 11396
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11992 10266 12020 10474
rect 12096 10364 12404 10373
rect 12096 10362 12102 10364
rect 12158 10362 12182 10364
rect 12238 10362 12262 10364
rect 12318 10362 12342 10364
rect 12398 10362 12404 10364
rect 12158 10310 12160 10362
rect 12340 10310 12342 10362
rect 12096 10308 12102 10310
rect 12158 10308 12182 10310
rect 12238 10308 12262 10310
rect 12318 10308 12342 10310
rect 12398 10308 12404 10310
rect 12096 10299 12404 10308
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11900 9674 11928 10202
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11900 9646 12020 9674
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11756 9132 11836 9160
rect 11704 9114 11756 9120
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11436 8732 11744 8741
rect 11436 8730 11442 8732
rect 11498 8730 11522 8732
rect 11578 8730 11602 8732
rect 11658 8730 11682 8732
rect 11738 8730 11744 8732
rect 11498 8678 11500 8730
rect 11680 8678 11682 8730
rect 11436 8676 11442 8678
rect 11498 8676 11522 8678
rect 11578 8676 11602 8678
rect 11658 8676 11682 8678
rect 11738 8676 11744 8678
rect 11436 8667 11744 8676
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10152 7342 10180 7890
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10244 7342 10272 7822
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10704 6866 10732 7686
rect 10888 7342 10916 7686
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6866 11100 7142
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11164 6458 11192 7210
rect 11348 6934 11376 8230
rect 11716 7954 11744 8230
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11436 7644 11744 7653
rect 11436 7642 11442 7644
rect 11498 7642 11522 7644
rect 11578 7642 11602 7644
rect 11658 7642 11682 7644
rect 11738 7642 11744 7644
rect 11498 7590 11500 7642
rect 11680 7590 11682 7642
rect 11436 7588 11442 7590
rect 11498 7588 11522 7590
rect 11578 7588 11602 7590
rect 11658 7588 11682 7590
rect 11738 7588 11744 7590
rect 11436 7579 11744 7588
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11348 6746 11376 6870
rect 11532 6866 11560 7482
rect 11808 7290 11836 9132
rect 11900 9110 11928 9318
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11992 7886 12020 9646
rect 12084 9518 12112 9862
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12096 9276 12404 9285
rect 12096 9274 12102 9276
rect 12158 9274 12182 9276
rect 12238 9274 12262 9276
rect 12318 9274 12342 9276
rect 12398 9274 12404 9276
rect 12158 9222 12160 9274
rect 12340 9222 12342 9274
rect 12096 9220 12102 9222
rect 12158 9220 12182 9222
rect 12238 9220 12262 9222
rect 12318 9220 12342 9222
rect 12398 9220 12404 9222
rect 12096 9211 12404 9220
rect 12096 8188 12404 8197
rect 12096 8186 12102 8188
rect 12158 8186 12182 8188
rect 12238 8186 12262 8188
rect 12318 8186 12342 8188
rect 12398 8186 12404 8188
rect 12158 8134 12160 8186
rect 12340 8134 12342 8186
rect 12096 8132 12102 8134
rect 12158 8132 12182 8134
rect 12238 8132 12262 8134
rect 12318 8132 12342 8134
rect 12398 8132 12404 8134
rect 12096 8123 12404 8132
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11900 7410 11928 7822
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 12084 7290 12112 7958
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7478 12296 7686
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12452 7342 12480 11834
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 9178 12572 9454
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12636 8090 12664 11494
rect 12808 9988 12860 9994
rect 13004 9976 13032 12679
rect 13084 12650 13136 12656
rect 13096 11694 13124 12650
rect 13280 12306 13308 12718
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13464 10538 13492 12718
rect 13740 12714 13768 13398
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13096 10130 13124 10474
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 10130 13216 10406
rect 13648 10198 13676 12378
rect 13832 12102 13860 12854
rect 14016 12838 14320 12866
rect 14016 12782 14044 12838
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13740 10130 13768 10542
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 12860 9948 13032 9976
rect 12808 9930 12860 9936
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 9042 12756 9454
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12544 7546 12572 7958
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 11808 7262 12112 7290
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11256 6718 11376 6746
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11256 5778 11284 6718
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9416 5642 9444 5714
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9140 5166 9168 5510
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9508 5098 9536 5714
rect 11348 5370 11376 6598
rect 11436 6556 11744 6565
rect 11436 6554 11442 6556
rect 11498 6554 11522 6556
rect 11578 6554 11602 6556
rect 11658 6554 11682 6556
rect 11738 6554 11744 6556
rect 11498 6502 11500 6554
rect 11680 6502 11682 6554
rect 11436 6500 11442 6502
rect 11498 6500 11522 6502
rect 11578 6500 11602 6502
rect 11658 6500 11682 6502
rect 11738 6500 11744 6502
rect 11436 6491 11744 6500
rect 11808 6186 11836 7262
rect 12096 7100 12404 7109
rect 12096 7098 12102 7100
rect 12158 7098 12182 7100
rect 12238 7098 12262 7100
rect 12318 7098 12342 7100
rect 12398 7098 12404 7100
rect 12158 7046 12160 7098
rect 12340 7046 12342 7098
rect 12096 7044 12102 7046
rect 12158 7044 12182 7046
rect 12238 7044 12262 7046
rect 12318 7044 12342 7046
rect 12398 7044 12404 7046
rect 12096 7035 12404 7044
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6458 12204 6598
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12176 6254 12204 6394
rect 12360 6390 12388 6870
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12452 6322 12480 7278
rect 12544 7002 12572 7482
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12544 6254 12572 6938
rect 12820 6866 12848 9930
rect 13464 9722 13492 10066
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 8430 13584 8774
rect 13740 8430 13768 10066
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 7886 13032 8230
rect 13740 7954 13768 8366
rect 14016 7993 14044 12582
rect 14108 12442 14136 12718
rect 14096 12436 14148 12442
rect 14292 12424 14320 12838
rect 14384 12782 14412 13126
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14372 12436 14424 12442
rect 14292 12396 14372 12424
rect 14096 12378 14148 12384
rect 14372 12378 14424 12384
rect 14568 12306 14596 14418
rect 14660 13938 14688 15302
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14660 13444 14688 13874
rect 14752 13870 14780 17983
rect 14936 17746 14964 18770
rect 15198 18320 15254 18329
rect 15198 18255 15254 18264
rect 15014 18184 15070 18193
rect 15014 18119 15016 18128
rect 15068 18119 15070 18128
rect 15016 18090 15068 18096
rect 15028 17882 15056 18090
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 15212 17746 15240 18255
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 14844 16726 14872 17206
rect 14936 17134 14964 17478
rect 15212 17202 15240 17478
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14936 15570 14964 15914
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14844 14618 14872 15506
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 15014 14376 15070 14385
rect 15014 14311 15070 14320
rect 15028 14074 15056 14311
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14740 13456 14792 13462
rect 14660 13416 14740 13444
rect 14740 13398 14792 13404
rect 14556 12300 14608 12306
rect 14476 12260 14556 12288
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10606 14320 10950
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 9926 14320 10542
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 9518 14320 9862
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14476 9042 14504 12260
rect 14556 12242 14608 12248
rect 14936 11354 14964 13942
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15120 12889 15148 12922
rect 15106 12880 15162 12889
rect 15106 12815 15162 12824
rect 15304 12306 15332 19306
rect 15488 18358 15516 19654
rect 15856 19446 15884 20295
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15580 18358 15608 18770
rect 15672 18766 15700 19110
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15672 18170 15700 18702
rect 15764 18222 15792 18906
rect 15948 18834 15976 19314
rect 16040 19242 16068 19722
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15936 18828 15988 18834
rect 15856 18788 15936 18816
rect 15856 18630 15884 18788
rect 15936 18770 15988 18776
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15856 18222 15884 18566
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15580 18142 15700 18170
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15580 17746 15608 18142
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15672 17746 15700 18022
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15580 15638 15608 17682
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 14822 15792 15438
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14482 15792 14758
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15396 12170 15424 13330
rect 15488 12782 15516 13738
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15580 12986 15608 13126
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15476 12776 15528 12782
rect 15528 12736 15608 12764
rect 15476 12718 15528 12724
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15488 11762 15516 12582
rect 15580 12442 15608 12736
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15764 12374 15792 14418
rect 15752 12368 15804 12374
rect 15566 12336 15622 12345
rect 15752 12310 15804 12316
rect 15566 12271 15622 12280
rect 15660 12300 15712 12306
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15212 10606 15240 11494
rect 15580 11354 15608 12271
rect 15660 12242 15712 12248
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 9586 14596 10406
rect 14660 10266 14688 10542
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 15014 10160 15070 10169
rect 15212 10130 15240 10542
rect 15014 10095 15016 10104
rect 15068 10095 15070 10104
rect 15200 10124 15252 10130
rect 15016 10066 15068 10072
rect 15200 10066 15252 10072
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14568 9110 14596 9386
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 9178 14780 9318
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14002 7984 14058 7993
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13728 7948 13780 7954
rect 14002 7919 14058 7928
rect 13728 7890 13780 7896
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13096 7410 13124 7822
rect 13188 7410 13216 7890
rect 14292 7886 14320 8842
rect 14568 8090 14596 9046
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 8430 14872 8774
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 15028 8129 15056 10066
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 9602 15148 9862
rect 15120 9574 15240 9602
rect 15212 9450 15240 9574
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15014 8120 15070 8129
rect 14556 8084 14608 8090
rect 15014 8055 15016 8064
rect 14556 8026 14608 8032
rect 15068 8055 15070 8064
rect 15016 8026 15068 8032
rect 14568 7993 14596 8026
rect 14648 8016 14700 8022
rect 14554 7984 14610 7993
rect 14700 7976 14780 8004
rect 14648 7958 14700 7964
rect 14554 7919 14610 7928
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13096 6866 13124 7346
rect 13464 6866 13492 7686
rect 13740 7410 13768 7686
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 14016 7342 14044 7686
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 6934 13860 7210
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 12808 6860 12860 6866
rect 13084 6860 13136 6866
rect 12808 6802 12860 6808
rect 13004 6820 13084 6848
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11436 5468 11744 5477
rect 11436 5466 11442 5468
rect 11498 5466 11522 5468
rect 11578 5466 11602 5468
rect 11658 5466 11682 5468
rect 11738 5466 11744 5468
rect 11498 5414 11500 5466
rect 11680 5414 11682 5466
rect 11436 5412 11442 5414
rect 11498 5412 11522 5414
rect 11578 5412 11602 5414
rect 11658 5412 11682 5414
rect 11738 5412 11744 5414
rect 11436 5403 11744 5412
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11808 5114 11836 6122
rect 12096 6012 12404 6021
rect 12096 6010 12102 6012
rect 12158 6010 12182 6012
rect 12238 6010 12262 6012
rect 12318 6010 12342 6012
rect 12398 6010 12404 6012
rect 12158 5958 12160 6010
rect 12340 5958 12342 6010
rect 12096 5956 12102 5958
rect 12158 5956 12182 5958
rect 12238 5956 12262 5958
rect 12318 5956 12342 5958
rect 12398 5956 12404 5958
rect 12096 5947 12404 5956
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 5370 12204 5510
rect 12530 5400 12586 5409
rect 12164 5364 12216 5370
rect 12530 5335 12532 5344
rect 12164 5306 12216 5312
rect 12584 5335 12586 5344
rect 12532 5306 12584 5312
rect 12440 5160 12492 5166
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 8956 4758 8984 4966
rect 9048 4950 9168 4978
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 9140 4214 9168 4950
rect 9508 4826 9536 5034
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8496 2922 8524 3334
rect 8956 2990 8984 3402
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7300 2106 7328 2382
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7024 1822 7144 1850
rect 7024 1494 7052 1822
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 7012 1488 7064 1494
rect 7012 1430 7064 1436
rect 6920 1012 6972 1018
rect 6920 954 6972 960
rect 5816 876 5868 882
rect 5816 818 5868 824
rect 7116 814 7144 1702
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 7208 1018 7236 1294
rect 7484 1290 7512 2382
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 8036 1494 8064 2042
rect 8312 1970 8340 2382
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8312 1562 8340 1906
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 8024 1488 8076 1494
rect 8024 1430 8076 1436
rect 7472 1284 7524 1290
rect 7472 1226 7524 1232
rect 7196 1012 7248 1018
rect 7196 954 7248 960
rect 7104 808 7156 814
rect 7104 750 7156 756
rect 7484 746 7512 1226
rect 8036 1018 8064 1430
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8024 1012 8076 1018
rect 8024 954 8076 960
rect 8404 814 8432 1362
rect 8588 1222 8616 2790
rect 8956 2310 8984 2926
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8852 1828 8904 1834
rect 8852 1770 8904 1776
rect 8864 1562 8892 1770
rect 8852 1556 8904 1562
rect 8852 1498 8904 1504
rect 8668 1488 8720 1494
rect 8956 1442 8984 2246
rect 8668 1430 8720 1436
rect 8576 1216 8628 1222
rect 8576 1158 8628 1164
rect 8588 882 8616 1158
rect 8680 1018 8708 1430
rect 8864 1426 8984 1442
rect 9048 1426 9076 2994
rect 9140 2446 9168 4150
rect 9508 4146 9536 4762
rect 10980 4690 11008 4966
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 11164 4078 11192 5102
rect 11808 5086 11928 5114
rect 12440 5102 12492 5108
rect 11900 5030 11928 5086
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11256 4758 11284 4966
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11436 4380 11744 4389
rect 11436 4378 11442 4380
rect 11498 4378 11522 4380
rect 11578 4378 11602 4380
rect 11658 4378 11682 4380
rect 11738 4378 11744 4380
rect 11498 4326 11500 4378
rect 11680 4326 11682 4378
rect 11436 4324 11442 4326
rect 11498 4324 11522 4326
rect 11578 4324 11602 4326
rect 11658 4324 11682 4326
rect 11738 4324 11744 4326
rect 11436 4315 11744 4324
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3194 9352 3878
rect 9600 3210 9628 4014
rect 11808 4010 11836 4966
rect 11900 4758 11928 4966
rect 12096 4924 12404 4933
rect 12096 4922 12102 4924
rect 12158 4922 12182 4924
rect 12238 4922 12262 4924
rect 12318 4922 12342 4924
rect 12398 4922 12404 4924
rect 12158 4870 12160 4922
rect 12340 4870 12342 4922
rect 12096 4868 12102 4870
rect 12158 4868 12182 4870
rect 12238 4868 12262 4870
rect 12318 4868 12342 4870
rect 12398 4868 12404 4870
rect 12096 4859 12404 4868
rect 12452 4826 12480 5102
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 12544 4554 12572 5306
rect 12820 5098 12848 6190
rect 13004 5846 13032 6820
rect 13084 6802 13136 6808
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 14476 6798 14504 7482
rect 14568 7206 14596 7919
rect 14752 7546 14780 7976
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 15028 6322 15056 7890
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12820 4758 12848 5034
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12912 4690 12940 5578
rect 13004 5234 13032 5782
rect 13188 5710 13216 6122
rect 13280 5778 13308 6122
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5370 13124 5510
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4690 13032 4966
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 12636 3942 12664 4422
rect 13188 4078 13216 5646
rect 13648 5166 13676 5782
rect 13924 5370 13952 6054
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 13648 4690 13676 5102
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13832 4078 13860 4966
rect 14292 4758 14320 4966
rect 14384 4826 14412 5102
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14384 4486 14412 4626
rect 14476 4554 14504 5306
rect 15212 5234 15240 9386
rect 15672 9042 15700 12242
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 15764 11150 15792 12106
rect 15856 12102 15884 18022
rect 15948 17882 15976 18226
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16040 17746 16068 19178
rect 16132 18630 16160 20402
rect 16224 19904 16252 20402
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 16304 19916 16356 19922
rect 16224 19876 16304 19904
rect 16304 19858 16356 19864
rect 16316 19514 16344 19858
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16408 19394 16436 20334
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16224 19366 16436 19394
rect 16500 19394 16528 19654
rect 16592 19514 16620 19654
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16500 19366 16620 19394
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16132 18329 16160 18566
rect 16118 18320 16174 18329
rect 16118 18255 16174 18264
rect 16224 18222 16252 19366
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16316 18222 16344 19246
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16500 18834 16528 18906
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16212 18216 16264 18222
rect 16132 18176 16212 18204
rect 16132 17785 16160 18176
rect 16212 18158 16264 18164
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16212 17808 16264 17814
rect 16118 17776 16174 17785
rect 16028 17740 16080 17746
rect 16212 17750 16264 17756
rect 16118 17711 16120 17720
rect 16028 17682 16080 17688
rect 16172 17711 16174 17720
rect 16120 17682 16172 17688
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15948 17066 15976 17274
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 16132 13716 16160 17682
rect 16224 17338 16252 17750
rect 16316 17746 16344 18158
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16316 17134 16344 17682
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16316 16794 16344 17070
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16500 15473 16528 18158
rect 16592 17954 16620 19366
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16684 18970 16712 19246
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16776 18766 16804 19654
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16868 18222 16896 19722
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16960 18698 16988 19314
rect 17052 18902 17080 19450
rect 17512 19378 17540 20334
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17222 19272 17278 19281
rect 17222 19207 17224 19216
rect 17276 19207 17278 19216
rect 17316 19236 17368 19242
rect 17224 19178 17276 19184
rect 17316 19178 17368 19184
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17052 18290 17080 18566
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16592 17926 16988 17954
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17066 16804 17614
rect 16960 17134 16988 17926
rect 17144 17882 17172 19110
rect 17224 18828 17276 18834
rect 17328 18816 17356 19178
rect 17276 18788 17356 18816
rect 17224 18770 17276 18776
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16776 15570 16804 17002
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17144 16046 17172 16594
rect 17236 16250 17264 18770
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 16486 15464 16542 15473
rect 16486 15399 16542 15408
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16316 13870 16344 14010
rect 16500 14006 16528 15399
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16578 14512 16634 14521
rect 16578 14447 16634 14456
rect 16592 14414 16620 14447
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16132 13688 16344 13716
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16040 12850 16068 12922
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15856 11558 15884 12038
rect 16132 11676 16160 12038
rect 16224 11830 16252 12242
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16132 11648 16252 11676
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15856 10810 15884 11154
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15752 10124 15804 10130
rect 15856 10112 15884 10746
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15804 10084 15884 10112
rect 15752 10066 15804 10072
rect 15856 9518 15884 10084
rect 15948 9586 15976 10202
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15304 8090 15332 8978
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15658 8120 15714 8129
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15384 8084 15436 8090
rect 15658 8055 15714 8064
rect 15384 8026 15436 8032
rect 15396 7970 15424 8026
rect 15304 7954 15424 7970
rect 15292 7948 15424 7954
rect 15344 7942 15424 7948
rect 15566 7984 15622 7993
rect 15672 7954 15700 8055
rect 15856 7954 15884 8230
rect 15566 7919 15568 7928
rect 15292 7890 15344 7896
rect 15620 7919 15622 7928
rect 15660 7948 15712 7954
rect 15568 7890 15620 7896
rect 15660 7890 15712 7896
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15396 7342 15424 7754
rect 15580 7342 15608 7890
rect 15672 7342 15700 7890
rect 15384 7336 15436 7342
rect 15568 7336 15620 7342
rect 15384 7278 15436 7284
rect 15488 7296 15568 7324
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15304 6730 15332 7210
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4758 14780 5034
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 15488 4690 15516 7296
rect 15568 7278 15620 7284
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15580 6254 15608 6802
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15016 4616 15068 4622
rect 14936 4576 15016 4604
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14936 4486 14964 4576
rect 15016 4558 15068 4564
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14568 4282 14596 4422
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14568 4185 14596 4218
rect 14554 4176 14610 4185
rect 14554 4111 14610 4120
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12096 3836 12404 3845
rect 12096 3834 12102 3836
rect 12158 3834 12182 3836
rect 12238 3834 12262 3836
rect 12318 3834 12342 3836
rect 12398 3834 12404 3836
rect 12158 3782 12160 3834
rect 12340 3782 12342 3834
rect 12096 3780 12102 3782
rect 12158 3780 12182 3782
rect 12238 3780 12262 3782
rect 12318 3780 12342 3782
rect 12398 3780 12404 3782
rect 12096 3771 12404 3780
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 9312 3188 9364 3194
rect 9600 3182 9720 3210
rect 9312 3130 9364 3136
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9232 1494 9260 3062
rect 9588 3052 9640 3058
rect 9508 3012 9588 3040
rect 9508 2446 9536 3012
rect 9588 2994 9640 3000
rect 9692 2938 9720 3182
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 9600 2910 9720 2938
rect 9876 3046 10364 3074
rect 9600 2650 9628 2910
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9876 2582 9904 3046
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2650 10088 2790
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 10152 2378 10180 2926
rect 10244 2582 10272 2926
rect 10336 2854 10364 3046
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10244 2310 10272 2518
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 9416 1766 9444 2246
rect 10244 2106 10272 2246
rect 10428 2106 10456 3130
rect 10520 3126 10548 3470
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10980 2650 11008 3606
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10416 2100 10468 2106
rect 10416 2042 10468 2048
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 9404 1760 9456 1766
rect 9404 1702 9456 1708
rect 9220 1488 9272 1494
rect 9220 1430 9272 1436
rect 8852 1420 8984 1426
rect 8904 1414 8984 1420
rect 9036 1420 9088 1426
rect 8852 1362 8904 1368
rect 9036 1362 9088 1368
rect 8668 1012 8720 1018
rect 8668 954 8720 960
rect 8576 876 8628 882
rect 8576 818 8628 824
rect 9048 814 9076 1362
rect 9784 1018 9812 1838
rect 10612 1834 10640 2382
rect 11072 1902 11100 3334
rect 11436 3292 11744 3301
rect 11436 3290 11442 3292
rect 11498 3290 11522 3292
rect 11578 3290 11602 3292
rect 11658 3290 11682 3292
rect 11738 3290 11744 3292
rect 11498 3238 11500 3290
rect 11680 3238 11682 3290
rect 11436 3236 11442 3238
rect 11498 3236 11522 3238
rect 11578 3236 11602 3238
rect 11658 3236 11682 3238
rect 11738 3236 11744 3238
rect 11436 3227 11744 3236
rect 11808 3126 11836 3402
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11256 2514 11284 2926
rect 11348 2854 11376 2926
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11348 2514 11376 2790
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11808 2310 11836 3062
rect 13188 3058 13216 4014
rect 14936 3602 14964 4422
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12096 2748 12404 2757
rect 12096 2746 12102 2748
rect 12158 2746 12182 2748
rect 12238 2746 12262 2748
rect 12318 2746 12342 2748
rect 12398 2746 12404 2748
rect 12158 2694 12160 2746
rect 12340 2694 12342 2746
rect 12096 2692 12102 2694
rect 12158 2692 12182 2694
rect 12238 2692 12262 2694
rect 12318 2692 12342 2694
rect 12398 2692 12404 2694
rect 12096 2683 12404 2692
rect 12452 2582 12480 2790
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11436 2204 11744 2213
rect 11436 2202 11442 2204
rect 11498 2202 11522 2204
rect 11578 2202 11602 2204
rect 11658 2202 11682 2204
rect 11738 2202 11744 2204
rect 11498 2150 11500 2202
rect 11680 2150 11682 2202
rect 11436 2148 11442 2150
rect 11498 2148 11522 2150
rect 11578 2148 11602 2150
rect 11658 2148 11682 2150
rect 11738 2148 11744 2150
rect 11436 2139 11744 2148
rect 11808 1970 11836 2246
rect 11900 2106 11928 2382
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 12348 2100 12400 2106
rect 12348 2042 12400 2048
rect 11796 1964 11848 1970
rect 11796 1906 11848 1912
rect 11060 1896 11112 1902
rect 11060 1838 11112 1844
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 10612 1562 10640 1770
rect 10600 1556 10652 1562
rect 10600 1498 10652 1504
rect 11808 1290 11836 1906
rect 12360 1902 12388 2042
rect 12544 1970 12572 2994
rect 14108 2990 14136 3062
rect 14384 2990 14412 3334
rect 15028 3058 15056 4014
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 12532 1964 12584 1970
rect 12532 1906 12584 1912
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11992 1426 12020 1702
rect 12096 1660 12404 1669
rect 12096 1658 12102 1660
rect 12158 1658 12182 1660
rect 12238 1658 12262 1660
rect 12318 1658 12342 1660
rect 12398 1658 12404 1660
rect 12158 1606 12160 1658
rect 12340 1606 12342 1658
rect 12096 1604 12102 1606
rect 12158 1604 12182 1606
rect 12238 1604 12262 1606
rect 12318 1604 12342 1606
rect 12398 1604 12404 1606
rect 12096 1595 12404 1604
rect 12636 1494 12664 2926
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13004 2514 13032 2790
rect 13740 2650 13768 2858
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 12820 2088 12848 2450
rect 13636 2304 13688 2310
rect 13740 2258 13768 2586
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 13688 2252 13768 2258
rect 13636 2246 13768 2252
rect 13648 2230 13768 2246
rect 12900 2100 12952 2106
rect 12820 2060 12900 2088
rect 12900 2042 12952 2048
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 13648 1902 13676 2042
rect 13740 1902 13768 2230
rect 13636 1896 13688 1902
rect 13636 1838 13688 1844
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 14004 1896 14056 1902
rect 14004 1838 14056 1844
rect 13360 1760 13412 1766
rect 13360 1702 13412 1708
rect 13728 1760 13780 1766
rect 13728 1702 13780 1708
rect 13372 1494 13400 1702
rect 12624 1488 12676 1494
rect 12624 1430 12676 1436
rect 13360 1488 13412 1494
rect 13360 1430 13412 1436
rect 13740 1426 13768 1702
rect 14016 1562 14044 1838
rect 14004 1556 14056 1562
rect 14004 1498 14056 1504
rect 14108 1426 14136 2314
rect 14844 1970 14872 2858
rect 15028 2650 15056 2994
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 15580 2514 15608 6190
rect 15856 5914 15884 7278
rect 15948 7002 15976 9522
rect 16040 7342 16068 11494
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 10266 16160 10542
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16132 9178 16160 9454
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16224 8378 16252 11648
rect 16132 8350 16252 8378
rect 16132 7954 16160 8350
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 8022 16252 8230
rect 16316 8090 16344 13688
rect 16500 13326 16528 13806
rect 16684 13530 16712 15098
rect 16776 13734 16804 15506
rect 17052 15162 17080 15506
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 16960 14958 16988 15098
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14822 16988 14894
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 13802 17080 14214
rect 17040 13796 17092 13802
rect 17040 13738 17092 13744
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16500 12918 16528 13262
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16592 12374 16620 13126
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16684 11762 16712 12582
rect 17052 11812 17080 13738
rect 17144 13394 17172 15982
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15570 17264 15846
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17222 15056 17278 15065
rect 17222 14991 17278 15000
rect 17236 14482 17264 14991
rect 17328 14521 17356 18090
rect 17788 17134 17816 20538
rect 17880 20466 17908 20810
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17972 20330 18000 21100
rect 18052 21082 18104 21088
rect 18064 20806 18092 21082
rect 18248 21078 18276 21286
rect 18236 21072 18288 21078
rect 18236 21014 18288 21020
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 18156 20058 18184 20334
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 17958 19952 18014 19961
rect 17958 19887 17960 19896
rect 18012 19887 18014 19896
rect 17960 19858 18012 19864
rect 18064 19825 18092 19994
rect 18050 19816 18106 19825
rect 18050 19751 18106 19760
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19310 18092 19654
rect 18340 19310 18368 20946
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 20602 18552 20742
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18708 20534 18736 20878
rect 18800 20602 18828 21626
rect 22204 21486 22232 21791
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19536 21049 19564 21082
rect 19522 21040 19578 21049
rect 19064 21004 19116 21010
rect 19522 20975 19524 20984
rect 19064 20946 19116 20952
rect 19576 20975 19578 20984
rect 19524 20946 19576 20952
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18800 20369 18828 20538
rect 18984 20505 19012 20538
rect 18970 20496 19026 20505
rect 18880 20460 18932 20466
rect 19076 20466 19104 20946
rect 19210 20700 19518 20709
rect 19210 20698 19216 20700
rect 19272 20698 19296 20700
rect 19352 20698 19376 20700
rect 19432 20698 19456 20700
rect 19512 20698 19518 20700
rect 19272 20646 19274 20698
rect 19454 20646 19456 20698
rect 19210 20644 19216 20646
rect 19272 20644 19296 20646
rect 19352 20644 19376 20646
rect 19432 20644 19456 20646
rect 19512 20644 19518 20646
rect 19210 20635 19518 20644
rect 18970 20431 19026 20440
rect 19064 20460 19116 20466
rect 18880 20402 18932 20408
rect 19064 20402 19116 20408
rect 18786 20360 18842 20369
rect 18512 20324 18564 20330
rect 18892 20346 18920 20402
rect 18892 20318 19012 20346
rect 18786 20295 18842 20304
rect 18512 20266 18564 20272
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18156 18970 18184 19246
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18326 18048 18382 18057
rect 18326 17983 18382 17992
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17696 16454 17724 16594
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17512 15638 17540 16390
rect 17696 16182 17724 16390
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17314 14512 17370 14521
rect 17224 14476 17276 14482
rect 17314 14447 17370 14456
rect 17224 14418 17276 14424
rect 17420 14346 17448 14894
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17512 14482 17540 14826
rect 17604 14618 17632 15982
rect 17696 15892 17724 16118
rect 17788 16046 17816 17070
rect 18156 16658 18184 17614
rect 17868 16652 17920 16658
rect 18144 16652 18196 16658
rect 17920 16612 18000 16640
rect 17868 16594 17920 16600
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17776 15904 17828 15910
rect 17696 15864 17776 15892
rect 17776 15846 17828 15852
rect 17788 15706 17816 15846
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17696 14618 17724 14758
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17512 14006 17540 14418
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17604 13870 17632 14554
rect 17788 14414 17816 15642
rect 17776 14408 17828 14414
rect 17696 14356 17776 14362
rect 17696 14350 17828 14356
rect 17696 14334 17816 14350
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17316 13728 17368 13734
rect 17696 13682 17724 14334
rect 17880 14006 17908 15982
rect 17972 15366 18000 16612
rect 18144 16594 18196 16600
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 14822 18000 15302
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17316 13670 17368 13676
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 12306 17172 13126
rect 17328 12782 17356 13670
rect 17512 13654 17724 13682
rect 17512 12918 17540 13654
rect 17788 13190 17816 13874
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17604 12782 17632 13126
rect 17880 13002 17908 13738
rect 17972 13716 18000 14418
rect 18064 14385 18092 15506
rect 18156 15162 18184 15914
rect 18340 15638 18368 17983
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18432 16250 18460 17682
rect 18524 16658 18552 20266
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18708 18834 18736 19722
rect 18800 19514 18828 19858
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18892 19689 18920 19722
rect 18878 19680 18934 19689
rect 18878 19615 18934 19624
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18984 19174 19012 20318
rect 19156 20256 19208 20262
rect 19076 20216 19156 20244
rect 19076 19922 19104 20216
rect 19156 20198 19208 20204
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19352 19922 19380 19994
rect 19628 19922 19656 21422
rect 19870 21244 20178 21253
rect 19870 21242 19876 21244
rect 19932 21242 19956 21244
rect 20012 21242 20036 21244
rect 20092 21242 20116 21244
rect 20172 21242 20178 21244
rect 19932 21190 19934 21242
rect 20114 21190 20116 21242
rect 19870 21188 19876 21190
rect 19932 21188 19956 21190
rect 20012 21188 20036 21190
rect 20092 21188 20116 21190
rect 20172 21188 20178 21190
rect 19706 21176 19762 21185
rect 19870 21179 20178 21188
rect 19706 21111 19762 21120
rect 19720 21010 19748 21111
rect 20640 21010 20668 21422
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 21284 21010 21312 21286
rect 21836 21010 21864 21286
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 19720 20534 19748 20946
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19708 20528 19760 20534
rect 19708 20470 19760 20476
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18602 17640 18658 17649
rect 18602 17575 18658 17584
rect 18616 17202 18644 17575
rect 18708 17542 18736 18022
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18708 17134 18736 17478
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18432 15910 18460 16186
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18144 15020 18196 15026
rect 18248 15008 18276 15506
rect 18326 15464 18382 15473
rect 18326 15399 18328 15408
rect 18380 15399 18382 15408
rect 18328 15370 18380 15376
rect 18196 14980 18276 15008
rect 18144 14962 18196 14968
rect 18248 14482 18276 14980
rect 18524 14550 18552 15574
rect 18708 14958 18736 15846
rect 18800 15638 18828 18770
rect 18984 18358 19012 19110
rect 19076 18834 19104 19858
rect 19352 19825 19380 19858
rect 19338 19816 19394 19825
rect 19338 19751 19394 19760
rect 19210 19612 19518 19621
rect 19210 19610 19216 19612
rect 19272 19610 19296 19612
rect 19352 19610 19376 19612
rect 19432 19610 19456 19612
rect 19512 19610 19518 19612
rect 19272 19558 19274 19610
rect 19454 19558 19456 19610
rect 19210 19556 19216 19558
rect 19272 19556 19296 19558
rect 19352 19556 19376 19558
rect 19432 19556 19456 19558
rect 19512 19556 19518 19558
rect 19210 19547 19518 19556
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 19076 18306 19104 18566
rect 19210 18524 19518 18533
rect 19210 18522 19216 18524
rect 19272 18522 19296 18524
rect 19352 18522 19376 18524
rect 19432 18522 19456 18524
rect 19512 18522 19518 18524
rect 19272 18470 19274 18522
rect 19454 18470 19456 18522
rect 19210 18468 19216 18470
rect 19272 18468 19296 18470
rect 19352 18468 19376 18470
rect 19432 18468 19456 18470
rect 19512 18468 19518 18470
rect 19210 18459 19518 18468
rect 18984 18222 19012 18294
rect 19076 18278 19196 18306
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18892 17660 18920 18158
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 19168 18034 19196 18278
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19246 18048 19302 18057
rect 19076 17746 19104 18022
rect 19168 18006 19246 18034
rect 19246 17983 19302 17992
rect 19260 17746 19288 17983
rect 19352 17882 19380 18158
rect 19628 18154 19656 19858
rect 19812 19786 19840 20810
rect 19996 20602 20024 20878
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 20732 20482 20760 20878
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20916 20505 20944 20538
rect 20548 20454 20760 20482
rect 20902 20496 20958 20505
rect 20548 20398 20576 20454
rect 20902 20431 20958 20440
rect 21008 20398 21036 20742
rect 21560 20602 21588 20878
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21546 20496 21602 20505
rect 21088 20460 21140 20466
rect 21546 20431 21602 20440
rect 21088 20402 21140 20408
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21100 20346 21128 20402
rect 21560 20398 21588 20431
rect 21272 20392 21324 20398
rect 19870 20156 20178 20165
rect 19870 20154 19876 20156
rect 19932 20154 19956 20156
rect 20012 20154 20036 20156
rect 20092 20154 20116 20156
rect 20172 20154 20178 20156
rect 19932 20102 19934 20154
rect 20114 20102 20116 20154
rect 19870 20100 19876 20102
rect 19932 20100 19956 20102
rect 20012 20100 20036 20102
rect 20092 20100 20116 20102
rect 20172 20100 20178 20102
rect 19870 20091 20178 20100
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 20364 19718 20392 20334
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 19720 19378 19748 19654
rect 20456 19446 20484 19790
rect 20548 19514 20576 20334
rect 20732 20058 20760 20334
rect 21100 20318 21220 20346
rect 21272 20334 21324 20340
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20640 19378 20668 19994
rect 21192 19922 21220 20318
rect 21284 20058 21312 20334
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21100 19786 21128 19858
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 19870 19068 20178 19077
rect 19870 19066 19876 19068
rect 19932 19066 19956 19068
rect 20012 19066 20036 19068
rect 20092 19066 20116 19068
rect 20172 19066 20178 19068
rect 19932 19014 19934 19066
rect 20114 19014 20116 19066
rect 19870 19012 19876 19014
rect 19932 19012 19956 19014
rect 20012 19012 20036 19014
rect 20092 19012 20116 19014
rect 20172 19012 20178 19014
rect 19870 19003 20178 19012
rect 20640 18986 20668 19314
rect 21100 19310 21128 19722
rect 21560 19310 21588 20334
rect 21836 19922 21864 20946
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21928 20058 21956 20198
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21824 19916 21876 19922
rect 21824 19858 21876 19864
rect 21652 19514 21680 19858
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 20272 18958 20668 18986
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19444 17814 19472 18022
rect 19536 17814 19564 18090
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 18972 17672 19024 17678
rect 18892 17632 18972 17660
rect 18972 17614 19024 17620
rect 18984 17513 19012 17614
rect 18970 17504 19026 17513
rect 18970 17439 19026 17448
rect 19210 17436 19518 17445
rect 19210 17434 19216 17436
rect 19272 17434 19296 17436
rect 19352 17434 19376 17436
rect 19432 17434 19456 17436
rect 19512 17434 19518 17436
rect 19272 17382 19274 17434
rect 19454 17382 19456 17434
rect 19210 17380 19216 17382
rect 19272 17380 19296 17382
rect 19352 17380 19376 17382
rect 19432 17380 19456 17382
rect 19512 17380 19518 17382
rect 19210 17371 19518 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18696 14952 18748 14958
rect 18788 14952 18840 14958
rect 18696 14894 18748 14900
rect 18786 14920 18788 14929
rect 18892 14940 18920 16934
rect 18984 16658 19012 17070
rect 19076 16794 19104 17070
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19168 16794 19196 17002
rect 19444 16998 19472 17206
rect 19628 17134 19656 17682
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18984 15094 19012 16594
rect 19444 16522 19472 16934
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19536 16658 19564 16730
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19076 16250 19104 16458
rect 19210 16348 19518 16357
rect 19210 16346 19216 16348
rect 19272 16346 19296 16348
rect 19352 16346 19376 16348
rect 19432 16346 19456 16348
rect 19512 16346 19518 16348
rect 19272 16294 19274 16346
rect 19454 16294 19456 16346
rect 19210 16292 19216 16294
rect 19272 16292 19296 16294
rect 19352 16292 19376 16294
rect 19432 16292 19456 16294
rect 19512 16292 19518 16294
rect 19210 16283 19518 16292
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19536 16114 19564 16186
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19628 15994 19656 16934
rect 19720 16726 19748 17682
rect 19812 17134 19840 18090
rect 19870 17980 20178 17989
rect 19870 17978 19876 17980
rect 19932 17978 19956 17980
rect 20012 17978 20036 17980
rect 20092 17978 20116 17980
rect 20172 17978 20178 17980
rect 19932 17926 19934 17978
rect 20114 17926 20116 17978
rect 19870 17924 19876 17926
rect 19932 17924 19956 17926
rect 20012 17924 20036 17926
rect 20092 17924 20116 17926
rect 20172 17924 20178 17926
rect 19870 17915 20178 17924
rect 20272 17354 20300 18958
rect 21100 18902 21128 19246
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20640 18426 20668 18770
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20180 17326 20300 17354
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 20180 16980 20208 17326
rect 20260 17264 20312 17270
rect 20258 17232 20260 17241
rect 20312 17232 20314 17241
rect 20258 17167 20314 17176
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20180 16952 20300 16980
rect 19870 16892 20178 16901
rect 19870 16890 19876 16892
rect 19932 16890 19956 16892
rect 20012 16890 20036 16892
rect 20092 16890 20116 16892
rect 20172 16890 20178 16892
rect 19932 16838 19934 16890
rect 20114 16838 20116 16890
rect 19870 16836 19876 16838
rect 19932 16836 19956 16838
rect 20012 16836 20036 16838
rect 20092 16836 20116 16838
rect 20172 16836 20178 16838
rect 19870 16827 20178 16836
rect 19708 16720 19760 16726
rect 19708 16662 19760 16668
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19720 16114 19748 16458
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19904 16046 19932 16662
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 19892 16040 19944 16046
rect 19628 15966 19748 15994
rect 19616 15632 19668 15638
rect 19616 15574 19668 15580
rect 19210 15260 19518 15269
rect 19210 15258 19216 15260
rect 19272 15258 19296 15260
rect 19352 15258 19376 15260
rect 19432 15258 19456 15260
rect 19512 15258 19518 15260
rect 19272 15206 19274 15258
rect 19454 15206 19456 15258
rect 19210 15204 19216 15206
rect 19272 15204 19296 15206
rect 19352 15204 19376 15206
rect 19432 15204 19456 15206
rect 19512 15204 19518 15206
rect 19210 15195 19518 15204
rect 19628 15162 19656 15574
rect 19720 15570 19748 15966
rect 19812 15988 19892 15994
rect 19812 15982 19944 15988
rect 19812 15966 19932 15982
rect 20088 15978 20116 16594
rect 20272 16538 20300 16952
rect 20364 16658 20392 17002
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20180 16510 20300 16538
rect 20180 16250 20208 16510
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20076 15972 20128 15978
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 19260 15026 19288 15098
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 18972 14952 19024 14958
rect 18840 14920 18842 14929
rect 18892 14912 18972 14940
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18616 14482 18644 14894
rect 18972 14894 19024 14900
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 18786 14855 18842 14864
rect 19156 14816 19208 14822
rect 19352 14804 19380 14894
rect 19208 14776 19380 14804
rect 19156 14758 19208 14764
rect 19720 14618 19748 15302
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 18236 14476 18288 14482
rect 18156 14436 18236 14464
rect 18050 14376 18106 14385
rect 18050 14311 18106 14320
rect 18064 13870 18092 14311
rect 18156 14074 18184 14436
rect 18236 14418 18288 14424
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17972 13688 18092 13716
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17788 12974 17908 13002
rect 17224 12776 17276 12782
rect 17316 12776 17368 12782
rect 17224 12718 17276 12724
rect 17314 12744 17316 12753
rect 17592 12776 17644 12782
rect 17368 12744 17370 12753
rect 17236 12442 17264 12718
rect 17592 12718 17644 12724
rect 17314 12679 17370 12688
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17132 11824 17184 11830
rect 17052 11784 17132 11812
rect 17132 11766 17184 11772
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16408 10266 16436 11154
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9518 16436 10066
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16224 7342 16252 7958
rect 16408 7478 16436 9454
rect 16500 8022 16528 10746
rect 16592 10538 16620 10950
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16776 10198 16804 10474
rect 16868 10198 16896 10950
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16856 10192 16908 10198
rect 16948 10192 17000 10198
rect 16856 10134 16908 10140
rect 16946 10160 16948 10169
rect 17000 10160 17002 10169
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16684 9926 16712 10066
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16592 7886 16620 8366
rect 16776 8090 16804 8366
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16868 8022 16896 10134
rect 17144 10130 17172 11766
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10266 17264 10406
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 16946 10095 17002 10104
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17328 9654 17356 10134
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17420 9042 17448 12378
rect 17604 11014 17632 12718
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17696 10606 17724 11698
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17408 8628 17460 8634
rect 17328 8588 17408 8616
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 16856 8016 16908 8022
rect 16854 7984 16856 7993
rect 16908 7984 16910 7993
rect 17236 7954 17264 8230
rect 16854 7919 16910 7928
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15948 5681 15976 6598
rect 15934 5672 15990 5681
rect 15934 5607 15990 5616
rect 16132 4826 16160 6938
rect 16224 6322 16252 7278
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16500 5642 16528 6258
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16132 4690 16160 4762
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16500 4672 16528 4762
rect 16580 4684 16632 4690
rect 16500 4644 16580 4672
rect 16224 4282 16252 4626
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16132 3738 16160 3946
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16316 3602 16344 4422
rect 16500 3602 16528 4644
rect 16580 4626 16632 4632
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16776 3602 16804 3878
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16960 2854 16988 4422
rect 17144 3670 17172 6734
rect 17328 6186 17356 8588
rect 17408 8570 17460 8576
rect 17512 7410 17540 10406
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17604 9654 17632 10134
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17590 8120 17646 8129
rect 17590 8055 17646 8064
rect 17604 8022 17632 8055
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17788 7954 17816 12974
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17880 11762 17908 12718
rect 17972 12442 18000 13330
rect 18064 12782 18092 13688
rect 18156 13172 18184 14010
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18236 13320 18288 13326
rect 18340 13308 18368 13670
rect 18288 13280 18368 13308
rect 18236 13262 18288 13268
rect 18156 13144 18276 13172
rect 18248 12986 18276 13144
rect 18340 12986 18368 13280
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18144 12912 18196 12918
rect 18142 12880 18144 12889
rect 18196 12880 18198 12889
rect 18142 12815 18198 12824
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18156 11830 18184 12718
rect 18432 12374 18460 13126
rect 18524 12714 18552 14350
rect 18616 14278 18644 14418
rect 19628 14362 19656 14486
rect 19628 14334 19748 14362
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18616 13190 18644 14214
rect 19210 14172 19518 14181
rect 19210 14170 19216 14172
rect 19272 14170 19296 14172
rect 19352 14170 19376 14172
rect 19432 14170 19456 14172
rect 19512 14170 19518 14172
rect 19272 14118 19274 14170
rect 19454 14118 19456 14170
rect 19210 14116 19216 14118
rect 19272 14116 19296 14118
rect 19352 14116 19376 14118
rect 19432 14116 19456 14118
rect 19512 14116 19518 14118
rect 19210 14107 19518 14116
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 13841 19472 13874
rect 19430 13832 19486 13841
rect 19430 13767 19486 13776
rect 19616 13796 19668 13802
rect 19616 13738 19668 13744
rect 19628 13394 19656 13738
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19720 13326 19748 14334
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 19076 12986 19104 13262
rect 19210 13084 19518 13093
rect 19210 13082 19216 13084
rect 19272 13082 19296 13084
rect 19352 13082 19376 13084
rect 19432 13082 19456 13084
rect 19512 13082 19518 13084
rect 19272 13030 19274 13082
rect 19454 13030 19456 13082
rect 19210 13028 19216 13030
rect 19272 13028 19296 13030
rect 19352 13028 19376 13030
rect 19432 13028 19456 13030
rect 19512 13028 19518 13030
rect 19210 13019 19518 13028
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 18420 12368 18472 12374
rect 19628 12345 19656 12378
rect 18420 12310 18472 12316
rect 19614 12336 19670 12345
rect 19064 12300 19116 12306
rect 19614 12271 19670 12280
rect 19708 12300 19760 12306
rect 19064 12242 19116 12248
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 18144 11688 18196 11694
rect 17866 11656 17922 11665
rect 18144 11630 18196 11636
rect 17866 11591 17868 11600
rect 17920 11591 17922 11600
rect 17868 11562 17920 11568
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17972 8430 18000 8842
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17972 7886 18000 8230
rect 18064 7886 18092 9998
rect 18156 9586 18184 11630
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18800 10606 18828 11562
rect 18892 10996 18920 12174
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18984 11694 19012 12106
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 19076 11354 19104 12242
rect 19210 11996 19518 12005
rect 19210 11994 19216 11996
rect 19272 11994 19296 11996
rect 19352 11994 19376 11996
rect 19432 11994 19456 11996
rect 19512 11994 19518 11996
rect 19272 11942 19274 11994
rect 19454 11942 19456 11994
rect 19210 11940 19216 11942
rect 19272 11940 19296 11942
rect 19352 11940 19376 11942
rect 19432 11940 19456 11942
rect 19512 11940 19518 11942
rect 19210 11931 19518 11940
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19524 11348 19576 11354
rect 19628 11336 19656 12271
rect 19708 12242 19760 12248
rect 19720 11642 19748 12242
rect 19812 11898 19840 15966
rect 20076 15914 20128 15920
rect 19870 15804 20178 15813
rect 19870 15802 19876 15804
rect 19932 15802 19956 15804
rect 20012 15802 20036 15804
rect 20092 15802 20116 15804
rect 20172 15802 20178 15804
rect 19932 15750 19934 15802
rect 20114 15750 20116 15802
rect 19870 15748 19876 15750
rect 19932 15748 19956 15750
rect 20012 15748 20036 15750
rect 20092 15748 20116 15750
rect 20172 15748 20178 15750
rect 19870 15739 20178 15748
rect 20272 15638 20300 16390
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19996 15094 20024 15370
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 20364 14872 20392 16118
rect 20456 15570 20484 18022
rect 20640 17814 20668 18090
rect 20628 17808 20680 17814
rect 20628 17750 20680 17756
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20732 17338 20760 17682
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20732 16674 20760 17274
rect 20548 16646 20760 16674
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20272 14844 20392 14872
rect 19870 14716 20178 14725
rect 19870 14714 19876 14716
rect 19932 14714 19956 14716
rect 20012 14714 20036 14716
rect 20092 14714 20116 14716
rect 20172 14714 20178 14716
rect 19932 14662 19934 14714
rect 20114 14662 20116 14714
rect 19870 14660 19876 14662
rect 19932 14660 19956 14662
rect 20012 14660 20036 14662
rect 20092 14660 20116 14662
rect 20172 14660 20178 14662
rect 19870 14651 20178 14660
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19904 14006 19932 14486
rect 20272 14482 20300 14844
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20456 14362 20484 15506
rect 20548 14550 20576 16646
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 14890 20668 16186
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20732 15706 20760 16050
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20732 15162 20760 15642
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 19996 14334 20484 14362
rect 19892 14000 19944 14006
rect 19890 13968 19892 13977
rect 19944 13968 19946 13977
rect 19890 13903 19946 13912
rect 19996 13802 20024 14334
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 20272 13734 20300 13806
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 19870 13628 20178 13637
rect 19870 13626 19876 13628
rect 19932 13626 19956 13628
rect 20012 13626 20036 13628
rect 20092 13626 20116 13628
rect 20172 13626 20178 13628
rect 19932 13574 19934 13626
rect 20114 13574 20116 13626
rect 19870 13572 19876 13574
rect 19932 13572 19956 13574
rect 20012 13572 20036 13574
rect 20092 13572 20116 13574
rect 20172 13572 20178 13574
rect 19870 13563 20178 13572
rect 20456 13530 20484 14214
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20548 13841 20576 13942
rect 20534 13832 20590 13841
rect 20534 13767 20590 13776
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20640 13410 20668 14826
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14482 20760 14758
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20824 13734 20852 17614
rect 20916 17202 20944 18294
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 17202 21128 17682
rect 21284 17610 21312 18566
rect 21376 18222 21404 18566
rect 21836 18222 21864 19858
rect 22112 19854 22140 19994
rect 22204 19922 22232 21082
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22388 18902 22416 21286
rect 23676 20942 23704 21490
rect 23860 21486 23888 21791
rect 24412 21486 24440 21927
rect 26422 21856 26478 21865
rect 26422 21791 26478 21800
rect 26698 21856 26754 21865
rect 26698 21791 26754 21800
rect 25318 21720 25374 21729
rect 25318 21655 25374 21664
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24676 21412 24728 21418
rect 24676 21354 24728 21360
rect 25136 21412 25188 21418
rect 25136 21354 25188 21360
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24044 21078 24072 21286
rect 24032 21072 24084 21078
rect 24032 21014 24084 21020
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23676 20466 23704 20878
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22466 20088 22522 20097
rect 22466 20023 22468 20032
rect 22520 20023 22522 20032
rect 22468 19994 22520 20000
rect 22940 19990 22968 20198
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 23400 19922 23428 20334
rect 24596 20330 24624 21286
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 22376 18896 22428 18902
rect 22376 18838 22428 18844
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22020 18358 22048 18770
rect 23480 18760 23532 18766
rect 24032 18760 24084 18766
rect 23480 18702 23532 18708
rect 24030 18728 24032 18737
rect 24084 18728 24086 18737
rect 22008 18352 22060 18358
rect 22008 18294 22060 18300
rect 23492 18222 23520 18702
rect 24030 18663 24086 18672
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21824 18216 21876 18222
rect 21824 18158 21876 18164
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 21454 17912 21510 17921
rect 21454 17847 21510 17856
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21468 17202 21496 17847
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22008 17536 22060 17542
rect 22204 17513 22232 17682
rect 22008 17478 22060 17484
rect 22190 17504 22246 17513
rect 20904 17196 20956 17202
rect 21088 17196 21140 17202
rect 20904 17138 20956 17144
rect 21008 17156 21088 17184
rect 21008 16794 21036 17156
rect 21088 17138 21140 17144
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21008 15570 21036 16730
rect 21192 16538 21220 17070
rect 21468 16998 21496 17138
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21100 16510 21220 16538
rect 21100 16182 21128 16510
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15609 21312 15846
rect 21376 15706 21404 16594
rect 21824 16176 21876 16182
rect 21824 16118 21876 16124
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 15706 21772 15846
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 21270 15600 21326 15609
rect 20996 15564 21048 15570
rect 21270 15535 21272 15544
rect 20996 15506 21048 15512
rect 21324 15535 21326 15544
rect 21272 15506 21324 15512
rect 21836 15502 21864 16118
rect 22020 16046 22048 17478
rect 22190 17439 22246 17448
rect 22204 16726 22232 17439
rect 22296 16998 22324 18022
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22192 16720 22244 16726
rect 22192 16662 22244 16668
rect 22296 16250 22324 16934
rect 22480 16590 22508 18158
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 22560 17808 22612 17814
rect 22612 17768 22692 17796
rect 22560 17750 22612 17756
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22572 17202 22600 17614
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22664 16794 22692 17768
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22940 16658 22968 17478
rect 23216 16658 23244 17478
rect 23308 17134 23336 18022
rect 23492 17134 23520 18158
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 24136 17882 24164 18090
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23676 16726 23704 17274
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22008 16040 22060 16046
rect 22006 16008 22008 16017
rect 22100 16040 22152 16046
rect 22060 16008 22062 16017
rect 22100 15982 22152 15988
rect 22006 15943 22062 15952
rect 21088 15496 21140 15502
rect 21086 15464 21088 15473
rect 21824 15496 21876 15502
rect 21140 15464 21142 15473
rect 20904 15428 20956 15434
rect 21824 15438 21876 15444
rect 21086 15399 21142 15408
rect 20904 15370 20956 15376
rect 20916 14278 20944 15370
rect 21364 15156 21416 15162
rect 22020 15144 22048 15943
rect 22112 15706 22140 15982
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22296 15638 22324 16186
rect 22572 16046 22600 16458
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22468 15972 22520 15978
rect 22468 15914 22520 15920
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22020 15116 22232 15144
rect 21364 15098 21416 15104
rect 21376 15065 21404 15098
rect 21362 15056 21418 15065
rect 21362 14991 21418 15000
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 21008 13802 21036 14826
rect 21100 14550 21128 14894
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 21100 14006 21128 14486
rect 21376 14482 21404 14894
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21560 14618 21588 14758
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 22112 14482 22140 14894
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 21928 14346 21956 14418
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21284 14074 21312 14214
rect 21744 14113 21772 14214
rect 21730 14104 21786 14113
rect 21272 14068 21324 14074
rect 21730 14039 21786 14048
rect 21272 14010 21324 14016
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 21730 13832 21786 13841
rect 20996 13796 21048 13802
rect 21730 13767 21786 13776
rect 20996 13738 21048 13744
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20272 13382 20668 13410
rect 19870 12540 20178 12549
rect 19870 12538 19876 12540
rect 19932 12538 19956 12540
rect 20012 12538 20036 12540
rect 20092 12538 20116 12540
rect 20172 12538 20178 12540
rect 19932 12486 19934 12538
rect 20114 12486 20116 12538
rect 19870 12484 19876 12486
rect 19932 12484 19956 12486
rect 20012 12484 20036 12486
rect 20092 12484 20116 12486
rect 20172 12484 20178 12486
rect 19870 12475 20178 12484
rect 20272 12434 20300 13382
rect 21744 13326 21772 13767
rect 21928 13394 21956 14282
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 20180 12406 20300 12434
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19904 11762 19932 12174
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19720 11614 19840 11642
rect 20180 11626 20208 12406
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19576 11308 19656 11336
rect 19524 11290 19576 11296
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19338 11112 19394 11121
rect 19444 11098 19472 11154
rect 19720 11098 19748 11494
rect 19812 11336 19840 11614
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 19870 11452 20178 11461
rect 19870 11450 19876 11452
rect 19932 11450 19956 11452
rect 20012 11450 20036 11452
rect 20092 11450 20116 11452
rect 20172 11450 20178 11452
rect 19932 11398 19934 11450
rect 20114 11398 20116 11450
rect 19870 11396 19876 11398
rect 19932 11396 19956 11398
rect 20012 11396 20036 11398
rect 20092 11396 20116 11398
rect 20172 11396 20178 11398
rect 19870 11387 20178 11396
rect 19812 11308 19932 11336
rect 19444 11070 19748 11098
rect 19338 11047 19340 11056
rect 19392 11047 19394 11056
rect 19340 11018 19392 11024
rect 19616 11008 19668 11014
rect 18892 10968 19012 10996
rect 18984 10606 19012 10968
rect 19616 10950 19668 10956
rect 19210 10908 19518 10917
rect 19210 10906 19216 10908
rect 19272 10906 19296 10908
rect 19352 10906 19376 10908
rect 19432 10906 19456 10908
rect 19512 10906 19518 10908
rect 19272 10854 19274 10906
rect 19454 10854 19456 10906
rect 19210 10852 19216 10854
rect 19272 10852 19296 10854
rect 19352 10852 19376 10854
rect 19432 10852 19456 10854
rect 19512 10852 19518 10854
rect 19210 10843 19518 10852
rect 19628 10606 19656 10950
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18340 9518 18368 10474
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18156 8022 18184 8910
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17972 7546 18000 7822
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17592 7540 17644 7546
rect 17960 7540 18012 7546
rect 17644 7500 17908 7528
rect 17592 7482 17644 7488
rect 17880 7426 17908 7500
rect 17960 7482 18012 7488
rect 17500 7404 17552 7410
rect 17420 7364 17500 7392
rect 17420 6322 17448 7364
rect 17880 7398 18000 7426
rect 17500 7346 17552 7352
rect 17972 7206 18000 7398
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 18064 7018 18092 7686
rect 17972 6990 18092 7018
rect 18156 7002 18184 7958
rect 18340 7886 18368 9454
rect 18800 9110 18828 10542
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18432 8022 18460 8910
rect 18524 8090 18552 8978
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8566 18736 8774
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18800 8362 18828 9046
rect 18984 8906 19012 10542
rect 19210 9820 19518 9829
rect 19210 9818 19216 9820
rect 19272 9818 19296 9820
rect 19352 9818 19376 9820
rect 19432 9818 19456 9820
rect 19512 9818 19518 9820
rect 19272 9766 19274 9818
rect 19454 9766 19456 9818
rect 19210 9764 19216 9766
rect 19272 9764 19296 9766
rect 19352 9764 19376 9766
rect 19432 9764 19456 9766
rect 19512 9764 19518 9766
rect 19210 9755 19518 9764
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18892 7546 18920 8774
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18984 8022 19012 8570
rect 19076 8362 19104 9522
rect 19338 9480 19394 9489
rect 19338 9415 19340 9424
rect 19392 9415 19394 9424
rect 19340 9386 19392 9392
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19210 8732 19518 8741
rect 19210 8730 19216 8732
rect 19272 8730 19296 8732
rect 19352 8730 19376 8732
rect 19432 8730 19456 8732
rect 19512 8730 19518 8732
rect 19272 8678 19274 8730
rect 19454 8678 19456 8730
rect 19210 8676 19216 8678
rect 19272 8676 19296 8678
rect 19352 8676 19376 8678
rect 19432 8676 19456 8678
rect 19512 8676 19518 8678
rect 19210 8667 19518 8676
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 19076 7970 19104 8298
rect 19628 8090 19656 9318
rect 19720 8906 19748 11070
rect 19904 10470 19932 11308
rect 19982 11248 20038 11257
rect 20272 11218 20300 12106
rect 20364 11694 20392 12854
rect 20548 12434 20576 13262
rect 20548 12406 20668 12434
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20548 12238 20576 12310
rect 20536 12232 20588 12238
rect 20442 12200 20498 12209
rect 20536 12174 20588 12180
rect 20442 12135 20444 12144
rect 20496 12135 20498 12144
rect 20444 12106 20496 12112
rect 20548 11830 20576 12174
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20548 11354 20576 11766
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20640 11234 20668 12406
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 19982 11183 19984 11192
rect 20036 11183 20038 11192
rect 20076 11212 20128 11218
rect 19984 11154 20036 11160
rect 20076 11154 20128 11160
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20548 11206 20668 11234
rect 19996 11014 20024 11154
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 20088 10520 20116 11154
rect 20180 11082 20208 11154
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20088 10492 20300 10520
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19870 10364 20178 10373
rect 19870 10362 19876 10364
rect 19932 10362 19956 10364
rect 20012 10362 20036 10364
rect 20092 10362 20116 10364
rect 20172 10362 20178 10364
rect 19932 10310 19934 10362
rect 20114 10310 20116 10362
rect 19870 10308 19876 10310
rect 19932 10308 19956 10310
rect 20012 10308 20036 10310
rect 20092 10308 20116 10310
rect 20172 10308 20178 10310
rect 19870 10299 20178 10308
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19996 9722 20024 10066
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 20272 9674 20300 10492
rect 20364 10266 20392 11154
rect 20548 11150 20576 11206
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20548 9722 20576 11086
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20916 10810 20944 11018
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20536 9716 20588 9722
rect 20272 9646 20392 9674
rect 20536 9658 20588 9664
rect 20364 9518 20392 9646
rect 20732 9518 20760 10202
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20824 9586 20852 9930
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20352 9512 20404 9518
rect 20720 9512 20772 9518
rect 20404 9472 20484 9500
rect 20352 9454 20404 9460
rect 19870 9276 20178 9285
rect 19870 9274 19876 9276
rect 19932 9274 19956 9276
rect 20012 9274 20036 9276
rect 20092 9274 20116 9276
rect 20172 9274 20178 9276
rect 19932 9222 19934 9274
rect 20114 9222 20116 9274
rect 19870 9220 19876 9222
rect 19932 9220 19956 9222
rect 20012 9220 20036 9222
rect 20092 9220 20116 9222
rect 20172 9220 20178 9222
rect 19870 9211 20178 9220
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19870 8188 20178 8197
rect 19870 8186 19876 8188
rect 19932 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20178 8188
rect 19932 8134 19934 8186
rect 20114 8134 20116 8186
rect 19870 8132 19876 8134
rect 19932 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20178 8134
rect 19870 8123 20178 8132
rect 20364 8090 20392 8978
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18800 7426 18828 7482
rect 18800 7398 18920 7426
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18144 6996 18196 7002
rect 17972 6798 18000 6990
rect 18144 6938 18196 6944
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 18142 6216 18198 6225
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17500 6180 17552 6186
rect 18142 6151 18144 6160
rect 17500 6122 17552 6128
rect 18196 6151 18198 6160
rect 18144 6122 18196 6128
rect 17236 4622 17264 6122
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17328 4690 17356 4966
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 1970 15332 2246
rect 15580 2106 15608 2450
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 14832 1964 14884 1970
rect 14832 1906 14884 1912
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 15568 1828 15620 1834
rect 15568 1770 15620 1776
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 15488 1562 15516 1702
rect 15580 1562 15608 1770
rect 15476 1556 15528 1562
rect 15476 1498 15528 1504
rect 15568 1556 15620 1562
rect 15568 1498 15620 1504
rect 15764 1426 15792 2246
rect 16316 1426 16344 2246
rect 16500 1494 16528 2246
rect 16580 1964 16632 1970
rect 16580 1906 16632 1912
rect 16488 1488 16540 1494
rect 16488 1430 16540 1436
rect 11980 1420 12032 1426
rect 11980 1362 12032 1368
rect 13728 1420 13780 1426
rect 13728 1362 13780 1368
rect 14096 1420 14148 1426
rect 14096 1362 14148 1368
rect 15752 1420 15804 1426
rect 15752 1362 15804 1368
rect 16304 1420 16356 1426
rect 16304 1362 16356 1368
rect 11796 1284 11848 1290
rect 11796 1226 11848 1232
rect 16592 1222 16620 1906
rect 16960 1902 16988 2790
rect 17236 2650 17264 4558
rect 17420 4146 17448 4694
rect 17512 4690 17540 6122
rect 18248 4826 18276 6870
rect 18708 6866 18736 7278
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18708 6730 18736 6802
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18800 6458 18828 6734
rect 18892 6474 18920 7398
rect 18984 6934 19012 7958
rect 19076 7954 19196 7970
rect 20456 7954 20484 9472
rect 20534 9480 20590 9489
rect 20720 9454 20772 9460
rect 20534 9415 20536 9424
rect 20588 9415 20590 9424
rect 20536 9386 20588 9392
rect 20732 8514 20760 9454
rect 20916 8922 20944 10746
rect 21008 9674 21036 11562
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 21192 10606 21220 11154
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21100 10198 21128 10406
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 21008 9646 21128 9674
rect 20916 8894 21036 8922
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20732 8486 20852 8514
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 19076 7948 19208 7954
rect 19076 7942 19156 7948
rect 19156 7890 19208 7896
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20456 7818 20484 7890
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20640 7750 20668 7890
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 19210 7644 19518 7653
rect 19210 7642 19216 7644
rect 19272 7642 19296 7644
rect 19352 7642 19376 7644
rect 19432 7642 19456 7644
rect 19512 7642 19518 7644
rect 19272 7590 19274 7642
rect 19454 7590 19456 7642
rect 19210 7588 19216 7590
rect 19272 7588 19296 7590
rect 19352 7588 19376 7590
rect 19432 7588 19456 7590
rect 19512 7588 19518 7590
rect 19210 7579 19518 7588
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20732 7324 20760 8298
rect 20824 8022 20852 8486
rect 20916 8430 20944 8774
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 21008 7868 21036 8894
rect 21100 8022 21128 9646
rect 21192 9586 21220 10542
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21192 9042 21220 9522
rect 21284 9042 21312 11834
rect 21468 11694 21496 12038
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 21744 11354 21772 11630
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21180 9036 21232 9042
rect 21180 8978 21232 8984
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21284 8634 21312 8978
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21088 7880 21140 7886
rect 21008 7840 21088 7868
rect 20812 7336 20864 7342
rect 20732 7296 20812 7324
rect 19154 7032 19210 7041
rect 19154 6967 19210 6976
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 19168 6798 19196 6967
rect 19246 6896 19302 6905
rect 19352 6866 19380 7278
rect 19870 7100 20178 7109
rect 19870 7098 19876 7100
rect 19932 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20178 7100
rect 19932 7046 19934 7098
rect 20114 7046 20116 7098
rect 19870 7044 19876 7046
rect 19932 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20178 7046
rect 19870 7035 20178 7044
rect 19246 6831 19248 6840
rect 19300 6831 19302 6840
rect 19340 6860 19392 6866
rect 19248 6802 19300 6808
rect 19340 6802 19392 6808
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19156 6792 19208 6798
rect 18970 6760 19026 6769
rect 19156 6734 19208 6740
rect 18970 6695 19026 6704
rect 18984 6662 19012 6695
rect 19352 6662 19380 6802
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19210 6556 19518 6565
rect 19210 6554 19216 6556
rect 19272 6554 19296 6556
rect 19352 6554 19376 6556
rect 19432 6554 19456 6556
rect 19512 6554 19518 6556
rect 19272 6502 19274 6554
rect 19454 6502 19456 6554
rect 19210 6500 19216 6502
rect 19272 6500 19296 6502
rect 19352 6500 19376 6502
rect 19432 6500 19456 6502
rect 19512 6500 19518 6502
rect 19210 6491 19518 6500
rect 18788 6452 18840 6458
rect 18892 6446 19012 6474
rect 18788 6394 18840 6400
rect 18880 6316 18932 6322
rect 18708 6276 18880 6304
rect 18708 6118 18736 6276
rect 18880 6258 18932 6264
rect 18984 6186 19012 6446
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19154 6352 19210 6361
rect 19536 6322 19564 6394
rect 19154 6287 19210 6296
rect 19524 6316 19576 6322
rect 19168 6254 19196 6287
rect 19524 6258 19576 6264
rect 19628 6254 19656 6802
rect 19982 6352 20038 6361
rect 19982 6287 20038 6296
rect 19996 6254 20024 6287
rect 20364 6254 20392 7278
rect 20732 6934 20760 7296
rect 20812 7278 20864 7284
rect 21008 7274 21036 7840
rect 21088 7822 21140 7828
rect 20996 7268 21048 7274
rect 20996 7210 21048 7216
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19708 6248 19760 6254
rect 19984 6248 20036 6254
rect 19708 6190 19760 6196
rect 19798 6216 19854 6225
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 18696 6112 18748 6118
rect 18984 6089 19012 6122
rect 18696 6054 18748 6060
rect 18970 6080 19026 6089
rect 18970 6015 19026 6024
rect 19076 5953 19104 6122
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19062 5944 19118 5953
rect 18892 5902 19062 5930
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17880 4078 17908 4422
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17972 3942 18000 4626
rect 18156 4282 18184 4626
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18234 4176 18290 4185
rect 18234 4111 18290 4120
rect 18248 4078 18276 4111
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 18248 3738 18276 4014
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18340 2774 18368 5238
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4146 18552 4558
rect 18616 4214 18644 5102
rect 18708 4826 18736 5510
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18432 3670 18460 4014
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18524 3602 18552 4082
rect 18616 4078 18644 4150
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18892 3602 18920 5902
rect 19062 5879 19118 5888
rect 19168 5710 19196 6054
rect 18972 5704 19024 5710
rect 19156 5704 19208 5710
rect 18972 5646 19024 5652
rect 19076 5664 19156 5692
rect 18984 5409 19012 5646
rect 18970 5400 19026 5409
rect 18970 5335 19026 5344
rect 18984 4146 19012 5335
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19076 4010 19104 5664
rect 19156 5646 19208 5652
rect 19260 5642 19288 6122
rect 19616 6112 19668 6118
rect 19338 6080 19394 6089
rect 19616 6054 19668 6060
rect 19338 6015 19394 6024
rect 19352 5642 19380 6015
rect 19628 5846 19656 6054
rect 19720 5914 19748 6190
rect 19984 6190 20036 6196
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 19798 6151 19854 6160
rect 19812 5914 19840 6151
rect 19870 6012 20178 6021
rect 19870 6010 19876 6012
rect 19932 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20178 6012
rect 19932 5958 19934 6010
rect 20114 5958 20116 6010
rect 19870 5956 19876 5958
rect 19932 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20178 5958
rect 19870 5947 20178 5956
rect 20364 5914 20392 6190
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 19616 5840 19668 5846
rect 19720 5817 19748 5850
rect 19616 5782 19668 5788
rect 19706 5808 19762 5817
rect 19706 5743 19762 5752
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19210 5468 19518 5477
rect 19210 5466 19216 5468
rect 19272 5466 19296 5468
rect 19352 5466 19376 5468
rect 19432 5466 19456 5468
rect 19512 5466 19518 5468
rect 19272 5414 19274 5466
rect 19454 5414 19456 5466
rect 19210 5412 19216 5414
rect 19272 5412 19296 5414
rect 19352 5412 19376 5414
rect 19432 5412 19456 5414
rect 19512 5412 19518 5414
rect 19210 5403 19518 5412
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19444 4486 19472 4626
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19210 4380 19518 4389
rect 19210 4378 19216 4380
rect 19272 4378 19296 4380
rect 19352 4378 19376 4380
rect 19432 4378 19456 4380
rect 19512 4378 19518 4380
rect 19272 4326 19274 4378
rect 19454 4326 19456 4378
rect 19210 4324 19216 4326
rect 19272 4324 19296 4326
rect 19352 4324 19376 4326
rect 19432 4324 19456 4326
rect 19512 4324 19518 4326
rect 19210 4315 19518 4324
rect 19628 4282 19656 4762
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 18984 3738 19012 3946
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 19076 3194 19104 3946
rect 19210 3292 19518 3301
rect 19210 3290 19216 3292
rect 19272 3290 19296 3292
rect 19352 3290 19376 3292
rect 19432 3290 19456 3292
rect 19512 3290 19518 3292
rect 19272 3238 19274 3290
rect 19454 3238 19456 3290
rect 19210 3236 19216 3238
rect 19272 3236 19296 3238
rect 19352 3236 19376 3238
rect 19432 3236 19456 3238
rect 19512 3236 19518 3238
rect 19210 3227 19518 3236
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18340 2746 18460 2774
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17236 2514 17264 2586
rect 18432 2514 18460 2746
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 17052 1970 17080 2450
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17144 1970 17172 2314
rect 17040 1964 17092 1970
rect 17040 1906 17092 1912
rect 17132 1964 17184 1970
rect 17132 1906 17184 1912
rect 16948 1896 17000 1902
rect 16948 1838 17000 1844
rect 17236 1562 17264 2450
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17684 1828 17736 1834
rect 17684 1770 17736 1776
rect 17696 1562 17724 1770
rect 17224 1556 17276 1562
rect 17224 1498 17276 1504
rect 17684 1556 17736 1562
rect 17684 1498 17736 1504
rect 17880 1494 17908 2246
rect 17960 1828 18012 1834
rect 17960 1770 18012 1776
rect 17868 1488 17920 1494
rect 17868 1430 17920 1436
rect 17972 1426 18000 1770
rect 17960 1420 18012 1426
rect 17960 1362 18012 1368
rect 16580 1216 16632 1222
rect 16580 1158 16632 1164
rect 11436 1116 11744 1125
rect 11436 1114 11442 1116
rect 11498 1114 11522 1116
rect 11578 1114 11602 1116
rect 11658 1114 11682 1116
rect 11738 1114 11744 1116
rect 11498 1062 11500 1114
rect 11680 1062 11682 1114
rect 11436 1060 11442 1062
rect 11498 1060 11522 1062
rect 11578 1060 11602 1062
rect 11658 1060 11682 1062
rect 11738 1060 11744 1062
rect 11436 1051 11744 1060
rect 9772 1012 9824 1018
rect 9772 954 9824 960
rect 18340 814 18368 2382
rect 18616 2378 18644 2926
rect 19812 2774 19840 5850
rect 20626 5536 20682 5545
rect 20626 5471 20682 5480
rect 19870 4924 20178 4933
rect 19870 4922 19876 4924
rect 19932 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20178 4924
rect 19932 4870 19934 4922
rect 20114 4870 20116 4922
rect 19870 4868 19876 4870
rect 19932 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20178 4870
rect 19870 4859 20178 4868
rect 20640 4690 20668 5471
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 19870 3836 20178 3845
rect 19870 3834 19876 3836
rect 19932 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20178 3836
rect 19932 3782 19934 3834
rect 20114 3782 20116 3834
rect 19870 3780 19876 3782
rect 19932 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20178 3782
rect 19870 3771 20178 3780
rect 20732 3058 20760 6870
rect 21284 6866 21312 8570
rect 21468 7954 21496 9862
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21652 8634 21680 9318
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21836 7954 21864 8842
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21456 7948 21508 7954
rect 21640 7948 21692 7954
rect 21456 7890 21508 7896
rect 21560 7908 21640 7936
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21192 5409 21220 6802
rect 21376 5914 21404 6802
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21178 5400 21234 5409
rect 21178 5335 21234 5344
rect 21376 5273 21404 5510
rect 21362 5264 21418 5273
rect 21468 5234 21496 7890
rect 21560 7206 21588 7908
rect 21640 7890 21692 7896
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 21640 7744 21692 7750
rect 21928 7732 21956 8230
rect 21692 7704 21956 7732
rect 21640 7686 21692 7692
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21362 5199 21418 5208
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21560 5098 21588 5238
rect 21652 5098 21680 7686
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21744 6186 21772 6666
rect 22020 6458 22048 8434
rect 22112 8430 22140 14418
rect 22204 13394 22232 15116
rect 22296 14482 22324 15438
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22296 14249 22324 14418
rect 22282 14240 22338 14249
rect 22282 14175 22338 14184
rect 22388 13870 22416 15846
rect 22480 15706 22508 15914
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22480 14074 22508 14418
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22572 13326 22600 15982
rect 22664 15434 22692 15982
rect 22928 15904 22980 15910
rect 23032 15881 23060 16594
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23400 16250 23428 16458
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23400 15910 23428 16186
rect 23492 15978 23520 16594
rect 23676 16046 23704 16662
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23388 15904 23440 15910
rect 22928 15846 22980 15852
rect 23018 15872 23074 15881
rect 22940 15473 22968 15846
rect 23388 15846 23440 15852
rect 23018 15807 23074 15816
rect 23204 15496 23256 15502
rect 22926 15464 22982 15473
rect 22652 15428 22704 15434
rect 23204 15438 23256 15444
rect 22926 15399 22982 15408
rect 22652 15370 22704 15376
rect 22664 14822 22692 15370
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22756 14550 22784 14962
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22664 13258 22692 14418
rect 22940 13841 22968 15399
rect 23216 15162 23244 15438
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23308 14482 23336 15302
rect 23492 15094 23520 15914
rect 23676 15162 23704 15982
rect 23952 15609 23980 17818
rect 24412 17746 24440 18158
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24400 17740 24452 17746
rect 24400 17682 24452 17688
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24044 16658 24072 17274
rect 24136 16658 24164 17682
rect 24308 17604 24360 17610
rect 24308 17546 24360 17552
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 23938 15600 23994 15609
rect 23938 15535 23940 15544
rect 23992 15535 23994 15544
rect 23940 15506 23992 15512
rect 24044 15366 24072 16594
rect 24136 16182 24164 16594
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 23676 14958 23704 15098
rect 24044 15065 24072 15302
rect 24030 15056 24086 15065
rect 24030 14991 24086 15000
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 23480 14884 23532 14890
rect 23480 14826 23532 14832
rect 23756 14884 23808 14890
rect 23756 14826 23808 14832
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23400 14482 23428 14758
rect 23492 14618 23520 14826
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23584 13870 23612 14758
rect 23768 14074 23796 14826
rect 24044 14618 24072 14894
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24136 14482 24164 16118
rect 24214 15872 24270 15881
rect 24214 15807 24270 15816
rect 24228 14958 24256 15807
rect 24320 15706 24348 17546
rect 24412 17116 24440 17682
rect 24492 17128 24544 17134
rect 24412 17088 24492 17116
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23768 13870 23796 14010
rect 23388 13864 23440 13870
rect 22926 13832 22982 13841
rect 22926 13767 22982 13776
rect 23386 13832 23388 13841
rect 23572 13864 23624 13870
rect 23440 13832 23442 13841
rect 23572 13806 23624 13812
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23386 13767 23442 13776
rect 23860 13530 23888 13806
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 24228 13258 24256 14894
rect 24320 14482 24348 15642
rect 24412 15570 24440 17088
rect 24492 17070 24544 17076
rect 24596 16810 24624 18362
rect 24688 17746 24716 21354
rect 25148 21146 25176 21354
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25332 21010 25360 21655
rect 25502 21584 25558 21593
rect 25502 21519 25558 21528
rect 25516 21010 25544 21519
rect 26436 21486 26464 21791
rect 26712 21486 26740 21791
rect 26984 21788 27292 21797
rect 26984 21786 26990 21788
rect 27046 21786 27070 21788
rect 27126 21786 27150 21788
rect 27206 21786 27230 21788
rect 27286 21786 27292 21788
rect 27046 21734 27048 21786
rect 27228 21734 27230 21786
rect 26984 21732 26990 21734
rect 27046 21732 27070 21734
rect 27126 21732 27150 21734
rect 27206 21732 27230 21734
rect 27286 21732 27292 21734
rect 26984 21723 27292 21732
rect 27356 21486 27384 21927
rect 27724 21486 27752 21927
rect 28262 21856 28318 21865
rect 28262 21791 28318 21800
rect 28276 21486 28304 21791
rect 29276 21684 29328 21690
rect 29276 21626 29328 21632
rect 26424 21480 26476 21486
rect 26424 21422 26476 21428
rect 26700 21480 26752 21486
rect 26700 21422 26752 21428
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 29000 21480 29052 21486
rect 29000 21422 29052 21428
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 27068 21344 27120 21350
rect 27068 21286 27120 21292
rect 27344 21344 27396 21350
rect 27344 21286 27396 21292
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25504 21004 25556 21010
rect 25504 20946 25556 20952
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25332 19922 25360 20742
rect 25884 20602 25912 20878
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25412 20256 25464 20262
rect 25412 20198 25464 20204
rect 25424 19922 25452 20198
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24952 19916 25004 19922
rect 25228 19916 25280 19922
rect 24952 19858 25004 19864
rect 25148 19876 25228 19904
rect 24872 19446 24900 19858
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24872 18970 24900 19382
rect 24964 19174 24992 19858
rect 25148 19417 25176 19876
rect 25228 19858 25280 19864
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25516 19786 25544 19926
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25608 19514 25636 19654
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25134 19408 25190 19417
rect 25884 19378 25912 20538
rect 25976 20398 26004 20742
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25964 19916 26016 19922
rect 26068 19904 26096 21286
rect 27080 21010 27108 21286
rect 27356 21146 27384 21286
rect 27644 21244 27952 21253
rect 27644 21242 27650 21244
rect 27706 21242 27730 21244
rect 27786 21242 27810 21244
rect 27866 21242 27890 21244
rect 27946 21242 27952 21244
rect 27706 21190 27708 21242
rect 27888 21190 27890 21242
rect 27644 21188 27650 21190
rect 27706 21188 27730 21190
rect 27786 21188 27810 21190
rect 27866 21188 27890 21190
rect 27946 21188 27952 21190
rect 27644 21179 27952 21188
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 28356 20800 28408 20806
rect 28356 20742 28408 20748
rect 26984 20700 27292 20709
rect 26984 20698 26990 20700
rect 27046 20698 27070 20700
rect 27126 20698 27150 20700
rect 27206 20698 27230 20700
rect 27286 20698 27292 20700
rect 27046 20646 27048 20698
rect 27228 20646 27230 20698
rect 26984 20644 26990 20646
rect 27046 20644 27070 20646
rect 27126 20644 27150 20646
rect 27206 20644 27230 20646
rect 27286 20644 27292 20646
rect 26984 20635 27292 20644
rect 26608 20256 26660 20262
rect 26608 20198 26660 20204
rect 26700 20256 26752 20262
rect 26700 20198 26752 20204
rect 26514 20088 26570 20097
rect 26332 20052 26384 20058
rect 26620 20058 26648 20198
rect 26514 20023 26570 20032
rect 26608 20052 26660 20058
rect 26332 19994 26384 20000
rect 26016 19876 26096 19904
rect 25964 19858 26016 19864
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 25134 19343 25190 19352
rect 25872 19372 25924 19378
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24872 18154 24900 18702
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24872 17882 24900 18090
rect 24964 18086 24992 18702
rect 25148 18193 25176 19343
rect 25872 19314 25924 19320
rect 25976 19310 26004 19450
rect 25688 19304 25740 19310
rect 25688 19246 25740 19252
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25134 18184 25190 18193
rect 25134 18119 25190 18128
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 24688 17649 24716 17682
rect 24674 17640 24730 17649
rect 24674 17575 24730 17584
rect 24780 17134 24808 17682
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24964 17202 24992 17614
rect 25148 17524 25176 18022
rect 25240 17921 25268 18634
rect 25226 17912 25282 17921
rect 25226 17847 25282 17856
rect 25228 17536 25280 17542
rect 25148 17496 25228 17524
rect 25228 17478 25280 17484
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24950 17096 25006 17105
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24504 16782 24624 16810
rect 24504 16522 24532 16782
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24320 14385 24348 14418
rect 24306 14376 24362 14385
rect 24306 14311 24362 14320
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24320 13462 24348 13738
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 24596 13394 24624 15438
rect 24688 14958 24716 16934
rect 24780 16522 24808 17070
rect 24950 17031 25006 17040
rect 25136 17060 25188 17066
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24872 16726 24900 16934
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 24780 16046 24808 16458
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24964 15978 24992 17031
rect 25136 17002 25188 17008
rect 25148 16250 25176 17002
rect 25240 16998 25268 17478
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25240 16658 25268 16934
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25240 16114 25268 16594
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24872 14482 24900 15302
rect 24964 14958 24992 15506
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 25228 14952 25280 14958
rect 25332 14929 25360 19110
rect 25700 18970 25728 19246
rect 26056 19236 26108 19242
rect 26056 19178 26108 19184
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 25412 17808 25464 17814
rect 25412 17750 25464 17756
rect 25424 15978 25452 17750
rect 25516 16250 25544 18158
rect 25608 17338 25636 18158
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25608 17066 25636 17274
rect 25596 17060 25648 17066
rect 25596 17002 25648 17008
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25412 15972 25464 15978
rect 25412 15914 25464 15920
rect 25424 15881 25452 15914
rect 25700 15892 25728 18906
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25792 18222 25820 18362
rect 25884 18329 25912 18702
rect 25870 18320 25926 18329
rect 25870 18255 25926 18264
rect 25884 18222 25912 18255
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 25792 17785 25820 18158
rect 25778 17776 25834 17785
rect 25778 17711 25834 17720
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25792 17338 25820 17614
rect 25780 17332 25832 17338
rect 25780 17274 25832 17280
rect 25884 17134 25912 18158
rect 26068 17898 26096 19178
rect 26252 19174 26280 19654
rect 26344 19378 26372 19994
rect 26528 19922 26556 20023
rect 26608 19994 26660 20000
rect 26712 19990 26740 20198
rect 27644 20156 27952 20165
rect 27644 20154 27650 20156
rect 27706 20154 27730 20156
rect 27786 20154 27810 20156
rect 27866 20154 27890 20156
rect 27946 20154 27952 20156
rect 27706 20102 27708 20154
rect 27888 20102 27890 20154
rect 27644 20100 27650 20102
rect 27706 20100 27730 20102
rect 27786 20100 27810 20102
rect 27866 20100 27890 20102
rect 27946 20100 27952 20102
rect 27644 20091 27952 20100
rect 28368 20058 28396 20742
rect 29012 20398 29040 21422
rect 29184 21072 29236 21078
rect 29184 21014 29236 21020
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 26700 19984 26752 19990
rect 26700 19926 26752 19932
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 27988 19916 28040 19922
rect 27988 19858 28040 19864
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 26804 19514 26832 19858
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 26984 19612 27292 19621
rect 26984 19610 26990 19612
rect 27046 19610 27070 19612
rect 27126 19610 27150 19612
rect 27206 19610 27230 19612
rect 27286 19610 27292 19612
rect 27046 19558 27048 19610
rect 27228 19558 27230 19610
rect 26984 19556 26990 19558
rect 27046 19556 27070 19558
rect 27126 19556 27150 19558
rect 27206 19556 27230 19558
rect 27286 19556 27292 19558
rect 26984 19547 27292 19556
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 27724 19446 27752 19654
rect 27712 19440 27764 19446
rect 27712 19382 27764 19388
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 25976 17870 26096 17898
rect 25976 17202 26004 17870
rect 26056 17808 26108 17814
rect 26056 17750 26108 17756
rect 26068 17513 26096 17750
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 26054 17504 26110 17513
rect 26054 17439 26110 17448
rect 25964 17196 26016 17202
rect 25964 17138 26016 17144
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25792 16046 25820 16730
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 25780 16040 25832 16046
rect 25780 15982 25832 15988
rect 25410 15872 25466 15881
rect 25700 15864 25820 15892
rect 25410 15807 25466 15816
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25228 14894 25280 14900
rect 25318 14920 25374 14929
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24780 14362 24808 14418
rect 24780 14334 24900 14362
rect 24872 14278 24900 14334
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24964 13841 24992 14894
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24950 13832 25006 13841
rect 24950 13767 25006 13776
rect 25056 13462 25084 14758
rect 25240 14113 25268 14894
rect 25318 14855 25374 14864
rect 25320 14816 25372 14822
rect 25320 14758 25372 14764
rect 25332 14550 25360 14758
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25226 14104 25282 14113
rect 25148 14048 25226 14056
rect 25148 14028 25228 14048
rect 25044 13456 25096 13462
rect 25044 13398 25096 13404
rect 25148 13394 25176 14028
rect 25280 14039 25282 14048
rect 25228 14010 25280 14016
rect 25424 13938 25452 15098
rect 25516 15026 25544 15098
rect 25596 15088 25648 15094
rect 25596 15030 25648 15036
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25504 14816 25556 14822
rect 25504 14758 25556 14764
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25228 13388 25280 13394
rect 25332 13376 25360 13670
rect 25424 13462 25452 13874
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25516 13394 25544 14758
rect 25608 13394 25636 15030
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25700 13870 25728 14010
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25280 13348 25360 13376
rect 25504 13388 25556 13394
rect 25228 13330 25280 13336
rect 25504 13330 25556 13336
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 22192 12368 22244 12374
rect 22244 12328 22324 12356
rect 22192 12310 22244 12316
rect 22192 12232 22244 12238
rect 22296 12209 22324 12328
rect 22192 12174 22244 12180
rect 22282 12200 22338 12209
rect 22204 11626 22232 12174
rect 22282 12135 22338 12144
rect 22192 11620 22244 11626
rect 22192 11562 22244 11568
rect 22388 10810 22416 13194
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22848 12434 22876 13126
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 22756 12406 22968 12434
rect 22468 12368 22520 12374
rect 22560 12368 22612 12374
rect 22468 12310 22520 12316
rect 22558 12336 22560 12345
rect 22612 12336 22614 12345
rect 22480 11880 22508 12310
rect 22558 12271 22614 12280
rect 22756 12238 22784 12406
rect 22744 12232 22796 12238
rect 22836 12232 22888 12238
rect 22744 12174 22796 12180
rect 22834 12200 22836 12209
rect 22888 12200 22890 12209
rect 22834 12135 22890 12144
rect 22652 11892 22704 11898
rect 22480 11852 22652 11880
rect 22652 11834 22704 11840
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22480 11082 22508 11630
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22204 9110 22232 9522
rect 22388 9178 22416 10066
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22192 9104 22244 9110
rect 22190 9072 22192 9081
rect 22244 9072 22246 9081
rect 22190 9007 22246 9016
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22296 8673 22324 8910
rect 22282 8664 22338 8673
rect 22388 8634 22416 8978
rect 22282 8599 22338 8608
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22112 7206 22140 7754
rect 22296 7750 22324 7958
rect 22480 7750 22508 11018
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 22572 9518 22600 9862
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22572 8430 22600 9114
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22572 8090 22600 8366
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22664 7954 22692 11834
rect 22742 10160 22798 10169
rect 22848 10146 22876 12135
rect 22798 10118 22876 10146
rect 22742 10095 22798 10104
rect 22756 9178 22784 10095
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22848 9042 22876 9114
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22756 8430 22784 8570
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22848 8294 22876 8978
rect 22940 8974 22968 12406
rect 23110 12336 23166 12345
rect 23020 12300 23072 12306
rect 23110 12271 23112 12280
rect 23020 12242 23072 12248
rect 23164 12271 23166 12280
rect 24032 12300 24084 12306
rect 23112 12242 23164 12248
rect 24032 12242 24084 12248
rect 23032 11694 23060 12242
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23020 11688 23072 11694
rect 23308 11642 23336 11698
rect 23400 11694 23428 12038
rect 23020 11630 23072 11636
rect 23124 11614 23336 11642
rect 23388 11688 23440 11694
rect 23388 11630 23440 11636
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23124 11558 23152 11614
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23216 11286 23244 11494
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23308 10062 23336 11614
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23492 11218 23520 11494
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22926 8664 22982 8673
rect 22926 8599 22928 8608
rect 22980 8599 22982 8608
rect 22928 8570 22980 8576
rect 23400 8430 23428 9862
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23584 9042 23612 9386
rect 23676 9081 23704 11630
rect 24044 11218 24072 12242
rect 24872 11762 24900 12650
rect 25688 12368 25740 12374
rect 25688 12310 25740 12316
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24032 11212 24084 11218
rect 24032 11154 24084 11160
rect 24044 10606 24072 11154
rect 24872 10674 24900 11698
rect 25056 11694 25084 12038
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 25332 11354 25360 12242
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25516 11218 25544 12242
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25608 11218 25636 11494
rect 25504 11212 25556 11218
rect 25424 11172 25504 11200
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 23952 10130 23980 10406
rect 23940 10124 23992 10130
rect 23940 10066 23992 10072
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23662 9072 23718 9081
rect 23572 9036 23624 9042
rect 23662 9007 23718 9016
rect 23572 8978 23624 8984
rect 23676 8430 23704 9007
rect 23768 8906 23796 9318
rect 24044 9042 24072 10406
rect 24228 9489 24256 10610
rect 24492 9512 24544 9518
rect 24214 9480 24270 9489
rect 24492 9454 24544 9460
rect 24214 9415 24270 9424
rect 24308 9444 24360 9450
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 23756 8900 23808 8906
rect 23756 8842 23808 8848
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 24136 8362 24164 8978
rect 24228 8974 24256 9415
rect 24308 9386 24360 9392
rect 24320 8974 24348 9386
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24504 8838 24532 9454
rect 24872 9042 24900 10610
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25148 9926 25176 10542
rect 25424 10130 25452 11172
rect 25504 11154 25556 11160
rect 25596 11212 25648 11218
rect 25700 11200 25728 12310
rect 25792 12102 25820 15864
rect 25870 15056 25926 15065
rect 25870 14991 25926 15000
rect 25884 14958 25912 14991
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25976 14822 26004 16390
rect 26068 16046 26096 17439
rect 26160 17338 26188 17682
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26160 16182 26188 17138
rect 26148 16176 26200 16182
rect 26148 16118 26200 16124
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25964 14816 26016 14822
rect 25964 14758 26016 14764
rect 25872 13728 25924 13734
rect 25872 13670 25924 13676
rect 25884 13462 25912 13670
rect 26068 13462 26096 14894
rect 26160 14414 26188 16118
rect 26252 15910 26280 17682
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26252 15094 26280 15846
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26160 14278 26188 14350
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 13938 26188 14214
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 25872 13456 25924 13462
rect 25872 13398 25924 13404
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 26344 12782 26372 19314
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 26436 18834 26464 19110
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26528 18426 26556 18770
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 26896 18222 26924 19110
rect 26984 18524 27292 18533
rect 26984 18522 26990 18524
rect 27046 18522 27070 18524
rect 27126 18522 27150 18524
rect 27206 18522 27230 18524
rect 27286 18522 27292 18524
rect 27046 18470 27048 18522
rect 27228 18470 27230 18522
rect 26984 18468 26990 18470
rect 27046 18468 27070 18470
rect 27126 18468 27150 18470
rect 27206 18468 27230 18470
rect 27286 18468 27292 18470
rect 26984 18459 27292 18468
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 26712 17882 26740 18158
rect 26792 18148 26844 18154
rect 26792 18090 26844 18096
rect 26700 17876 26752 17882
rect 26700 17818 26752 17824
rect 26804 17202 26832 18090
rect 26896 17649 26924 18158
rect 27356 17814 27384 19246
rect 27644 19068 27952 19077
rect 27644 19066 27650 19068
rect 27706 19066 27730 19068
rect 27786 19066 27810 19068
rect 27866 19066 27890 19068
rect 27946 19066 27952 19068
rect 27706 19014 27708 19066
rect 27888 19014 27890 19066
rect 27644 19012 27650 19014
rect 27706 19012 27730 19014
rect 27786 19012 27810 19014
rect 27866 19012 27890 19014
rect 27946 19012 27952 19014
rect 27644 19003 27952 19012
rect 28000 18970 28028 19858
rect 28184 19514 28212 19858
rect 28172 19508 28224 19514
rect 28172 19450 28224 19456
rect 28446 19408 28502 19417
rect 28446 19343 28502 19352
rect 28460 19242 28488 19343
rect 29012 19310 29040 20334
rect 29092 20256 29144 20262
rect 29092 20198 29144 20204
rect 29104 19990 29132 20198
rect 29092 19984 29144 19990
rect 29092 19926 29144 19932
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 28448 19236 28500 19242
rect 28448 19178 28500 19184
rect 29000 19168 29052 19174
rect 29104 19122 29132 19654
rect 29196 19446 29224 21014
rect 29288 20398 29316 21626
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 29460 20868 29512 20874
rect 29460 20810 29512 20816
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29380 19922 29408 20742
rect 29472 19922 29500 20810
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 29734 19952 29790 19961
rect 29368 19916 29420 19922
rect 29368 19858 29420 19864
rect 29460 19916 29512 19922
rect 29734 19887 29736 19896
rect 29460 19858 29512 19864
rect 29788 19887 29790 19896
rect 29736 19858 29788 19864
rect 29184 19440 29236 19446
rect 30024 19417 30052 20742
rect 30116 19990 30144 21286
rect 30392 21146 30420 21286
rect 30380 21140 30432 21146
rect 30380 21082 30432 21088
rect 30104 19984 30156 19990
rect 30104 19926 30156 19932
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 29184 19382 29236 19388
rect 30010 19408 30066 19417
rect 30010 19343 30066 19352
rect 29552 19236 29604 19242
rect 29552 19178 29604 19184
rect 29052 19116 29132 19122
rect 29000 19110 29132 19116
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29460 19168 29512 19174
rect 29460 19110 29512 19116
rect 29012 19094 29132 19110
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27724 18154 27752 18566
rect 27986 18320 28042 18329
rect 28092 18290 28120 18906
rect 28724 18896 28776 18902
rect 28724 18838 28776 18844
rect 28736 18630 28764 18838
rect 29380 18834 29408 19110
rect 29472 18902 29500 19110
rect 29564 18970 29592 19178
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29460 18896 29512 18902
rect 29460 18838 29512 18844
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 29368 18828 29420 18834
rect 29368 18770 29420 18776
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 28368 18358 28396 18566
rect 28356 18352 28408 18358
rect 28356 18294 28408 18300
rect 27986 18255 28042 18264
rect 28080 18284 28132 18290
rect 28000 18222 28028 18255
rect 28080 18226 28132 18232
rect 28448 18284 28500 18290
rect 28448 18226 28500 18232
rect 27988 18216 28040 18222
rect 27988 18158 28040 18164
rect 28172 18216 28224 18222
rect 28224 18176 28304 18204
rect 28172 18158 28224 18164
rect 27712 18148 27764 18154
rect 27712 18090 27764 18096
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 27644 17980 27952 17989
rect 27644 17978 27650 17980
rect 27706 17978 27730 17980
rect 27786 17978 27810 17980
rect 27866 17978 27890 17980
rect 27946 17978 27952 17980
rect 27706 17926 27708 17978
rect 27888 17926 27890 17978
rect 27644 17924 27650 17926
rect 27706 17924 27730 17926
rect 27786 17924 27810 17926
rect 27866 17924 27890 17926
rect 27946 17924 27952 17926
rect 27644 17915 27952 17924
rect 28092 17814 28120 18022
rect 27344 17808 27396 17814
rect 27344 17750 27396 17756
rect 28080 17808 28132 17814
rect 28080 17750 28132 17756
rect 26882 17640 26938 17649
rect 26882 17575 26938 17584
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 26712 15978 26740 16594
rect 26700 15972 26752 15978
rect 26700 15914 26752 15920
rect 26712 15570 26740 15914
rect 26700 15564 26752 15570
rect 26700 15506 26752 15512
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26422 14240 26478 14249
rect 26422 14175 26478 14184
rect 26436 13394 26464 14175
rect 26516 13796 26568 13802
rect 26516 13738 26568 13744
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 26148 12776 26200 12782
rect 26332 12776 26384 12782
rect 26148 12718 26200 12724
rect 26252 12736 26332 12764
rect 25976 12442 26004 12718
rect 25964 12436 26016 12442
rect 25964 12378 26016 12384
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 25884 12170 25912 12242
rect 25976 12186 26004 12242
rect 26160 12238 26188 12718
rect 26252 12481 26280 12736
rect 26332 12718 26384 12724
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26238 12472 26294 12481
rect 26238 12407 26294 12416
rect 26344 12306 26372 12582
rect 26332 12300 26384 12306
rect 26332 12242 26384 12248
rect 26148 12232 26200 12238
rect 25872 12164 25924 12170
rect 25976 12158 26096 12186
rect 26148 12174 26200 12180
rect 25872 12106 25924 12112
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25780 11212 25832 11218
rect 25700 11172 25780 11200
rect 25596 11154 25648 11160
rect 25780 11154 25832 11160
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25516 10198 25544 10406
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23032 7954 23060 8230
rect 23584 8022 23612 8230
rect 24320 8090 24348 8434
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 23572 8016 23624 8022
rect 23572 7958 23624 7964
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22388 7478 22416 7686
rect 22572 7546 22600 7890
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22480 7002 22508 7346
rect 22664 7002 22692 7890
rect 23296 7744 23348 7750
rect 23348 7704 23428 7732
rect 23296 7686 23348 7692
rect 22836 7268 22888 7274
rect 22836 7210 22888 7216
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22284 6656 22336 6662
rect 22336 6604 22416 6610
rect 22284 6598 22416 6604
rect 22296 6582 22416 6598
rect 22282 6488 22338 6497
rect 22008 6452 22060 6458
rect 22282 6423 22338 6432
rect 22008 6394 22060 6400
rect 22296 6390 22324 6423
rect 22284 6384 22336 6390
rect 22284 6326 22336 6332
rect 22008 6248 22060 6254
rect 22006 6216 22008 6225
rect 22192 6248 22244 6254
rect 22060 6216 22062 6225
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21824 6180 21876 6186
rect 22192 6190 22244 6196
rect 22006 6151 22062 6160
rect 21824 6122 21876 6128
rect 21744 5953 21772 6122
rect 21730 5944 21786 5953
rect 21730 5879 21786 5888
rect 21836 5710 21864 6122
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21744 5370 21772 5510
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 22020 5302 22048 5714
rect 22008 5296 22060 5302
rect 22008 5238 22060 5244
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 22020 4486 22048 5238
rect 22112 5166 22140 5714
rect 22204 5574 22232 6190
rect 22388 6186 22416 6582
rect 22480 6254 22508 6938
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6662 22600 6734
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22376 6180 22428 6186
rect 22376 6122 22428 6128
rect 22388 5846 22416 6122
rect 22284 5840 22336 5846
rect 22284 5782 22336 5788
rect 22376 5840 22428 5846
rect 22376 5782 22428 5788
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22296 5370 22324 5782
rect 22376 5704 22428 5710
rect 22572 5692 22600 6394
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22428 5664 22600 5692
rect 22376 5646 22428 5652
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22112 4078 22140 4558
rect 22388 4554 22416 5034
rect 22664 5001 22692 5714
rect 22756 5574 22784 6802
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 22756 5273 22784 5510
rect 22742 5264 22798 5273
rect 22742 5199 22798 5208
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22650 4992 22706 5001
rect 22650 4927 22706 4936
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 22192 4208 22244 4214
rect 22192 4150 22244 4156
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21560 3534 21588 3674
rect 22112 3670 22140 4014
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 19720 2746 19840 2774
rect 19870 2748 20178 2757
rect 19870 2746 19876 2748
rect 19932 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20178 2748
rect 19720 2650 19748 2746
rect 19932 2694 19934 2746
rect 20114 2694 20116 2746
rect 19870 2692 19876 2694
rect 19932 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20178 2694
rect 19870 2683 20178 2692
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 18616 2106 18644 2314
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 18800 1834 18828 2518
rect 18788 1828 18840 1834
rect 18788 1770 18840 1776
rect 18696 1352 18748 1358
rect 18696 1294 18748 1300
rect 18708 1018 18736 1294
rect 18696 1012 18748 1018
rect 18696 954 18748 960
rect 18800 898 18828 1770
rect 18892 1018 18920 2586
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 18880 1012 18932 1018
rect 18880 954 18932 960
rect 18800 870 18920 898
rect 8392 808 8444 814
rect 8392 750 8444 756
rect 9036 808 9088 814
rect 9036 750 9088 756
rect 18328 808 18380 814
rect 18328 750 18380 756
rect 18892 746 18920 870
rect 18984 746 19012 2450
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19076 1562 19104 2246
rect 19210 2204 19518 2213
rect 19210 2202 19216 2204
rect 19272 2202 19296 2204
rect 19352 2202 19376 2204
rect 19432 2202 19456 2204
rect 19512 2202 19518 2204
rect 19272 2150 19274 2202
rect 19454 2150 19456 2202
rect 19210 2148 19216 2150
rect 19272 2148 19296 2150
rect 19352 2148 19376 2150
rect 19432 2148 19456 2150
rect 19512 2148 19518 2150
rect 19210 2139 19518 2148
rect 19720 1902 19748 2586
rect 20364 2446 20392 2926
rect 20916 2514 20944 3334
rect 22112 3194 22140 3606
rect 22204 3602 22232 4150
rect 22664 3738 22692 4626
rect 22756 4146 22784 5102
rect 22848 4690 22876 7210
rect 23020 6996 23072 7002
rect 23020 6938 23072 6944
rect 23032 6390 23060 6938
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23308 6730 23336 6802
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23110 6488 23166 6497
rect 23110 6423 23166 6432
rect 23124 6390 23152 6423
rect 23020 6384 23072 6390
rect 23020 6326 23072 6332
rect 23112 6384 23164 6390
rect 23112 6326 23164 6332
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 22940 5710 22968 5850
rect 23020 5840 23072 5846
rect 23020 5782 23072 5788
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22928 5568 22980 5574
rect 23032 5556 23060 5782
rect 22980 5528 23060 5556
rect 22928 5510 22980 5516
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 22940 4826 22968 5102
rect 23032 4826 23060 5528
rect 23124 5302 23152 6054
rect 23216 5778 23244 6054
rect 23294 5944 23350 5953
rect 23294 5879 23350 5888
rect 23204 5772 23256 5778
rect 23204 5714 23256 5720
rect 23308 5574 23336 5879
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23216 5234 23244 5510
rect 23204 5228 23256 5234
rect 23400 5216 23428 7704
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 23480 6860 23532 6866
rect 23532 6820 23612 6848
rect 23480 6802 23532 6808
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23492 5914 23520 6598
rect 23584 6458 23612 6820
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23664 6724 23716 6730
rect 23664 6666 23716 6672
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23676 5846 23704 6666
rect 23768 6390 23796 6734
rect 23860 6662 23888 7142
rect 24044 6866 24072 7346
rect 24320 6934 24348 8026
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24308 6928 24360 6934
rect 24308 6870 24360 6876
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23756 6384 23808 6390
rect 23756 6326 23808 6332
rect 23860 6118 23888 6598
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 23204 5170 23256 5176
rect 23308 5188 23428 5216
rect 23202 5128 23258 5137
rect 23202 5063 23204 5072
rect 23256 5063 23258 5072
rect 23204 5034 23256 5040
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23308 4706 23336 5188
rect 23388 5092 23440 5098
rect 23388 5034 23440 5040
rect 23400 4826 23428 5034
rect 23492 5030 23520 5578
rect 23584 5030 23612 5714
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23662 5400 23718 5409
rect 23768 5370 23796 5510
rect 23662 5335 23718 5344
rect 23756 5364 23808 5370
rect 23676 5302 23704 5335
rect 23756 5306 23808 5312
rect 23664 5296 23716 5302
rect 23664 5238 23716 5244
rect 23860 5166 23888 6054
rect 23952 5930 23980 6802
rect 23952 5902 24164 5930
rect 23940 5840 23992 5846
rect 23940 5782 23992 5788
rect 23952 5642 23980 5782
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23572 5024 23624 5030
rect 23952 5001 23980 5102
rect 23572 4966 23624 4972
rect 23938 4992 23994 5001
rect 23938 4927 23994 4936
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 24044 4758 24072 5714
rect 24136 5166 24164 5902
rect 24412 5778 24440 7142
rect 24596 6866 24624 8842
rect 24872 8498 24900 8978
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 25148 8362 25176 9862
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25136 8356 25188 8362
rect 25136 8298 25188 8304
rect 25148 7342 25176 8298
rect 25240 7410 25268 9318
rect 25332 9110 25360 9318
rect 25320 9104 25372 9110
rect 25320 9046 25372 9052
rect 25608 8616 25636 11154
rect 25792 10538 25820 11154
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25884 10169 25912 11290
rect 25976 11218 26004 12038
rect 26068 11830 26096 12158
rect 26344 12084 26372 12242
rect 26252 12056 26372 12084
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 26252 11218 26280 12056
rect 26436 11218 26464 12582
rect 26528 12374 26556 13738
rect 26620 13394 26648 14758
rect 26712 14618 26740 14894
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26804 14346 26832 15506
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26712 13462 26740 14214
rect 26804 14006 26832 14282
rect 26792 14000 26844 14006
rect 26792 13942 26844 13948
rect 26896 13954 26924 17575
rect 26984 17436 27292 17445
rect 26984 17434 26990 17436
rect 27046 17434 27070 17436
rect 27126 17434 27150 17436
rect 27206 17434 27230 17436
rect 27286 17434 27292 17436
rect 27046 17382 27048 17434
rect 27228 17382 27230 17434
rect 26984 17380 26990 17382
rect 27046 17380 27070 17382
rect 27126 17380 27150 17382
rect 27206 17380 27230 17382
rect 27286 17380 27292 17382
rect 26984 17371 27292 17380
rect 27356 17134 27384 17750
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28080 17604 28132 17610
rect 28080 17546 28132 17552
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27434 17368 27490 17377
rect 27434 17303 27490 17312
rect 27344 17128 27396 17134
rect 27344 17070 27396 17076
rect 27344 16516 27396 16522
rect 27344 16458 27396 16464
rect 26984 16348 27292 16357
rect 26984 16346 26990 16348
rect 27046 16346 27070 16348
rect 27126 16346 27150 16348
rect 27206 16346 27230 16348
rect 27286 16346 27292 16348
rect 27046 16294 27048 16346
rect 27228 16294 27230 16346
rect 26984 16292 26990 16294
rect 27046 16292 27070 16294
rect 27126 16292 27150 16294
rect 27206 16292 27230 16294
rect 27286 16292 27292 16294
rect 26984 16283 27292 16292
rect 27356 15978 27384 16458
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 26984 15260 27292 15269
rect 26984 15258 26990 15260
rect 27046 15258 27070 15260
rect 27126 15258 27150 15260
rect 27206 15258 27230 15260
rect 27286 15258 27292 15260
rect 27046 15206 27048 15258
rect 27228 15206 27230 15258
rect 26984 15204 26990 15206
rect 27046 15204 27070 15206
rect 27126 15204 27150 15206
rect 27206 15204 27230 15206
rect 27286 15204 27292 15206
rect 26984 15195 27292 15204
rect 26984 14172 27292 14181
rect 26984 14170 26990 14172
rect 27046 14170 27070 14172
rect 27126 14170 27150 14172
rect 27206 14170 27230 14172
rect 27286 14170 27292 14172
rect 27046 14118 27048 14170
rect 27228 14118 27230 14170
rect 26984 14116 26990 14118
rect 27046 14116 27070 14118
rect 27126 14116 27150 14118
rect 27206 14116 27230 14118
rect 27286 14116 27292 14118
rect 26984 14107 27292 14116
rect 27356 13977 27384 15914
rect 27448 15638 27476 17303
rect 27632 17134 27660 17478
rect 27986 17232 28042 17241
rect 27986 17167 27988 17176
rect 28040 17167 28042 17176
rect 27988 17138 28040 17144
rect 27620 17128 27672 17134
rect 27896 17128 27948 17134
rect 27620 17070 27672 17076
rect 27894 17096 27896 17105
rect 27948 17096 27950 17105
rect 27894 17031 27950 17040
rect 27988 17060 28040 17066
rect 27988 17002 28040 17008
rect 27644 16892 27952 16901
rect 27644 16890 27650 16892
rect 27706 16890 27730 16892
rect 27786 16890 27810 16892
rect 27866 16890 27890 16892
rect 27946 16890 27952 16892
rect 27706 16838 27708 16890
rect 27888 16838 27890 16890
rect 27644 16836 27650 16838
rect 27706 16836 27730 16838
rect 27786 16836 27810 16838
rect 27866 16836 27890 16838
rect 27946 16836 27952 16838
rect 27644 16827 27952 16836
rect 28000 16674 28028 17002
rect 27908 16658 28028 16674
rect 27896 16652 28028 16658
rect 27948 16646 28028 16652
rect 27896 16594 27948 16600
rect 27620 16516 27672 16522
rect 27620 16458 27672 16464
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27436 15632 27488 15638
rect 27436 15574 27488 15580
rect 27448 14958 27476 15574
rect 27540 15570 27568 16390
rect 27632 16046 27660 16458
rect 27620 16040 27672 16046
rect 27804 16040 27856 16046
rect 27620 15982 27672 15988
rect 27802 16008 27804 16017
rect 27856 16008 27858 16017
rect 27802 15943 27858 15952
rect 28092 15910 28120 17546
rect 28184 17066 28212 17614
rect 28172 17060 28224 17066
rect 28172 17002 28224 17008
rect 28184 16114 28212 17002
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 27644 15804 27952 15813
rect 27644 15802 27650 15804
rect 27706 15802 27730 15804
rect 27786 15802 27810 15804
rect 27866 15802 27890 15804
rect 27946 15802 27952 15804
rect 27706 15750 27708 15802
rect 27888 15750 27890 15802
rect 27644 15748 27650 15750
rect 27706 15748 27730 15750
rect 27786 15748 27810 15750
rect 27866 15748 27890 15750
rect 27946 15748 27952 15750
rect 27644 15739 27952 15748
rect 27804 15632 27856 15638
rect 27804 15574 27856 15580
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27816 15434 27844 15574
rect 28184 15570 28212 15846
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27908 15162 27936 15506
rect 27988 15428 28040 15434
rect 27988 15370 28040 15376
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27448 14414 27476 14758
rect 27540 14618 27568 14894
rect 27644 14716 27952 14725
rect 27644 14714 27650 14716
rect 27706 14714 27730 14716
rect 27786 14714 27810 14716
rect 27866 14714 27890 14716
rect 27946 14714 27952 14716
rect 27706 14662 27708 14714
rect 27888 14662 27890 14714
rect 27644 14660 27650 14662
rect 27706 14660 27730 14662
rect 27786 14660 27810 14662
rect 27866 14660 27890 14662
rect 27946 14660 27952 14662
rect 27644 14651 27952 14660
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 28000 14482 28028 15370
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 27988 14476 28040 14482
rect 28040 14436 28120 14464
rect 27988 14418 28040 14424
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27342 13968 27398 13977
rect 26896 13926 27292 13954
rect 26884 13864 26936 13870
rect 26976 13864 27028 13870
rect 26884 13806 26936 13812
rect 26974 13832 26976 13841
rect 27028 13832 27030 13841
rect 26896 13546 26924 13806
rect 27264 13818 27292 13926
rect 27342 13903 27398 13912
rect 27264 13790 27384 13818
rect 27448 13802 27476 14350
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 27620 13932 27672 13938
rect 27620 13874 27672 13880
rect 27632 13818 27660 13874
rect 26974 13767 27030 13776
rect 26896 13518 27016 13546
rect 26988 13462 27016 13518
rect 26700 13456 26752 13462
rect 26700 13398 26752 13404
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 26984 13084 27292 13093
rect 26984 13082 26990 13084
rect 27046 13082 27070 13084
rect 27126 13082 27150 13084
rect 27206 13082 27230 13084
rect 27286 13082 27292 13084
rect 27046 13030 27048 13082
rect 27228 13030 27230 13082
rect 26984 13028 26990 13030
rect 27046 13028 27070 13030
rect 27126 13028 27150 13030
rect 27206 13028 27230 13030
rect 27286 13028 27292 13030
rect 26984 13019 27292 13028
rect 26700 12912 26752 12918
rect 26700 12854 26752 12860
rect 26516 12368 26568 12374
rect 26516 12310 26568 12316
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 26514 12200 26570 12209
rect 26514 12135 26570 12144
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 26056 11212 26108 11218
rect 26056 11154 26108 11160
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26068 11121 26096 11154
rect 26054 11112 26110 11121
rect 26054 11047 26110 11056
rect 26528 10742 26556 12135
rect 26620 11354 26648 12242
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 26712 11286 26740 12854
rect 27356 12434 27384 13790
rect 27436 13796 27488 13802
rect 27436 13738 27488 13744
rect 27540 13790 27660 13818
rect 27540 13410 27568 13790
rect 27644 13628 27952 13637
rect 27644 13626 27650 13628
rect 27706 13626 27730 13628
rect 27786 13626 27810 13628
rect 27866 13626 27890 13628
rect 27946 13626 27952 13628
rect 27706 13574 27708 13626
rect 27888 13574 27890 13626
rect 27644 13572 27650 13574
rect 27706 13572 27730 13574
rect 27786 13572 27810 13574
rect 27866 13572 27890 13574
rect 27946 13572 27952 13574
rect 27644 13563 27952 13572
rect 28000 13462 28028 14214
rect 27988 13456 28040 13462
rect 27540 13394 27660 13410
rect 27988 13398 28040 13404
rect 27540 13388 27672 13394
rect 27540 13382 27620 13388
rect 27620 13330 27672 13336
rect 28092 12782 28120 14436
rect 28184 14074 28212 14962
rect 28276 14958 28304 18176
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 28368 17338 28396 17682
rect 28460 17610 28488 18226
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28552 17882 28580 18158
rect 28540 17876 28592 17882
rect 28540 17818 28592 17824
rect 28630 17776 28686 17785
rect 28540 17740 28592 17746
rect 28736 17762 28764 18566
rect 28828 18426 28856 18770
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28906 18320 28962 18329
rect 29012 18306 29040 18770
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 28962 18278 29040 18306
rect 28906 18255 28962 18264
rect 29000 18148 29052 18154
rect 29000 18090 29052 18096
rect 29092 18148 29144 18154
rect 29092 18090 29144 18096
rect 29012 17882 29040 18090
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29104 17762 29132 18090
rect 28736 17746 29132 17762
rect 28630 17711 28632 17720
rect 28540 17682 28592 17688
rect 28684 17711 28686 17720
rect 28724 17740 29132 17746
rect 28632 17682 28684 17688
rect 28776 17734 29132 17740
rect 28724 17682 28776 17688
rect 28448 17604 28500 17610
rect 28448 17546 28500 17552
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28460 17184 28488 17546
rect 28552 17377 28580 17682
rect 28724 17604 28776 17610
rect 28724 17546 28776 17552
rect 28538 17368 28594 17377
rect 28538 17303 28594 17312
rect 28630 17232 28686 17241
rect 28460 17156 28580 17184
rect 28630 17167 28686 17176
rect 28448 17060 28500 17066
rect 28448 17002 28500 17008
rect 28460 16590 28488 17002
rect 28552 16998 28580 17156
rect 28644 17066 28672 17167
rect 28632 17060 28684 17066
rect 28632 17002 28684 17008
rect 28540 16992 28592 16998
rect 28540 16934 28592 16940
rect 28736 16658 28764 17546
rect 29196 17218 29224 18702
rect 29368 18352 29420 18358
rect 29368 18294 29420 18300
rect 29276 18080 29328 18086
rect 29276 18022 29328 18028
rect 29288 17814 29316 18022
rect 29276 17808 29328 17814
rect 29276 17750 29328 17756
rect 29380 17626 29408 18294
rect 29472 17882 29500 18838
rect 30208 18834 30236 19654
rect 29644 18828 29696 18834
rect 29644 18770 29696 18776
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 29656 18426 29684 18770
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29460 17876 29512 17882
rect 29460 17818 29512 17824
rect 29458 17776 29514 17785
rect 29458 17711 29514 17720
rect 28816 17196 28868 17202
rect 28816 17138 28868 17144
rect 29104 17190 29224 17218
rect 29288 17598 29408 17626
rect 28828 16658 28856 17138
rect 29104 17134 29132 17190
rect 29288 17134 29316 17598
rect 28908 17128 28960 17134
rect 28908 17070 28960 17076
rect 29092 17128 29144 17134
rect 29092 17070 29144 17076
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29276 17128 29328 17134
rect 29276 17070 29328 17076
rect 28920 16658 28948 17070
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 28816 16652 28868 16658
rect 28816 16594 28868 16600
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28644 16046 28672 16594
rect 28632 16040 28684 16046
rect 28632 15982 28684 15988
rect 28540 15972 28592 15978
rect 28540 15914 28592 15920
rect 28448 15360 28500 15366
rect 28448 15302 28500 15308
rect 28264 14952 28316 14958
rect 28264 14894 28316 14900
rect 28460 14482 28488 15302
rect 28552 14958 28580 15914
rect 28736 15162 28764 16594
rect 28828 16266 28856 16594
rect 29104 16538 29132 17070
rect 29012 16510 29132 16538
rect 29012 16454 29040 16510
rect 29000 16448 29052 16454
rect 29000 16390 29052 16396
rect 28828 16238 29132 16266
rect 29196 16250 29224 17070
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28920 15706 28948 15846
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 28540 14952 28592 14958
rect 28540 14894 28592 14900
rect 28816 14952 28868 14958
rect 28816 14894 28868 14900
rect 28828 14657 28856 14894
rect 28920 14822 28948 15642
rect 29012 15094 29040 15642
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 29104 14958 29132 16238
rect 29184 16244 29236 16250
rect 29184 16186 29236 16192
rect 29288 15994 29316 17070
rect 29196 15966 29316 15994
rect 29196 15366 29224 15966
rect 29276 15564 29328 15570
rect 29276 15506 29328 15512
rect 29184 15360 29236 15366
rect 29184 15302 29236 15308
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 28908 14816 28960 14822
rect 28908 14758 28960 14764
rect 28814 14648 28870 14657
rect 28920 14618 28948 14758
rect 28814 14583 28870 14592
rect 28908 14612 28960 14618
rect 28448 14476 28500 14482
rect 28448 14418 28500 14424
rect 28828 14385 28856 14583
rect 28908 14554 28960 14560
rect 29184 14476 29236 14482
rect 29184 14418 29236 14424
rect 28814 14376 28870 14385
rect 28814 14311 28870 14320
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 28172 14068 28224 14074
rect 28172 14010 28224 14016
rect 28170 13832 28226 13841
rect 28170 13767 28226 13776
rect 28184 13462 28212 13767
rect 28172 13456 28224 13462
rect 28172 13398 28224 13404
rect 28644 13394 28672 14214
rect 28724 13728 28776 13734
rect 28724 13670 28776 13676
rect 28736 13530 28764 13670
rect 28724 13524 28776 13530
rect 28724 13466 28776 13472
rect 28632 13388 28684 13394
rect 28632 13330 28684 13336
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 27644 12540 27952 12549
rect 27644 12538 27650 12540
rect 27706 12538 27730 12540
rect 27786 12538 27810 12540
rect 27866 12538 27890 12540
rect 27946 12538 27952 12540
rect 27706 12486 27708 12538
rect 27888 12486 27890 12538
rect 27644 12484 27650 12486
rect 27706 12484 27730 12486
rect 27786 12484 27810 12486
rect 27866 12484 27890 12486
rect 27946 12484 27952 12486
rect 27644 12475 27952 12484
rect 28632 12436 28684 12442
rect 27356 12406 27476 12434
rect 27448 12306 27476 12406
rect 28632 12378 28684 12384
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 26792 12164 26844 12170
rect 26792 12106 26844 12112
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26804 10810 26832 12106
rect 26896 11898 26924 12242
rect 26984 11996 27292 12005
rect 26984 11994 26990 11996
rect 27046 11994 27070 11996
rect 27126 11994 27150 11996
rect 27206 11994 27230 11996
rect 27286 11994 27292 11996
rect 27046 11942 27048 11994
rect 27228 11942 27230 11994
rect 26984 11940 26990 11942
rect 27046 11940 27070 11942
rect 27126 11940 27150 11942
rect 27206 11940 27230 11942
rect 27286 11940 27292 11942
rect 26984 11931 27292 11940
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 26984 10908 27292 10917
rect 26984 10906 26990 10908
rect 27046 10906 27070 10908
rect 27126 10906 27150 10908
rect 27206 10906 27230 10908
rect 27286 10906 27292 10908
rect 27046 10854 27048 10906
rect 27228 10854 27230 10906
rect 26984 10852 26990 10854
rect 27046 10852 27070 10854
rect 27126 10852 27150 10854
rect 27206 10852 27230 10854
rect 27286 10852 27292 10854
rect 26984 10843 27292 10852
rect 26792 10804 26844 10810
rect 26792 10746 26844 10752
rect 26516 10736 26568 10742
rect 26516 10678 26568 10684
rect 27160 10736 27212 10742
rect 27160 10678 27212 10684
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 26240 10532 26292 10538
rect 26240 10474 26292 10480
rect 26252 10198 26280 10474
rect 26240 10192 26292 10198
rect 25870 10160 25926 10169
rect 26240 10134 26292 10140
rect 25870 10095 25926 10104
rect 25780 9988 25832 9994
rect 25780 9930 25832 9936
rect 25792 9722 25820 9930
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 26068 9450 26096 9862
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 26056 9444 26108 9450
rect 26056 9386 26108 9392
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25688 8628 25740 8634
rect 25608 8588 25688 8616
rect 25688 8570 25740 8576
rect 25792 8430 25820 8774
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24492 6724 24544 6730
rect 24492 6666 24544 6672
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24228 5370 24256 5646
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24320 5234 24348 5510
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24124 5160 24176 5166
rect 24124 5102 24176 5108
rect 23756 4752 23808 4758
rect 23308 4690 23704 4706
rect 23756 4694 23808 4700
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 23296 4684 23716 4690
rect 23348 4678 23664 4684
rect 23296 4626 23348 4632
rect 23664 4626 23716 4632
rect 22848 4146 22876 4626
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23492 4282 23520 4558
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 23768 4078 23796 4694
rect 24044 4554 24072 4694
rect 24228 4690 24256 5170
rect 24216 4684 24268 4690
rect 24216 4626 24268 4632
rect 24320 4622 24348 5170
rect 24504 4758 24532 6666
rect 24596 5545 24624 6802
rect 24688 5778 24716 7278
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 6866 25268 7142
rect 25884 7002 25912 7482
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24582 5536 24638 5545
rect 24582 5471 24638 5480
rect 24688 5386 24716 5714
rect 24596 5358 24716 5386
rect 24768 5364 24820 5370
rect 24596 5137 24624 5358
rect 24768 5306 24820 5312
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24582 5128 24638 5137
rect 24582 5063 24638 5072
rect 24492 4752 24544 4758
rect 24492 4694 24544 4700
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24032 4548 24084 4554
rect 24032 4490 24084 4496
rect 24504 4282 24532 4694
rect 24492 4276 24544 4282
rect 24492 4218 24544 4224
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22388 3618 22416 3674
rect 22388 3602 22876 3618
rect 22192 3596 22244 3602
rect 22388 3596 22888 3602
rect 22388 3590 22836 3596
rect 22192 3538 22244 3544
rect 22836 3538 22888 3544
rect 22204 3482 22232 3538
rect 24596 3534 24624 5063
rect 24688 4486 24716 5238
rect 24780 4486 24808 5306
rect 24964 4554 24992 5782
rect 25056 5681 25084 6802
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25516 6361 25544 6598
rect 25502 6352 25558 6361
rect 25502 6287 25558 6296
rect 25136 6180 25188 6186
rect 25136 6122 25188 6128
rect 25042 5672 25098 5681
rect 25042 5607 25098 5616
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 25056 4758 25084 5102
rect 25044 4752 25096 4758
rect 25044 4694 25096 4700
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24780 4146 24808 4422
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 25148 3738 25176 6122
rect 25410 5808 25466 5817
rect 25410 5743 25412 5752
rect 25464 5743 25466 5752
rect 25412 5714 25464 5720
rect 25884 5302 25912 6938
rect 25872 5296 25924 5302
rect 25872 5238 25924 5244
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25240 4690 25268 5102
rect 25884 5098 25912 5238
rect 25872 5092 25924 5098
rect 25872 5034 25924 5040
rect 25976 4690 26004 8570
rect 26252 8430 26280 9658
rect 26344 8838 26372 10542
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26712 10130 26740 10406
rect 26700 10124 26752 10130
rect 26700 10066 26752 10072
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26804 9722 26832 10066
rect 27172 10062 27200 10678
rect 27356 10606 27384 11290
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27448 10266 27476 12242
rect 27712 12164 27764 12170
rect 27712 12106 27764 12112
rect 27724 11694 27752 12106
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 27712 11688 27764 11694
rect 27712 11630 27764 11636
rect 27644 11452 27952 11461
rect 27644 11450 27650 11452
rect 27706 11450 27730 11452
rect 27786 11450 27810 11452
rect 27866 11450 27890 11452
rect 27946 11450 27952 11452
rect 27706 11398 27708 11450
rect 27888 11398 27890 11450
rect 27644 11396 27650 11398
rect 27706 11396 27730 11398
rect 27786 11396 27810 11398
rect 27866 11396 27890 11398
rect 27946 11396 27952 11398
rect 27644 11387 27952 11396
rect 28000 10470 28028 11834
rect 28644 11218 28672 12378
rect 29012 12374 29040 14214
rect 29104 13394 29132 14214
rect 29196 13530 29224 14418
rect 29288 14414 29316 15506
rect 29472 15026 29500 17711
rect 29564 17678 29592 18226
rect 31036 18222 31064 18566
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 31024 18216 31076 18222
rect 31024 18158 31076 18164
rect 30288 17876 30340 17882
rect 30288 17818 30340 17824
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 29552 17672 29604 17678
rect 29552 17614 29604 17620
rect 30024 17626 30052 17682
rect 29564 17270 29592 17614
rect 30024 17598 30144 17626
rect 29552 17264 29604 17270
rect 29552 17206 29604 17212
rect 29564 16114 29592 17206
rect 30012 17060 30064 17066
rect 30012 17002 30064 17008
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29460 15020 29512 15026
rect 29460 14962 29512 14968
rect 29748 14958 29776 16730
rect 30024 16726 30052 17002
rect 30116 16794 30144 17598
rect 30208 17202 30236 17682
rect 30300 17270 30328 17818
rect 30392 17338 30420 18158
rect 30472 17536 30524 17542
rect 30472 17478 30524 17484
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30380 17332 30432 17338
rect 30380 17274 30432 17280
rect 30484 17270 30512 17478
rect 30288 17264 30340 17270
rect 30288 17206 30340 17212
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30196 16992 30248 16998
rect 30196 16934 30248 16940
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30012 16720 30064 16726
rect 30012 16662 30064 16668
rect 30024 16046 30052 16662
rect 30012 16040 30064 16046
rect 30012 15982 30064 15988
rect 29828 15904 29880 15910
rect 29828 15846 29880 15852
rect 29840 15570 29868 15846
rect 30116 15586 30144 16730
rect 30208 16726 30236 16934
rect 30196 16720 30248 16726
rect 30196 16662 30248 16668
rect 30300 16454 30328 17206
rect 30576 17134 30604 17478
rect 30564 17128 30616 17134
rect 30564 17070 30616 17076
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 30760 16794 30788 17070
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 30748 16788 30800 16794
rect 30748 16730 30800 16736
rect 31220 16658 31248 16934
rect 31208 16652 31260 16658
rect 31208 16594 31260 16600
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30300 15706 30328 16390
rect 30288 15700 30340 15706
rect 30288 15642 30340 15648
rect 29828 15564 29880 15570
rect 30116 15558 30328 15586
rect 29828 15506 29880 15512
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29564 14618 29592 14894
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 30104 14816 30156 14822
rect 30104 14758 30156 14764
rect 29552 14612 29604 14618
rect 29552 14554 29604 14560
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29288 13938 29316 14350
rect 29368 14000 29420 14006
rect 29564 13988 29592 14554
rect 29656 14550 29684 14758
rect 29644 14544 29696 14550
rect 29644 14486 29696 14492
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 29840 14074 29868 14418
rect 29828 14068 29880 14074
rect 29828 14010 29880 14016
rect 29564 13960 29684 13988
rect 29368 13942 29420 13948
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29380 13734 29408 13942
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 29564 12782 29592 13126
rect 29656 12986 29684 13960
rect 30116 13870 30144 14758
rect 30300 14482 30328 15558
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30760 14958 30788 15506
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 30562 14648 30618 14657
rect 30562 14583 30618 14592
rect 30576 14482 30604 14583
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30484 14074 30512 14418
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 30760 13734 30788 14894
rect 30930 14512 30986 14521
rect 30930 14447 30932 14456
rect 30984 14447 30986 14456
rect 30932 14418 30984 14424
rect 30748 13728 30800 13734
rect 30748 13670 30800 13676
rect 30760 13326 30788 13670
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 29000 12368 29052 12374
rect 29000 12310 29052 12316
rect 29104 12306 29132 12582
rect 30760 12442 30788 13262
rect 31036 12986 31064 13262
rect 31024 12980 31076 12986
rect 31024 12922 31076 12928
rect 30748 12436 30800 12442
rect 30748 12378 30800 12384
rect 29092 12300 29144 12306
rect 29092 12242 29144 12248
rect 29000 11688 29052 11694
rect 29000 11630 29052 11636
rect 30288 11688 30340 11694
rect 30288 11630 30340 11636
rect 30840 11688 30892 11694
rect 30840 11630 30892 11636
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28816 11212 28868 11218
rect 28816 11154 28868 11160
rect 28080 10736 28132 10742
rect 28080 10678 28132 10684
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 27644 10364 27952 10373
rect 27644 10362 27650 10364
rect 27706 10362 27730 10364
rect 27786 10362 27810 10364
rect 27866 10362 27890 10364
rect 27946 10362 27952 10364
rect 27706 10310 27708 10362
rect 27888 10310 27890 10362
rect 27644 10308 27650 10310
rect 27706 10308 27730 10310
rect 27786 10308 27810 10310
rect 27866 10308 27890 10310
rect 27946 10308 27952 10310
rect 27644 10299 27952 10308
rect 28000 10266 28028 10406
rect 27436 10260 27488 10266
rect 27436 10202 27488 10208
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 27434 10160 27490 10169
rect 28092 10146 28120 10678
rect 28644 10470 28672 11154
rect 28828 10810 28856 11154
rect 28816 10804 28868 10810
rect 28816 10746 28868 10752
rect 28632 10464 28684 10470
rect 28632 10406 28684 10412
rect 28644 10198 28672 10406
rect 27434 10095 27436 10104
rect 27488 10095 27490 10104
rect 27528 10124 27580 10130
rect 27436 10066 27488 10072
rect 27528 10066 27580 10072
rect 28000 10118 28120 10146
rect 28632 10192 28684 10198
rect 28632 10134 28684 10140
rect 28908 10192 28960 10198
rect 28908 10134 28960 10140
rect 28448 10124 28500 10130
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 26884 9988 26936 9994
rect 26884 9930 26936 9936
rect 26896 9722 26924 9930
rect 26984 9820 27292 9829
rect 26984 9818 26990 9820
rect 27046 9818 27070 9820
rect 27126 9818 27150 9820
rect 27206 9818 27230 9820
rect 27286 9818 27292 9820
rect 27046 9766 27048 9818
rect 27228 9766 27230 9818
rect 26984 9764 26990 9766
rect 27046 9764 27070 9766
rect 27126 9764 27150 9766
rect 27206 9764 27230 9766
rect 27286 9764 27292 9766
rect 26984 9755 27292 9764
rect 26792 9716 26844 9722
rect 26792 9658 26844 9664
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 26516 9104 26568 9110
rect 26516 9046 26568 9052
rect 26528 8906 26556 9046
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26252 6798 26280 8366
rect 26344 7478 26372 8774
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26436 8022 26464 8366
rect 26424 8016 26476 8022
rect 26424 7958 26476 7964
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 26344 6934 26372 7414
rect 26528 7002 26556 8842
rect 26984 8732 27292 8741
rect 26984 8730 26990 8732
rect 27046 8730 27070 8732
rect 27126 8730 27150 8732
rect 27206 8730 27230 8732
rect 27286 8730 27292 8732
rect 27046 8678 27048 8730
rect 27228 8678 27230 8730
rect 26984 8676 26990 8678
rect 27046 8676 27070 8678
rect 27126 8676 27150 8678
rect 27206 8676 27230 8678
rect 27286 8676 27292 8678
rect 26984 8667 27292 8676
rect 27448 8022 27476 9114
rect 27540 9110 27568 10066
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 27908 9518 27936 9862
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 28000 9466 28028 10118
rect 28448 10066 28500 10072
rect 28080 9988 28132 9994
rect 28080 9930 28132 9936
rect 28092 9674 28120 9930
rect 28092 9646 28212 9674
rect 28184 9518 28212 9646
rect 28172 9512 28224 9518
rect 28000 9438 28120 9466
rect 28172 9454 28224 9460
rect 27988 9376 28040 9382
rect 27988 9318 28040 9324
rect 27644 9276 27952 9285
rect 27644 9274 27650 9276
rect 27706 9274 27730 9276
rect 27786 9274 27810 9276
rect 27866 9274 27890 9276
rect 27946 9274 27952 9276
rect 27706 9222 27708 9274
rect 27888 9222 27890 9274
rect 27644 9220 27650 9222
rect 27706 9220 27730 9222
rect 27786 9220 27810 9222
rect 27866 9220 27890 9222
rect 27946 9220 27952 9222
rect 27644 9211 27952 9220
rect 28000 9110 28028 9318
rect 27528 9104 27580 9110
rect 27528 9046 27580 9052
rect 27988 9104 28040 9110
rect 27988 9046 28040 9052
rect 27644 8188 27952 8197
rect 27644 8186 27650 8188
rect 27706 8186 27730 8188
rect 27786 8186 27810 8188
rect 27866 8186 27890 8188
rect 27946 8186 27952 8188
rect 27706 8134 27708 8186
rect 27888 8134 27890 8186
rect 27644 8132 27650 8134
rect 27706 8132 27730 8134
rect 27786 8132 27810 8134
rect 27866 8132 27890 8134
rect 27946 8132 27952 8134
rect 27644 8123 27952 8132
rect 27436 8016 27488 8022
rect 27436 7958 27488 7964
rect 27896 7948 27948 7954
rect 27896 7890 27948 7896
rect 26984 7644 27292 7653
rect 26984 7642 26990 7644
rect 27046 7642 27070 7644
rect 27126 7642 27150 7644
rect 27206 7642 27230 7644
rect 27286 7642 27292 7644
rect 27046 7590 27048 7642
rect 27228 7590 27230 7642
rect 26984 7588 26990 7590
rect 27046 7588 27070 7590
rect 27126 7588 27150 7590
rect 27206 7588 27230 7590
rect 27286 7588 27292 7590
rect 26984 7579 27292 7588
rect 27908 7342 27936 7890
rect 28092 7886 28120 9438
rect 28264 8560 28316 8566
rect 28264 8502 28316 8508
rect 28276 8022 28304 8502
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28264 8016 28316 8022
rect 28264 7958 28316 7964
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28368 7342 28396 8434
rect 28460 8362 28488 10066
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28552 8634 28580 9454
rect 28644 8974 28672 10134
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28736 9042 28764 9318
rect 28724 9036 28776 9042
rect 28724 8978 28776 8984
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28644 8498 28672 8910
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28828 8430 28856 9658
rect 28920 8566 28948 10134
rect 29012 9722 29040 11630
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 29920 11552 29972 11558
rect 29920 11494 29972 11500
rect 29380 11218 29408 11494
rect 29932 11354 29960 11494
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 29368 11212 29420 11218
rect 29368 11154 29420 11160
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 29104 10606 29132 11086
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 29196 10674 29224 11018
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 30300 10606 30328 11630
rect 30852 11082 30880 11630
rect 30840 11076 30892 11082
rect 30840 11018 30892 11024
rect 30852 10742 30880 11018
rect 30840 10736 30892 10742
rect 30840 10678 30892 10684
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 30104 10600 30156 10606
rect 30104 10542 30156 10548
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 29288 10062 29316 10542
rect 30012 10464 30064 10470
rect 30012 10406 30064 10412
rect 30024 10198 30052 10406
rect 30116 10266 30144 10542
rect 30748 10464 30800 10470
rect 30748 10406 30800 10412
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 29920 10192 29972 10198
rect 29920 10134 29972 10140
rect 30012 10192 30064 10198
rect 30012 10134 30064 10140
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29276 10056 29328 10062
rect 29276 9998 29328 10004
rect 29184 9920 29236 9926
rect 29184 9862 29236 9868
rect 29000 9716 29052 9722
rect 29000 9658 29052 9664
rect 29196 9586 29224 9862
rect 29184 9580 29236 9586
rect 29184 9522 29236 9528
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29012 8634 29040 8978
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 28908 8560 28960 8566
rect 28908 8502 28960 8508
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 28448 8356 28500 8362
rect 28448 8298 28500 8304
rect 28460 8090 28488 8298
rect 28552 8090 28580 8366
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28448 8084 28500 8090
rect 28448 8026 28500 8032
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 28644 7954 28672 8230
rect 28816 8084 28868 8090
rect 28816 8026 28868 8032
rect 28540 7948 28592 7954
rect 28540 7890 28592 7896
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 27896 7336 27948 7342
rect 27896 7278 27948 7284
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 28356 7336 28408 7342
rect 28356 7278 28408 7284
rect 26608 7268 26660 7274
rect 26608 7210 26660 7216
rect 26516 6996 26568 7002
rect 26516 6938 26568 6944
rect 26332 6928 26384 6934
rect 26332 6870 26384 6876
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26620 6730 26648 7210
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 26792 7200 26844 7206
rect 26792 7142 26844 7148
rect 26608 6724 26660 6730
rect 26608 6666 26660 6672
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26056 5772 26108 5778
rect 26056 5714 26108 5720
rect 25228 4684 25280 4690
rect 25228 4626 25280 4632
rect 25964 4684 26016 4690
rect 25964 4626 26016 4632
rect 26068 4622 26096 5714
rect 26160 5234 26188 6258
rect 26344 6254 26372 6598
rect 26332 6248 26384 6254
rect 26332 6190 26384 6196
rect 26436 6186 26464 6598
rect 26424 6180 26476 6186
rect 26424 6122 26476 6128
rect 26620 5846 26648 6666
rect 26712 6458 26740 7142
rect 26804 6866 26832 7142
rect 27644 7100 27952 7109
rect 27644 7098 27650 7100
rect 27706 7098 27730 7100
rect 27786 7098 27810 7100
rect 27866 7098 27890 7100
rect 27946 7098 27952 7100
rect 27706 7046 27708 7098
rect 27888 7046 27890 7098
rect 27644 7044 27650 7046
rect 27706 7044 27730 7046
rect 27786 7044 27810 7046
rect 27866 7044 27890 7046
rect 27946 7044 27952 7046
rect 27644 7035 27952 7044
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 26984 6556 27292 6565
rect 26984 6554 26990 6556
rect 27046 6554 27070 6556
rect 27126 6554 27150 6556
rect 27206 6554 27230 6556
rect 27286 6554 27292 6556
rect 27046 6502 27048 6554
rect 27228 6502 27230 6554
rect 26984 6500 26990 6502
rect 27046 6500 27070 6502
rect 27126 6500 27150 6502
rect 27206 6500 27230 6502
rect 27286 6500 27292 6502
rect 26984 6491 27292 6500
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 27448 6254 27476 6598
rect 27436 6248 27488 6254
rect 26698 6216 26754 6225
rect 27436 6190 27488 6196
rect 26698 6151 26754 6160
rect 26712 6118 26740 6151
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 27644 6012 27952 6021
rect 27644 6010 27650 6012
rect 27706 6010 27730 6012
rect 27786 6010 27810 6012
rect 27866 6010 27890 6012
rect 27946 6010 27952 6012
rect 27706 5958 27708 6010
rect 27888 5958 27890 6010
rect 27644 5956 27650 5958
rect 27706 5956 27730 5958
rect 27786 5956 27810 5958
rect 27866 5956 27890 5958
rect 27946 5956 27952 5958
rect 27644 5947 27952 5956
rect 26608 5840 26660 5846
rect 26608 5782 26660 5788
rect 26984 5468 27292 5477
rect 26984 5466 26990 5468
rect 27046 5466 27070 5468
rect 27126 5466 27150 5468
rect 27206 5466 27230 5468
rect 27286 5466 27292 5468
rect 27046 5414 27048 5466
rect 27228 5414 27230 5466
rect 26984 5412 26990 5414
rect 27046 5412 27070 5414
rect 27126 5412 27150 5414
rect 27206 5412 27230 5414
rect 27286 5412 27292 5414
rect 26984 5403 27292 5412
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26056 4616 26108 4622
rect 26056 4558 26108 4564
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25240 3738 25268 4014
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25228 3732 25280 3738
rect 25228 3674 25280 3680
rect 24584 3528 24636 3534
rect 22204 3454 22324 3482
rect 24584 3470 24636 3476
rect 22296 3194 22324 3454
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21284 2650 21312 2858
rect 22112 2774 22140 3130
rect 22112 2746 22232 2774
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21638 2544 21694 2553
rect 20904 2508 20956 2514
rect 22204 2514 22232 2746
rect 21638 2479 21640 2488
rect 20904 2450 20956 2456
rect 21692 2479 21694 2488
rect 22192 2508 22244 2514
rect 21640 2450 21692 2456
rect 22192 2450 22244 2456
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 20088 2038 20116 2246
rect 20076 2032 20128 2038
rect 20076 1974 20128 1980
rect 20088 1902 20116 1974
rect 20364 1902 20392 2382
rect 20444 2032 20496 2038
rect 20444 1974 20496 1980
rect 20456 1902 20484 1974
rect 19156 1896 19208 1902
rect 19156 1838 19208 1844
rect 19708 1896 19760 1902
rect 19708 1838 19760 1844
rect 20076 1896 20128 1902
rect 20076 1838 20128 1844
rect 20352 1896 20404 1902
rect 20352 1838 20404 1844
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 19064 1556 19116 1562
rect 19064 1498 19116 1504
rect 19168 1426 19196 1838
rect 19432 1760 19484 1766
rect 19432 1702 19484 1708
rect 19616 1760 19668 1766
rect 19616 1702 19668 1708
rect 19444 1494 19472 1702
rect 19432 1488 19484 1494
rect 19432 1430 19484 1436
rect 19628 1426 19656 1702
rect 19720 1562 19748 1838
rect 22388 1834 22416 3402
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22664 2553 22692 3334
rect 22650 2544 22706 2553
rect 22650 2479 22652 2488
rect 22704 2479 22706 2488
rect 22652 2450 22704 2456
rect 22848 1902 22876 3334
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23112 2440 23164 2446
rect 23112 2382 23164 2388
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22836 1896 22888 1902
rect 22836 1838 22888 1844
rect 22376 1828 22428 1834
rect 22376 1770 22428 1776
rect 20628 1760 20680 1766
rect 20628 1702 20680 1708
rect 22652 1760 22704 1766
rect 22652 1702 22704 1708
rect 19870 1660 20178 1669
rect 19870 1658 19876 1660
rect 19932 1658 19956 1660
rect 20012 1658 20036 1660
rect 20092 1658 20116 1660
rect 20172 1658 20178 1660
rect 19932 1606 19934 1658
rect 20114 1606 20116 1658
rect 19870 1604 19876 1606
rect 19932 1604 19956 1606
rect 20012 1604 20036 1606
rect 20092 1604 20116 1606
rect 20172 1604 20178 1606
rect 19870 1595 20178 1604
rect 20640 1562 20668 1702
rect 19708 1556 19760 1562
rect 19708 1498 19760 1504
rect 20628 1556 20680 1562
rect 20628 1498 20680 1504
rect 22664 1426 22692 1702
rect 23032 1562 23060 2246
rect 23124 1902 23152 2382
rect 23308 2378 23336 2858
rect 23676 2378 23704 2926
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 23296 2372 23348 2378
rect 23296 2314 23348 2320
rect 23664 2372 23716 2378
rect 23664 2314 23716 2320
rect 23768 1970 23796 2450
rect 23756 1964 23808 1970
rect 23756 1906 23808 1912
rect 23112 1896 23164 1902
rect 23112 1838 23164 1844
rect 23204 1896 23256 1902
rect 23204 1838 23256 1844
rect 23020 1556 23072 1562
rect 23020 1498 23072 1504
rect 19156 1420 19208 1426
rect 19156 1362 19208 1368
rect 19616 1420 19668 1426
rect 19616 1362 19668 1368
rect 22652 1420 22704 1426
rect 22652 1362 22704 1368
rect 19168 1222 19196 1362
rect 23124 1290 23152 1838
rect 23216 1766 23244 1838
rect 23204 1760 23256 1766
rect 23204 1702 23256 1708
rect 23112 1284 23164 1290
rect 23112 1226 23164 1232
rect 23952 1222 23980 2450
rect 24044 2038 24072 2790
rect 24136 2514 24164 2790
rect 24412 2514 24440 2994
rect 24492 2576 24544 2582
rect 24492 2518 24544 2524
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 24032 2032 24084 2038
rect 24032 1974 24084 1980
rect 24044 1426 24072 1974
rect 24136 1562 24164 2450
rect 24504 2106 24532 2518
rect 24688 2514 24716 3674
rect 24952 3460 25004 3466
rect 24952 3402 25004 3408
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24216 2100 24268 2106
rect 24216 2042 24268 2048
rect 24492 2100 24544 2106
rect 24492 2042 24544 2048
rect 24228 1986 24256 2042
rect 24596 1986 24624 2382
rect 24872 1986 24900 2450
rect 24228 1958 24624 1986
rect 24688 1958 24900 1986
rect 24688 1902 24716 1958
rect 24676 1896 24728 1902
rect 24964 1850 24992 3402
rect 25148 2854 25176 3674
rect 25136 2848 25188 2854
rect 25136 2790 25188 2796
rect 25240 2774 25268 3674
rect 26160 3602 26188 5170
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 27172 4826 27200 5102
rect 27644 4924 27952 4933
rect 27644 4922 27650 4924
rect 27706 4922 27730 4924
rect 27786 4922 27810 4924
rect 27866 4922 27890 4924
rect 27946 4922 27952 4924
rect 27706 4870 27708 4922
rect 27888 4870 27890 4922
rect 27644 4868 27650 4870
rect 27706 4868 27730 4870
rect 27786 4868 27810 4870
rect 27866 4868 27890 4870
rect 27946 4868 27952 4870
rect 27644 4859 27952 4868
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 26896 4146 26924 4422
rect 26984 4380 27292 4389
rect 26984 4378 26990 4380
rect 27046 4378 27070 4380
rect 27126 4378 27150 4380
rect 27206 4378 27230 4380
rect 27286 4378 27292 4380
rect 27046 4326 27048 4378
rect 27228 4326 27230 4378
rect 26984 4324 26990 4326
rect 27046 4324 27070 4326
rect 27126 4324 27150 4326
rect 27206 4324 27230 4326
rect 27286 4324 27292 4326
rect 26984 4315 27292 4324
rect 27632 4282 27660 4422
rect 28000 4298 28028 5102
rect 28092 5098 28120 7278
rect 28552 7206 28580 7890
rect 28632 7744 28684 7750
rect 28632 7686 28684 7692
rect 28644 7342 28672 7686
rect 28828 7546 28856 8026
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 29104 7342 29132 8434
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 29012 5846 29040 6802
rect 29196 6798 29224 9522
rect 29276 9376 29328 9382
rect 29276 9318 29328 9324
rect 29288 9042 29316 9318
rect 29276 9036 29328 9042
rect 29276 8978 29328 8984
rect 29472 8838 29500 10066
rect 29932 9722 29960 10134
rect 30760 10130 30788 10406
rect 30748 10124 30800 10130
rect 30748 10066 30800 10072
rect 29920 9716 29972 9722
rect 29920 9658 29972 9664
rect 29460 8832 29512 8838
rect 29460 8774 29512 8780
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 29472 8430 29500 8774
rect 29460 8424 29512 8430
rect 29460 8366 29512 8372
rect 29276 8356 29328 8362
rect 29276 8298 29328 8304
rect 29288 8022 29316 8298
rect 29276 8016 29328 8022
rect 29276 7958 29328 7964
rect 29472 7954 29500 8366
rect 30668 8362 30696 8774
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 29460 7948 29512 7954
rect 29460 7890 29512 7896
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 7546 30144 7686
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 29920 7200 29972 7206
rect 29920 7142 29972 7148
rect 29644 6860 29696 6866
rect 29644 6802 29696 6808
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 29656 6458 29684 6802
rect 29840 6458 29868 6802
rect 29644 6452 29696 6458
rect 29644 6394 29696 6400
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 29932 6254 29960 7142
rect 30668 6866 30696 8298
rect 30748 8288 30800 8294
rect 30748 8230 30800 8236
rect 30760 8022 30788 8230
rect 30748 8016 30800 8022
rect 30748 7958 30800 7964
rect 30852 7954 30880 10678
rect 30840 7948 30892 7954
rect 30840 7890 30892 7896
rect 30104 6860 30156 6866
rect 30104 6802 30156 6808
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30116 6458 30144 6802
rect 30194 6760 30250 6769
rect 30194 6695 30196 6704
rect 30248 6695 30250 6704
rect 30196 6666 30248 6672
rect 30392 6662 30420 6802
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 30392 6186 30420 6598
rect 30668 6254 30696 6802
rect 30656 6248 30708 6254
rect 30656 6190 30708 6196
rect 30380 6180 30432 6186
rect 30380 6122 30432 6128
rect 28632 5840 28684 5846
rect 28632 5782 28684 5788
rect 29000 5840 29052 5846
rect 29000 5782 29052 5788
rect 28172 5772 28224 5778
rect 28172 5714 28224 5720
rect 28448 5772 28500 5778
rect 28448 5714 28500 5720
rect 28184 5370 28212 5714
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 28264 5160 28316 5166
rect 28264 5102 28316 5108
rect 28080 5092 28132 5098
rect 28080 5034 28132 5040
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27908 4270 28028 4298
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 26896 3670 26924 4082
rect 27252 4072 27304 4078
rect 27252 4014 27304 4020
rect 26884 3664 26936 3670
rect 26884 3606 26936 3612
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26160 2922 26188 3538
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26528 3194 26556 3470
rect 27264 3466 27292 4014
rect 27908 4010 27936 4270
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 27896 4004 27948 4010
rect 27896 3946 27948 3952
rect 27644 3836 27952 3845
rect 27644 3834 27650 3836
rect 27706 3834 27730 3836
rect 27786 3834 27810 3836
rect 27866 3834 27890 3836
rect 27946 3834 27952 3836
rect 27706 3782 27708 3834
rect 27888 3782 27890 3834
rect 27644 3780 27650 3782
rect 27706 3780 27730 3782
rect 27786 3780 27810 3782
rect 27866 3780 27890 3782
rect 27946 3780 27952 3782
rect 27644 3771 27952 3780
rect 28000 3670 28028 4014
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 28092 3534 28120 5034
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 28184 4486 28212 4966
rect 28276 4758 28304 5102
rect 28460 4758 28488 5714
rect 28540 5636 28592 5642
rect 28540 5578 28592 5584
rect 28552 4826 28580 5578
rect 28644 5030 28672 5782
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28736 5166 28764 5714
rect 29012 5302 29040 5782
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 28724 5160 28776 5166
rect 28724 5102 28776 5108
rect 28632 5024 28684 5030
rect 28632 4966 28684 4972
rect 28540 4820 28592 4826
rect 28540 4762 28592 4768
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 28448 4752 28500 4758
rect 28448 4694 28500 4700
rect 28460 4554 28488 4694
rect 28448 4548 28500 4554
rect 28448 4490 28500 4496
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 28644 4010 28672 4966
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28632 4004 28684 4010
rect 28632 3946 28684 3952
rect 28644 3618 28672 3946
rect 28920 3942 28948 4626
rect 29012 4486 29040 5238
rect 29104 4758 29132 5510
rect 29564 5370 29592 5510
rect 29552 5364 29604 5370
rect 29552 5306 29604 5312
rect 29092 4752 29144 4758
rect 29092 4694 29144 4700
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 29000 4072 29052 4078
rect 29000 4014 29052 4020
rect 28908 3936 28960 3942
rect 28908 3878 28960 3884
rect 29012 3738 29040 4014
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 30392 3670 30420 6122
rect 30932 5024 30984 5030
rect 30932 4966 30984 4972
rect 30944 4690 30972 4966
rect 30932 4684 30984 4690
rect 30932 4626 30984 4632
rect 28460 3590 28672 3618
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 28080 3528 28132 3534
rect 28080 3470 28132 3476
rect 27252 3460 27304 3466
rect 27252 3402 27304 3408
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26620 2990 26648 3334
rect 26984 3292 27292 3301
rect 26984 3290 26990 3292
rect 27046 3290 27070 3292
rect 27126 3290 27150 3292
rect 27206 3290 27230 3292
rect 27286 3290 27292 3292
rect 27046 3238 27048 3290
rect 27228 3238 27230 3290
rect 26984 3236 26990 3238
rect 27046 3236 27070 3238
rect 27126 3236 27150 3238
rect 27206 3236 27230 3238
rect 27286 3236 27292 3238
rect 26984 3227 27292 3236
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26700 3120 26752 3126
rect 26700 3062 26752 3068
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26148 2916 26200 2922
rect 26148 2858 26200 2864
rect 25240 2746 25360 2774
rect 25332 2514 25360 2746
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 25136 2372 25188 2378
rect 25136 2314 25188 2320
rect 25148 1902 25176 2314
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 25688 2304 25740 2310
rect 25688 2246 25740 2252
rect 25240 1970 25268 2246
rect 25700 2106 25728 2246
rect 25688 2100 25740 2106
rect 25688 2042 25740 2048
rect 25228 1964 25280 1970
rect 25228 1906 25280 1912
rect 24676 1838 24728 1844
rect 24872 1822 24992 1850
rect 25136 1896 25188 1902
rect 25136 1838 25188 1844
rect 25792 1834 25820 2450
rect 26160 2106 26188 2858
rect 26712 2650 26740 3062
rect 27080 2990 27108 3130
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 26792 2916 26844 2922
rect 26792 2858 26844 2864
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 26516 2576 26568 2582
rect 26516 2518 26568 2524
rect 26240 2372 26292 2378
rect 26240 2314 26292 2320
rect 26148 2100 26200 2106
rect 26148 2042 26200 2048
rect 25780 1828 25832 1834
rect 24872 1766 24900 1822
rect 25780 1770 25832 1776
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 25792 1562 25820 1770
rect 25872 1760 25924 1766
rect 25872 1702 25924 1708
rect 24124 1556 24176 1562
rect 24124 1498 24176 1504
rect 25780 1556 25832 1562
rect 25780 1498 25832 1504
rect 25884 1494 25912 1702
rect 25872 1488 25924 1494
rect 25872 1430 25924 1436
rect 24032 1420 24084 1426
rect 24032 1362 24084 1368
rect 26252 1358 26280 2314
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 26436 1970 26464 2246
rect 26424 1964 26476 1970
rect 26424 1906 26476 1912
rect 26528 1902 26556 2518
rect 26712 2378 26740 2586
rect 26700 2372 26752 2378
rect 26700 2314 26752 2320
rect 26516 1896 26568 1902
rect 26516 1838 26568 1844
rect 26804 1766 26832 2858
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26424 1760 26476 1766
rect 26424 1702 26476 1708
rect 26792 1760 26844 1766
rect 26792 1702 26844 1708
rect 26436 1358 26464 1702
rect 26896 1562 26924 2586
rect 27080 2514 27108 2926
rect 27448 2582 27476 2994
rect 28092 2990 28120 3470
rect 28356 3392 28408 3398
rect 28356 3334 28408 3340
rect 28368 3194 28396 3334
rect 28356 3188 28408 3194
rect 28356 3130 28408 3136
rect 28080 2984 28132 2990
rect 28080 2926 28132 2932
rect 27988 2848 28040 2854
rect 27988 2790 28040 2796
rect 27644 2748 27952 2757
rect 27644 2746 27650 2748
rect 27706 2746 27730 2748
rect 27786 2746 27810 2748
rect 27866 2746 27890 2748
rect 27946 2746 27952 2748
rect 27706 2694 27708 2746
rect 27888 2694 27890 2746
rect 27644 2692 27650 2694
rect 27706 2692 27730 2694
rect 27786 2692 27810 2694
rect 27866 2692 27890 2694
rect 27946 2692 27952 2694
rect 27644 2683 27952 2692
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 27068 2508 27120 2514
rect 27068 2450 27120 2456
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 27436 2304 27488 2310
rect 27436 2246 27488 2252
rect 26984 2204 27292 2213
rect 26984 2202 26990 2204
rect 27046 2202 27070 2204
rect 27126 2202 27150 2204
rect 27206 2202 27230 2204
rect 27286 2202 27292 2204
rect 27046 2150 27048 2202
rect 27228 2150 27230 2202
rect 26984 2148 26990 2150
rect 27046 2148 27070 2150
rect 27126 2148 27150 2150
rect 27206 2148 27230 2150
rect 27286 2148 27292 2150
rect 26984 2139 27292 2148
rect 26976 1828 27028 1834
rect 26976 1770 27028 1776
rect 26988 1562 27016 1770
rect 27356 1562 27384 2246
rect 26884 1556 26936 1562
rect 26884 1498 26936 1504
rect 26976 1556 27028 1562
rect 26976 1498 27028 1504
rect 27344 1556 27396 1562
rect 27344 1498 27396 1504
rect 26240 1352 26292 1358
rect 26240 1294 26292 1300
rect 26424 1352 26476 1358
rect 26424 1294 26476 1300
rect 27448 1222 27476 2246
rect 27632 2106 27660 2450
rect 28000 2378 28028 2790
rect 28092 2446 28120 2926
rect 28460 2922 28488 3590
rect 30392 3194 30420 3606
rect 30380 3188 30432 3194
rect 30380 3130 30432 3136
rect 28264 2916 28316 2922
rect 28264 2858 28316 2864
rect 28448 2916 28500 2922
rect 28448 2858 28500 2864
rect 28276 2650 28304 2858
rect 28264 2644 28316 2650
rect 28264 2586 28316 2592
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 27988 2372 28040 2378
rect 27988 2314 28040 2320
rect 27620 2100 27672 2106
rect 27620 2042 27672 2048
rect 28092 1902 28120 2382
rect 28908 2032 28960 2038
rect 28908 1974 28960 1980
rect 28080 1896 28132 1902
rect 28080 1838 28132 1844
rect 27988 1760 28040 1766
rect 27988 1702 28040 1708
rect 27644 1660 27952 1669
rect 27644 1658 27650 1660
rect 27706 1658 27730 1660
rect 27786 1658 27810 1660
rect 27866 1658 27890 1660
rect 27946 1658 27952 1660
rect 27706 1606 27708 1658
rect 27888 1606 27890 1658
rect 27644 1604 27650 1606
rect 27706 1604 27730 1606
rect 27786 1604 27810 1606
rect 27866 1604 27890 1606
rect 27946 1604 27952 1606
rect 27644 1595 27952 1604
rect 28000 1494 28028 1702
rect 28920 1562 28948 1974
rect 28908 1556 28960 1562
rect 28908 1498 28960 1504
rect 27988 1488 28040 1494
rect 27988 1430 28040 1436
rect 19156 1216 19208 1222
rect 19156 1158 19208 1164
rect 19616 1216 19668 1222
rect 19616 1158 19668 1164
rect 23940 1216 23992 1222
rect 23940 1158 23992 1164
rect 27436 1216 27488 1222
rect 27436 1158 27488 1164
rect 19210 1116 19518 1125
rect 19210 1114 19216 1116
rect 19272 1114 19296 1116
rect 19352 1114 19376 1116
rect 19432 1114 19456 1116
rect 19512 1114 19518 1116
rect 19272 1062 19274 1114
rect 19454 1062 19456 1114
rect 19210 1060 19216 1062
rect 19272 1060 19296 1062
rect 19352 1060 19376 1062
rect 19432 1060 19456 1062
rect 19512 1060 19518 1062
rect 19210 1051 19518 1060
rect 19628 814 19656 1158
rect 26984 1116 27292 1125
rect 26984 1114 26990 1116
rect 27046 1114 27070 1116
rect 27126 1114 27150 1116
rect 27206 1114 27230 1116
rect 27286 1114 27292 1116
rect 27046 1062 27048 1114
rect 27228 1062 27230 1114
rect 26984 1060 26990 1062
rect 27046 1060 27070 1062
rect 27126 1060 27150 1062
rect 27206 1060 27230 1062
rect 27286 1060 27292 1062
rect 26984 1051 27292 1060
rect 19616 808 19668 814
rect 19616 750 19668 756
rect 7472 740 7524 746
rect 7472 682 7524 688
rect 18880 740 18932 746
rect 18880 682 18932 688
rect 18972 740 19024 746
rect 18972 682 19024 688
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 12096 572 12404 581
rect 12096 570 12102 572
rect 12158 570 12182 572
rect 12238 570 12262 572
rect 12318 570 12342 572
rect 12398 570 12404 572
rect 12158 518 12160 570
rect 12340 518 12342 570
rect 12096 516 12102 518
rect 12158 516 12182 518
rect 12238 516 12262 518
rect 12318 516 12342 518
rect 12398 516 12404 518
rect 12096 507 12404 516
rect 19870 572 20178 581
rect 19870 570 19876 572
rect 19932 570 19956 572
rect 20012 570 20036 572
rect 20092 570 20116 572
rect 20172 570 20178 572
rect 19932 518 19934 570
rect 20114 518 20116 570
rect 19870 516 19876 518
rect 19932 516 19956 518
rect 20012 516 20036 518
rect 20092 516 20116 518
rect 20172 516 20178 518
rect 19870 507 20178 516
rect 27644 572 27952 581
rect 27644 570 27650 572
rect 27706 570 27730 572
rect 27786 570 27810 572
rect 27866 570 27890 572
rect 27946 570 27952 572
rect 27706 518 27708 570
rect 27888 518 27890 570
rect 27644 516 27650 518
rect 27706 516 27730 518
rect 27786 516 27810 518
rect 27866 516 27890 518
rect 27946 516 27952 518
rect 27644 507 27952 516
<< via2 >>
rect 11794 21936 11850 21992
rect 12254 21936 12310 21992
rect 24398 21936 24454 21992
rect 27342 21936 27398 21992
rect 27710 21936 27766 21992
rect 8666 21800 8722 21856
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 6090 21684 6146 21720
rect 6090 21664 6092 21684
rect 6092 21664 6144 21684
rect 6144 21664 6146 21684
rect 8022 21684 8078 21720
rect 8022 21664 8024 21684
rect 8024 21664 8076 21684
rect 8076 21664 8078 21684
rect 8390 21684 8446 21720
rect 11442 21786 11498 21788
rect 11522 21786 11578 21788
rect 11602 21786 11658 21788
rect 11682 21786 11738 21788
rect 11442 21734 11488 21786
rect 11488 21734 11498 21786
rect 11522 21734 11552 21786
rect 11552 21734 11564 21786
rect 11564 21734 11578 21786
rect 11602 21734 11616 21786
rect 11616 21734 11628 21786
rect 11628 21734 11658 21786
rect 11682 21734 11692 21786
rect 11692 21734 11738 21786
rect 11442 21732 11498 21734
rect 11522 21732 11578 21734
rect 11602 21732 11658 21734
rect 11682 21732 11738 21734
rect 22190 21800 22246 21856
rect 23846 21800 23902 21856
rect 19216 21786 19272 21788
rect 19296 21786 19352 21788
rect 19376 21786 19432 21788
rect 19456 21786 19512 21788
rect 19216 21734 19262 21786
rect 19262 21734 19272 21786
rect 19296 21734 19326 21786
rect 19326 21734 19338 21786
rect 19338 21734 19352 21786
rect 19376 21734 19390 21786
rect 19390 21734 19402 21786
rect 19402 21734 19432 21786
rect 19456 21734 19466 21786
rect 19466 21734 19512 21786
rect 19216 21732 19272 21734
rect 19296 21732 19352 21734
rect 19376 21732 19432 21734
rect 19456 21732 19512 21734
rect 8390 21664 8392 21684
rect 8392 21664 8444 21684
rect 8444 21664 8446 21684
rect 12990 21684 13046 21720
rect 12990 21664 12992 21684
rect 12992 21664 13044 21684
rect 13044 21664 13046 21684
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 6734 20324 6790 20360
rect 6734 20304 6736 20324
rect 6736 20304 6788 20324
rect 6788 20304 6790 20324
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 4158 17620 4160 17640
rect 4160 17620 4212 17640
rect 4212 17620 4214 17640
rect 4158 17584 4214 17620
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 4710 17584 4766 17640
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 4986 17584 5042 17640
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 4986 14864 5042 14920
rect 4986 14592 5042 14648
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 8942 21256 8998 21312
rect 8574 21140 8630 21176
rect 12102 21242 12158 21244
rect 12182 21242 12238 21244
rect 12262 21242 12318 21244
rect 12342 21242 12398 21244
rect 12102 21190 12148 21242
rect 12148 21190 12158 21242
rect 12182 21190 12212 21242
rect 12212 21190 12224 21242
rect 12224 21190 12238 21242
rect 12262 21190 12276 21242
rect 12276 21190 12288 21242
rect 12288 21190 12318 21242
rect 12342 21190 12352 21242
rect 12352 21190 12398 21242
rect 12102 21188 12158 21190
rect 12182 21188 12238 21190
rect 12262 21188 12318 21190
rect 12342 21188 12398 21190
rect 8574 21120 8576 21140
rect 8576 21120 8628 21140
rect 8628 21120 8630 21140
rect 9770 21140 9826 21176
rect 9770 21120 9772 21140
rect 9772 21120 9824 21140
rect 9824 21120 9826 21140
rect 7838 18808 7894 18864
rect 6090 17076 6092 17096
rect 6092 17076 6144 17096
rect 6144 17076 6146 17096
rect 6090 17040 6146 17076
rect 6458 17040 6514 17096
rect 5630 14320 5686 14376
rect 8206 19216 8262 19272
rect 8666 18672 8722 18728
rect 8942 19352 8998 19408
rect 11058 20576 11114 20632
rect 9954 20460 10010 20496
rect 9954 20440 9956 20460
rect 9956 20440 10008 20460
rect 10008 20440 10010 20460
rect 11442 20698 11498 20700
rect 11522 20698 11578 20700
rect 11602 20698 11658 20700
rect 11682 20698 11738 20700
rect 11442 20646 11488 20698
rect 11488 20646 11498 20698
rect 11522 20646 11552 20698
rect 11552 20646 11564 20698
rect 11564 20646 11578 20698
rect 11602 20646 11616 20698
rect 11616 20646 11628 20698
rect 11628 20646 11658 20698
rect 11682 20646 11692 20698
rect 11692 20646 11738 20698
rect 11442 20644 11498 20646
rect 11522 20644 11578 20646
rect 11602 20644 11658 20646
rect 11682 20644 11738 20646
rect 12102 20154 12158 20156
rect 12182 20154 12238 20156
rect 12262 20154 12318 20156
rect 12342 20154 12398 20156
rect 12102 20102 12148 20154
rect 12148 20102 12158 20154
rect 12182 20102 12212 20154
rect 12212 20102 12224 20154
rect 12224 20102 12238 20154
rect 12262 20102 12276 20154
rect 12276 20102 12288 20154
rect 12288 20102 12318 20154
rect 12342 20102 12352 20154
rect 12352 20102 12398 20154
rect 12102 20100 12158 20102
rect 12182 20100 12238 20102
rect 12262 20100 12318 20102
rect 12342 20100 12398 20102
rect 10690 19352 10746 19408
rect 10046 17856 10102 17912
rect 11442 19610 11498 19612
rect 11522 19610 11578 19612
rect 11602 19610 11658 19612
rect 11682 19610 11738 19612
rect 11442 19558 11488 19610
rect 11488 19558 11498 19610
rect 11522 19558 11552 19610
rect 11552 19558 11564 19610
rect 11564 19558 11578 19610
rect 11602 19558 11616 19610
rect 11616 19558 11628 19610
rect 11628 19558 11658 19610
rect 11682 19558 11692 19610
rect 11692 19558 11738 19610
rect 11442 19556 11498 19558
rect 11522 19556 11578 19558
rect 11602 19556 11658 19558
rect 11682 19556 11738 19558
rect 10782 17856 10838 17912
rect 10598 17720 10654 17776
rect 10414 17176 10470 17232
rect 12102 19066 12158 19068
rect 12182 19066 12238 19068
rect 12262 19066 12318 19068
rect 12342 19066 12398 19068
rect 12102 19014 12148 19066
rect 12148 19014 12158 19066
rect 12182 19014 12212 19066
rect 12212 19014 12224 19066
rect 12224 19014 12238 19066
rect 12262 19014 12276 19066
rect 12276 19014 12288 19066
rect 12288 19014 12318 19066
rect 12342 19014 12352 19066
rect 12352 19014 12398 19066
rect 12102 19012 12158 19014
rect 12182 19012 12238 19014
rect 12262 19012 12318 19014
rect 12342 19012 12398 19014
rect 13266 20576 13322 20632
rect 18050 21412 18106 21448
rect 18050 21392 18052 21412
rect 18052 21392 18104 21412
rect 18104 21392 18106 21412
rect 11442 18522 11498 18524
rect 11522 18522 11578 18524
rect 11602 18522 11658 18524
rect 11682 18522 11738 18524
rect 11442 18470 11488 18522
rect 11488 18470 11498 18522
rect 11522 18470 11552 18522
rect 11552 18470 11564 18522
rect 11564 18470 11578 18522
rect 11602 18470 11616 18522
rect 11616 18470 11628 18522
rect 11628 18470 11658 18522
rect 11682 18470 11692 18522
rect 11692 18470 11738 18522
rect 11442 18468 11498 18470
rect 11522 18468 11578 18470
rect 11602 18468 11658 18470
rect 11682 18468 11738 18470
rect 11610 17620 11612 17640
rect 11612 17620 11664 17640
rect 11664 17620 11666 17640
rect 11610 17584 11666 17620
rect 11442 17434 11498 17436
rect 11522 17434 11578 17436
rect 11602 17434 11658 17436
rect 11682 17434 11738 17436
rect 11442 17382 11488 17434
rect 11488 17382 11498 17434
rect 11522 17382 11552 17434
rect 11552 17382 11564 17434
rect 11564 17382 11578 17434
rect 11602 17382 11616 17434
rect 11616 17382 11628 17434
rect 11628 17382 11658 17434
rect 11682 17382 11692 17434
rect 11692 17382 11738 17434
rect 11442 17380 11498 17382
rect 11522 17380 11578 17382
rect 11602 17380 11658 17382
rect 11682 17380 11738 17382
rect 12102 17978 12158 17980
rect 12182 17978 12238 17980
rect 12262 17978 12318 17980
rect 12342 17978 12398 17980
rect 12102 17926 12148 17978
rect 12148 17926 12158 17978
rect 12182 17926 12212 17978
rect 12212 17926 12224 17978
rect 12224 17926 12238 17978
rect 12262 17926 12276 17978
rect 12276 17926 12288 17978
rect 12288 17926 12318 17978
rect 12342 17926 12352 17978
rect 12352 17926 12398 17978
rect 12102 17924 12158 17926
rect 12182 17924 12238 17926
rect 12262 17924 12318 17926
rect 12342 17924 12398 17926
rect 11426 17040 11482 17096
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 9494 13796 9550 13832
rect 9494 13776 9496 13796
rect 9496 13776 9548 13796
rect 9548 13776 9550 13796
rect 9954 13912 10010 13968
rect 12102 16890 12158 16892
rect 12182 16890 12238 16892
rect 12262 16890 12318 16892
rect 12342 16890 12398 16892
rect 12102 16838 12148 16890
rect 12148 16838 12158 16890
rect 12182 16838 12212 16890
rect 12212 16838 12224 16890
rect 12224 16838 12238 16890
rect 12262 16838 12276 16890
rect 12276 16838 12288 16890
rect 12288 16838 12318 16890
rect 12342 16838 12352 16890
rect 12352 16838 12398 16890
rect 12102 16836 12158 16838
rect 12182 16836 12238 16838
rect 12262 16836 12318 16838
rect 12342 16836 12398 16838
rect 11442 16346 11498 16348
rect 11522 16346 11578 16348
rect 11602 16346 11658 16348
rect 11682 16346 11738 16348
rect 11442 16294 11488 16346
rect 11488 16294 11498 16346
rect 11522 16294 11552 16346
rect 11552 16294 11564 16346
rect 11564 16294 11578 16346
rect 11602 16294 11616 16346
rect 11616 16294 11628 16346
rect 11628 16294 11658 16346
rect 11682 16294 11692 16346
rect 11692 16294 11738 16346
rect 11442 16292 11498 16294
rect 11522 16292 11578 16294
rect 11602 16292 11658 16294
rect 11682 16292 11738 16294
rect 11442 15258 11498 15260
rect 11522 15258 11578 15260
rect 11602 15258 11658 15260
rect 11682 15258 11738 15260
rect 11442 15206 11488 15258
rect 11488 15206 11498 15258
rect 11522 15206 11552 15258
rect 11552 15206 11564 15258
rect 11564 15206 11578 15258
rect 11602 15206 11616 15258
rect 11616 15206 11628 15258
rect 11628 15206 11658 15258
rect 11682 15206 11692 15258
rect 11692 15206 11738 15258
rect 11442 15204 11498 15206
rect 11522 15204 11578 15206
rect 11602 15204 11658 15206
rect 11682 15204 11738 15206
rect 12102 15802 12158 15804
rect 12182 15802 12238 15804
rect 12262 15802 12318 15804
rect 12342 15802 12398 15804
rect 12102 15750 12148 15802
rect 12148 15750 12158 15802
rect 12182 15750 12212 15802
rect 12212 15750 12224 15802
rect 12224 15750 12238 15802
rect 12262 15750 12276 15802
rect 12276 15750 12288 15802
rect 12288 15750 12318 15802
rect 12342 15750 12352 15802
rect 12352 15750 12398 15802
rect 12102 15748 12158 15750
rect 12182 15748 12238 15750
rect 12262 15748 12318 15750
rect 12342 15748 12398 15750
rect 11442 14170 11498 14172
rect 11522 14170 11578 14172
rect 11602 14170 11658 14172
rect 11682 14170 11738 14172
rect 11442 14118 11488 14170
rect 11488 14118 11498 14170
rect 11522 14118 11552 14170
rect 11552 14118 11564 14170
rect 11564 14118 11578 14170
rect 11602 14118 11616 14170
rect 11616 14118 11628 14170
rect 11628 14118 11658 14170
rect 11682 14118 11692 14170
rect 11692 14118 11738 14170
rect 11442 14116 11498 14118
rect 11522 14116 11578 14118
rect 11602 14116 11658 14118
rect 11682 14116 11738 14118
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 1766 4528 1822 4584
rect 2686 4528 2742 4584
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 9862 7948 9918 7984
rect 9862 7928 9864 7948
rect 9864 7928 9916 7948
rect 9916 7928 9918 7948
rect 12102 14714 12158 14716
rect 12182 14714 12238 14716
rect 12262 14714 12318 14716
rect 12342 14714 12398 14716
rect 12102 14662 12148 14714
rect 12148 14662 12158 14714
rect 12182 14662 12212 14714
rect 12212 14662 12224 14714
rect 12224 14662 12238 14714
rect 12262 14662 12276 14714
rect 12276 14662 12288 14714
rect 12288 14662 12318 14714
rect 12342 14662 12352 14714
rect 12352 14662 12398 14714
rect 12102 14660 12158 14662
rect 12182 14660 12238 14662
rect 12262 14660 12318 14662
rect 12342 14660 12398 14662
rect 12102 13626 12158 13628
rect 12182 13626 12238 13628
rect 12262 13626 12318 13628
rect 12342 13626 12398 13628
rect 12102 13574 12148 13626
rect 12148 13574 12158 13626
rect 12182 13574 12212 13626
rect 12212 13574 12224 13626
rect 12224 13574 12238 13626
rect 12262 13574 12276 13626
rect 12276 13574 12288 13626
rect 12288 13574 12318 13626
rect 12342 13574 12352 13626
rect 12352 13574 12398 13626
rect 12102 13572 12158 13574
rect 12182 13572 12238 13574
rect 12262 13572 12318 13574
rect 12342 13572 12398 13574
rect 11442 13082 11498 13084
rect 11522 13082 11578 13084
rect 11602 13082 11658 13084
rect 11682 13082 11738 13084
rect 11442 13030 11488 13082
rect 11488 13030 11498 13082
rect 11522 13030 11552 13082
rect 11552 13030 11564 13082
rect 11564 13030 11578 13082
rect 11602 13030 11616 13082
rect 11616 13030 11628 13082
rect 11628 13030 11658 13082
rect 11682 13030 11692 13082
rect 11692 13030 11738 13082
rect 11442 13028 11498 13030
rect 11522 13028 11578 13030
rect 11602 13028 11658 13030
rect 11682 13028 11738 13030
rect 12102 12538 12158 12540
rect 12182 12538 12238 12540
rect 12262 12538 12318 12540
rect 12342 12538 12398 12540
rect 12102 12486 12148 12538
rect 12148 12486 12158 12538
rect 12182 12486 12212 12538
rect 12212 12486 12224 12538
rect 12224 12486 12238 12538
rect 12262 12486 12276 12538
rect 12276 12486 12288 12538
rect 12288 12486 12318 12538
rect 12342 12486 12352 12538
rect 12352 12486 12398 12538
rect 12102 12484 12158 12486
rect 12182 12484 12238 12486
rect 12262 12484 12318 12486
rect 12342 12484 12398 12486
rect 11442 11994 11498 11996
rect 11522 11994 11578 11996
rect 11602 11994 11658 11996
rect 11682 11994 11738 11996
rect 11442 11942 11488 11994
rect 11488 11942 11498 11994
rect 11522 11942 11552 11994
rect 11552 11942 11564 11994
rect 11564 11942 11578 11994
rect 11602 11942 11616 11994
rect 11616 11942 11628 11994
rect 11628 11942 11658 11994
rect 11682 11942 11692 11994
rect 11692 11942 11738 11994
rect 11442 11940 11498 11942
rect 11522 11940 11578 11942
rect 11602 11940 11658 11942
rect 11682 11940 11738 11942
rect 12898 17992 12954 18048
rect 14278 20476 14280 20496
rect 14280 20476 14332 20496
rect 14332 20476 14334 20496
rect 14278 20440 14334 20476
rect 14830 19624 14886 19680
rect 15198 20848 15254 20904
rect 16210 20712 16266 20768
rect 15474 20576 15530 20632
rect 16486 20596 16542 20632
rect 16486 20576 16488 20596
rect 16488 20576 16540 20596
rect 16540 20576 16542 20596
rect 15842 20304 15898 20360
rect 15014 19252 15016 19272
rect 15016 19252 15068 19272
rect 15068 19252 15070 19272
rect 15014 19216 15070 19252
rect 15566 20032 15622 20088
rect 14738 17992 14794 18048
rect 14278 17448 14334 17504
rect 12990 12688 13046 12744
rect 13726 13912 13782 13968
rect 13634 13776 13690 13832
rect 11442 10906 11498 10908
rect 11522 10906 11578 10908
rect 11602 10906 11658 10908
rect 11682 10906 11738 10908
rect 11442 10854 11488 10906
rect 11488 10854 11498 10906
rect 11522 10854 11552 10906
rect 11552 10854 11564 10906
rect 11564 10854 11578 10906
rect 11602 10854 11616 10906
rect 11616 10854 11628 10906
rect 11628 10854 11658 10906
rect 11682 10854 11692 10906
rect 11692 10854 11738 10906
rect 11442 10852 11498 10854
rect 11522 10852 11578 10854
rect 11602 10852 11658 10854
rect 11682 10852 11738 10854
rect 11442 9818 11498 9820
rect 11522 9818 11578 9820
rect 11602 9818 11658 9820
rect 11682 9818 11738 9820
rect 11442 9766 11488 9818
rect 11488 9766 11498 9818
rect 11522 9766 11552 9818
rect 11552 9766 11564 9818
rect 11564 9766 11578 9818
rect 11602 9766 11616 9818
rect 11616 9766 11628 9818
rect 11628 9766 11658 9818
rect 11682 9766 11692 9818
rect 11692 9766 11738 9818
rect 11442 9764 11498 9766
rect 11522 9764 11578 9766
rect 11602 9764 11658 9766
rect 11682 9764 11738 9766
rect 12102 11450 12158 11452
rect 12182 11450 12238 11452
rect 12262 11450 12318 11452
rect 12342 11450 12398 11452
rect 12102 11398 12148 11450
rect 12148 11398 12158 11450
rect 12182 11398 12212 11450
rect 12212 11398 12224 11450
rect 12224 11398 12238 11450
rect 12262 11398 12276 11450
rect 12276 11398 12288 11450
rect 12288 11398 12318 11450
rect 12342 11398 12352 11450
rect 12352 11398 12398 11450
rect 12102 11396 12158 11398
rect 12182 11396 12238 11398
rect 12262 11396 12318 11398
rect 12342 11396 12398 11398
rect 12102 10362 12158 10364
rect 12182 10362 12238 10364
rect 12262 10362 12318 10364
rect 12342 10362 12398 10364
rect 12102 10310 12148 10362
rect 12148 10310 12158 10362
rect 12182 10310 12212 10362
rect 12212 10310 12224 10362
rect 12224 10310 12238 10362
rect 12262 10310 12276 10362
rect 12276 10310 12288 10362
rect 12288 10310 12318 10362
rect 12342 10310 12352 10362
rect 12352 10310 12398 10362
rect 12102 10308 12158 10310
rect 12182 10308 12238 10310
rect 12262 10308 12318 10310
rect 12342 10308 12398 10310
rect 11442 8730 11498 8732
rect 11522 8730 11578 8732
rect 11602 8730 11658 8732
rect 11682 8730 11738 8732
rect 11442 8678 11488 8730
rect 11488 8678 11498 8730
rect 11522 8678 11552 8730
rect 11552 8678 11564 8730
rect 11564 8678 11578 8730
rect 11602 8678 11616 8730
rect 11616 8678 11628 8730
rect 11628 8678 11658 8730
rect 11682 8678 11692 8730
rect 11692 8678 11738 8730
rect 11442 8676 11498 8678
rect 11522 8676 11578 8678
rect 11602 8676 11658 8678
rect 11682 8676 11738 8678
rect 11442 7642 11498 7644
rect 11522 7642 11578 7644
rect 11602 7642 11658 7644
rect 11682 7642 11738 7644
rect 11442 7590 11488 7642
rect 11488 7590 11498 7642
rect 11522 7590 11552 7642
rect 11552 7590 11564 7642
rect 11564 7590 11578 7642
rect 11602 7590 11616 7642
rect 11616 7590 11628 7642
rect 11628 7590 11658 7642
rect 11682 7590 11692 7642
rect 11692 7590 11738 7642
rect 11442 7588 11498 7590
rect 11522 7588 11578 7590
rect 11602 7588 11658 7590
rect 11682 7588 11738 7590
rect 12102 9274 12158 9276
rect 12182 9274 12238 9276
rect 12262 9274 12318 9276
rect 12342 9274 12398 9276
rect 12102 9222 12148 9274
rect 12148 9222 12158 9274
rect 12182 9222 12212 9274
rect 12212 9222 12224 9274
rect 12224 9222 12238 9274
rect 12262 9222 12276 9274
rect 12276 9222 12288 9274
rect 12288 9222 12318 9274
rect 12342 9222 12352 9274
rect 12352 9222 12398 9274
rect 12102 9220 12158 9222
rect 12182 9220 12238 9222
rect 12262 9220 12318 9222
rect 12342 9220 12398 9222
rect 12102 8186 12158 8188
rect 12182 8186 12238 8188
rect 12262 8186 12318 8188
rect 12342 8186 12398 8188
rect 12102 8134 12148 8186
rect 12148 8134 12158 8186
rect 12182 8134 12212 8186
rect 12212 8134 12224 8186
rect 12224 8134 12238 8186
rect 12262 8134 12276 8186
rect 12276 8134 12288 8186
rect 12288 8134 12318 8186
rect 12342 8134 12352 8186
rect 12352 8134 12398 8186
rect 12102 8132 12158 8134
rect 12182 8132 12238 8134
rect 12262 8132 12318 8134
rect 12342 8132 12398 8134
rect 11442 6554 11498 6556
rect 11522 6554 11578 6556
rect 11602 6554 11658 6556
rect 11682 6554 11738 6556
rect 11442 6502 11488 6554
rect 11488 6502 11498 6554
rect 11522 6502 11552 6554
rect 11552 6502 11564 6554
rect 11564 6502 11578 6554
rect 11602 6502 11616 6554
rect 11616 6502 11628 6554
rect 11628 6502 11658 6554
rect 11682 6502 11692 6554
rect 11692 6502 11738 6554
rect 11442 6500 11498 6502
rect 11522 6500 11578 6502
rect 11602 6500 11658 6502
rect 11682 6500 11738 6502
rect 12102 7098 12158 7100
rect 12182 7098 12238 7100
rect 12262 7098 12318 7100
rect 12342 7098 12398 7100
rect 12102 7046 12148 7098
rect 12148 7046 12158 7098
rect 12182 7046 12212 7098
rect 12212 7046 12224 7098
rect 12224 7046 12238 7098
rect 12262 7046 12276 7098
rect 12276 7046 12288 7098
rect 12288 7046 12318 7098
rect 12342 7046 12352 7098
rect 12352 7046 12398 7098
rect 12102 7044 12158 7046
rect 12182 7044 12238 7046
rect 12262 7044 12318 7046
rect 12342 7044 12398 7046
rect 15198 18264 15254 18320
rect 15014 18148 15070 18184
rect 15014 18128 15016 18148
rect 15016 18128 15068 18148
rect 15068 18128 15070 18148
rect 15014 14320 15070 14376
rect 15106 12824 15162 12880
rect 15566 12280 15622 12336
rect 15014 10124 15070 10160
rect 15014 10104 15016 10124
rect 15016 10104 15068 10124
rect 15068 10104 15070 10124
rect 14002 7928 14058 7984
rect 15014 8084 15070 8120
rect 15014 8064 15016 8084
rect 15016 8064 15068 8084
rect 15068 8064 15070 8084
rect 14554 7928 14610 7984
rect 11442 5466 11498 5468
rect 11522 5466 11578 5468
rect 11602 5466 11658 5468
rect 11682 5466 11738 5468
rect 11442 5414 11488 5466
rect 11488 5414 11498 5466
rect 11522 5414 11552 5466
rect 11552 5414 11564 5466
rect 11564 5414 11578 5466
rect 11602 5414 11616 5466
rect 11616 5414 11628 5466
rect 11628 5414 11658 5466
rect 11682 5414 11692 5466
rect 11692 5414 11738 5466
rect 11442 5412 11498 5414
rect 11522 5412 11578 5414
rect 11602 5412 11658 5414
rect 11682 5412 11738 5414
rect 12102 6010 12158 6012
rect 12182 6010 12238 6012
rect 12262 6010 12318 6012
rect 12342 6010 12398 6012
rect 12102 5958 12148 6010
rect 12148 5958 12158 6010
rect 12182 5958 12212 6010
rect 12212 5958 12224 6010
rect 12224 5958 12238 6010
rect 12262 5958 12276 6010
rect 12276 5958 12288 6010
rect 12288 5958 12318 6010
rect 12342 5958 12352 6010
rect 12352 5958 12398 6010
rect 12102 5956 12158 5958
rect 12182 5956 12238 5958
rect 12262 5956 12318 5958
rect 12342 5956 12398 5958
rect 12530 5364 12586 5400
rect 12530 5344 12532 5364
rect 12532 5344 12584 5364
rect 12584 5344 12586 5364
rect 11442 4378 11498 4380
rect 11522 4378 11578 4380
rect 11602 4378 11658 4380
rect 11682 4378 11738 4380
rect 11442 4326 11488 4378
rect 11488 4326 11498 4378
rect 11522 4326 11552 4378
rect 11552 4326 11564 4378
rect 11564 4326 11578 4378
rect 11602 4326 11616 4378
rect 11616 4326 11628 4378
rect 11628 4326 11658 4378
rect 11682 4326 11692 4378
rect 11692 4326 11738 4378
rect 11442 4324 11498 4326
rect 11522 4324 11578 4326
rect 11602 4324 11658 4326
rect 11682 4324 11738 4326
rect 12102 4922 12158 4924
rect 12182 4922 12238 4924
rect 12262 4922 12318 4924
rect 12342 4922 12398 4924
rect 12102 4870 12148 4922
rect 12148 4870 12158 4922
rect 12182 4870 12212 4922
rect 12212 4870 12224 4922
rect 12224 4870 12238 4922
rect 12262 4870 12276 4922
rect 12276 4870 12288 4922
rect 12288 4870 12318 4922
rect 12342 4870 12352 4922
rect 12352 4870 12398 4922
rect 12102 4868 12158 4870
rect 12182 4868 12238 4870
rect 12262 4868 12318 4870
rect 12342 4868 12398 4870
rect 16118 18264 16174 18320
rect 16118 17740 16174 17776
rect 16118 17720 16120 17740
rect 16120 17720 16172 17740
rect 16172 17720 16174 17740
rect 17222 19236 17278 19272
rect 17222 19216 17224 19236
rect 17224 19216 17276 19236
rect 17276 19216 17278 19236
rect 16486 15408 16542 15464
rect 16578 14456 16634 14512
rect 15658 8064 15714 8120
rect 15566 7948 15622 7984
rect 15566 7928 15568 7948
rect 15568 7928 15620 7948
rect 15620 7928 15622 7948
rect 14554 4120 14610 4176
rect 12102 3834 12158 3836
rect 12182 3834 12238 3836
rect 12262 3834 12318 3836
rect 12342 3834 12398 3836
rect 12102 3782 12148 3834
rect 12148 3782 12158 3834
rect 12182 3782 12212 3834
rect 12212 3782 12224 3834
rect 12224 3782 12238 3834
rect 12262 3782 12276 3834
rect 12276 3782 12288 3834
rect 12288 3782 12318 3834
rect 12342 3782 12352 3834
rect 12352 3782 12398 3834
rect 12102 3780 12158 3782
rect 12182 3780 12238 3782
rect 12262 3780 12318 3782
rect 12342 3780 12398 3782
rect 11442 3290 11498 3292
rect 11522 3290 11578 3292
rect 11602 3290 11658 3292
rect 11682 3290 11738 3292
rect 11442 3238 11488 3290
rect 11488 3238 11498 3290
rect 11522 3238 11552 3290
rect 11552 3238 11564 3290
rect 11564 3238 11578 3290
rect 11602 3238 11616 3290
rect 11616 3238 11628 3290
rect 11628 3238 11658 3290
rect 11682 3238 11692 3290
rect 11692 3238 11738 3290
rect 11442 3236 11498 3238
rect 11522 3236 11578 3238
rect 11602 3236 11658 3238
rect 11682 3236 11738 3238
rect 12102 2746 12158 2748
rect 12182 2746 12238 2748
rect 12262 2746 12318 2748
rect 12342 2746 12398 2748
rect 12102 2694 12148 2746
rect 12148 2694 12158 2746
rect 12182 2694 12212 2746
rect 12212 2694 12224 2746
rect 12224 2694 12238 2746
rect 12262 2694 12276 2746
rect 12276 2694 12288 2746
rect 12288 2694 12318 2746
rect 12342 2694 12352 2746
rect 12352 2694 12398 2746
rect 12102 2692 12158 2694
rect 12182 2692 12238 2694
rect 12262 2692 12318 2694
rect 12342 2692 12398 2694
rect 11442 2202 11498 2204
rect 11522 2202 11578 2204
rect 11602 2202 11658 2204
rect 11682 2202 11738 2204
rect 11442 2150 11488 2202
rect 11488 2150 11498 2202
rect 11522 2150 11552 2202
rect 11552 2150 11564 2202
rect 11564 2150 11578 2202
rect 11602 2150 11616 2202
rect 11616 2150 11628 2202
rect 11628 2150 11658 2202
rect 11682 2150 11692 2202
rect 11692 2150 11738 2202
rect 11442 2148 11498 2150
rect 11522 2148 11578 2150
rect 11602 2148 11658 2150
rect 11682 2148 11738 2150
rect 12102 1658 12158 1660
rect 12182 1658 12238 1660
rect 12262 1658 12318 1660
rect 12342 1658 12398 1660
rect 12102 1606 12148 1658
rect 12148 1606 12158 1658
rect 12182 1606 12212 1658
rect 12212 1606 12224 1658
rect 12224 1606 12238 1658
rect 12262 1606 12276 1658
rect 12276 1606 12288 1658
rect 12288 1606 12318 1658
rect 12342 1606 12352 1658
rect 12352 1606 12398 1658
rect 12102 1604 12158 1606
rect 12182 1604 12238 1606
rect 12262 1604 12318 1606
rect 12342 1604 12398 1606
rect 17222 15000 17278 15056
rect 17958 19916 18014 19952
rect 17958 19896 17960 19916
rect 17960 19896 18012 19916
rect 18012 19896 18014 19916
rect 18050 19760 18106 19816
rect 19522 21004 19578 21040
rect 19522 20984 19524 21004
rect 19524 20984 19576 21004
rect 19576 20984 19578 21004
rect 18970 20440 19026 20496
rect 19216 20698 19272 20700
rect 19296 20698 19352 20700
rect 19376 20698 19432 20700
rect 19456 20698 19512 20700
rect 19216 20646 19262 20698
rect 19262 20646 19272 20698
rect 19296 20646 19326 20698
rect 19326 20646 19338 20698
rect 19338 20646 19352 20698
rect 19376 20646 19390 20698
rect 19390 20646 19402 20698
rect 19402 20646 19432 20698
rect 19456 20646 19466 20698
rect 19466 20646 19512 20698
rect 19216 20644 19272 20646
rect 19296 20644 19352 20646
rect 19376 20644 19432 20646
rect 19456 20644 19512 20646
rect 18786 20304 18842 20360
rect 18326 17992 18382 18048
rect 17314 14456 17370 14512
rect 18878 19624 18934 19680
rect 19876 21242 19932 21244
rect 19956 21242 20012 21244
rect 20036 21242 20092 21244
rect 20116 21242 20172 21244
rect 19876 21190 19922 21242
rect 19922 21190 19932 21242
rect 19956 21190 19986 21242
rect 19986 21190 19998 21242
rect 19998 21190 20012 21242
rect 20036 21190 20050 21242
rect 20050 21190 20062 21242
rect 20062 21190 20092 21242
rect 20116 21190 20126 21242
rect 20126 21190 20172 21242
rect 19876 21188 19932 21190
rect 19956 21188 20012 21190
rect 20036 21188 20092 21190
rect 20116 21188 20172 21190
rect 19706 21120 19762 21176
rect 18602 17584 18658 17640
rect 18326 15428 18382 15464
rect 18326 15408 18328 15428
rect 18328 15408 18380 15428
rect 18380 15408 18382 15428
rect 19338 19760 19394 19816
rect 19216 19610 19272 19612
rect 19296 19610 19352 19612
rect 19376 19610 19432 19612
rect 19456 19610 19512 19612
rect 19216 19558 19262 19610
rect 19262 19558 19272 19610
rect 19296 19558 19326 19610
rect 19326 19558 19338 19610
rect 19338 19558 19352 19610
rect 19376 19558 19390 19610
rect 19390 19558 19402 19610
rect 19402 19558 19432 19610
rect 19456 19558 19466 19610
rect 19466 19558 19512 19610
rect 19216 19556 19272 19558
rect 19296 19556 19352 19558
rect 19376 19556 19432 19558
rect 19456 19556 19512 19558
rect 19216 18522 19272 18524
rect 19296 18522 19352 18524
rect 19376 18522 19432 18524
rect 19456 18522 19512 18524
rect 19216 18470 19262 18522
rect 19262 18470 19272 18522
rect 19296 18470 19326 18522
rect 19326 18470 19338 18522
rect 19338 18470 19352 18522
rect 19376 18470 19390 18522
rect 19390 18470 19402 18522
rect 19402 18470 19432 18522
rect 19456 18470 19466 18522
rect 19466 18470 19512 18522
rect 19216 18468 19272 18470
rect 19296 18468 19352 18470
rect 19376 18468 19432 18470
rect 19456 18468 19512 18470
rect 19246 17992 19302 18048
rect 20902 20440 20958 20496
rect 21546 20440 21602 20496
rect 19876 20154 19932 20156
rect 19956 20154 20012 20156
rect 20036 20154 20092 20156
rect 20116 20154 20172 20156
rect 19876 20102 19922 20154
rect 19922 20102 19932 20154
rect 19956 20102 19986 20154
rect 19986 20102 19998 20154
rect 19998 20102 20012 20154
rect 20036 20102 20050 20154
rect 20050 20102 20062 20154
rect 20062 20102 20092 20154
rect 20116 20102 20126 20154
rect 20126 20102 20172 20154
rect 19876 20100 19932 20102
rect 19956 20100 20012 20102
rect 20036 20100 20092 20102
rect 20116 20100 20172 20102
rect 19876 19066 19932 19068
rect 19956 19066 20012 19068
rect 20036 19066 20092 19068
rect 20116 19066 20172 19068
rect 19876 19014 19922 19066
rect 19922 19014 19932 19066
rect 19956 19014 19986 19066
rect 19986 19014 19998 19066
rect 19998 19014 20012 19066
rect 20036 19014 20050 19066
rect 20050 19014 20062 19066
rect 20062 19014 20092 19066
rect 20116 19014 20126 19066
rect 20126 19014 20172 19066
rect 19876 19012 19932 19014
rect 19956 19012 20012 19014
rect 20036 19012 20092 19014
rect 20116 19012 20172 19014
rect 18970 17448 19026 17504
rect 19216 17434 19272 17436
rect 19296 17434 19352 17436
rect 19376 17434 19432 17436
rect 19456 17434 19512 17436
rect 19216 17382 19262 17434
rect 19262 17382 19272 17434
rect 19296 17382 19326 17434
rect 19326 17382 19338 17434
rect 19338 17382 19352 17434
rect 19376 17382 19390 17434
rect 19390 17382 19402 17434
rect 19402 17382 19432 17434
rect 19456 17382 19466 17434
rect 19466 17382 19512 17434
rect 19216 17380 19272 17382
rect 19296 17380 19352 17382
rect 19376 17380 19432 17382
rect 19456 17380 19512 17382
rect 19216 16346 19272 16348
rect 19296 16346 19352 16348
rect 19376 16346 19432 16348
rect 19456 16346 19512 16348
rect 19216 16294 19262 16346
rect 19262 16294 19272 16346
rect 19296 16294 19326 16346
rect 19326 16294 19338 16346
rect 19338 16294 19352 16346
rect 19376 16294 19390 16346
rect 19390 16294 19402 16346
rect 19402 16294 19432 16346
rect 19456 16294 19466 16346
rect 19466 16294 19512 16346
rect 19216 16292 19272 16294
rect 19296 16292 19352 16294
rect 19376 16292 19432 16294
rect 19456 16292 19512 16294
rect 19876 17978 19932 17980
rect 19956 17978 20012 17980
rect 20036 17978 20092 17980
rect 20116 17978 20172 17980
rect 19876 17926 19922 17978
rect 19922 17926 19932 17978
rect 19956 17926 19986 17978
rect 19986 17926 19998 17978
rect 19998 17926 20012 17978
rect 20036 17926 20050 17978
rect 20050 17926 20062 17978
rect 20062 17926 20092 17978
rect 20116 17926 20126 17978
rect 20126 17926 20172 17978
rect 19876 17924 19932 17926
rect 19956 17924 20012 17926
rect 20036 17924 20092 17926
rect 20116 17924 20172 17926
rect 20258 17212 20260 17232
rect 20260 17212 20312 17232
rect 20312 17212 20314 17232
rect 20258 17176 20314 17212
rect 19876 16890 19932 16892
rect 19956 16890 20012 16892
rect 20036 16890 20092 16892
rect 20116 16890 20172 16892
rect 19876 16838 19922 16890
rect 19922 16838 19932 16890
rect 19956 16838 19986 16890
rect 19986 16838 19998 16890
rect 19998 16838 20012 16890
rect 20036 16838 20050 16890
rect 20050 16838 20062 16890
rect 20062 16838 20092 16890
rect 20116 16838 20126 16890
rect 20126 16838 20172 16890
rect 19876 16836 19932 16838
rect 19956 16836 20012 16838
rect 20036 16836 20092 16838
rect 20116 16836 20172 16838
rect 19216 15258 19272 15260
rect 19296 15258 19352 15260
rect 19376 15258 19432 15260
rect 19456 15258 19512 15260
rect 19216 15206 19262 15258
rect 19262 15206 19272 15258
rect 19296 15206 19326 15258
rect 19326 15206 19338 15258
rect 19338 15206 19352 15258
rect 19376 15206 19390 15258
rect 19390 15206 19402 15258
rect 19402 15206 19432 15258
rect 19456 15206 19466 15258
rect 19466 15206 19512 15258
rect 19216 15204 19272 15206
rect 19296 15204 19352 15206
rect 19376 15204 19432 15206
rect 19456 15204 19512 15206
rect 18786 14900 18788 14920
rect 18788 14900 18840 14920
rect 18840 14900 18842 14920
rect 18786 14864 18842 14900
rect 18050 14320 18106 14376
rect 17314 12724 17316 12744
rect 17316 12724 17368 12744
rect 17368 12724 17370 12744
rect 17314 12688 17370 12724
rect 16946 10140 16948 10160
rect 16948 10140 17000 10160
rect 17000 10140 17002 10160
rect 16946 10104 17002 10140
rect 16854 7964 16856 7984
rect 16856 7964 16908 7984
rect 16908 7964 16910 7984
rect 16854 7928 16910 7964
rect 15934 5616 15990 5672
rect 17590 8064 17646 8120
rect 18142 12860 18144 12880
rect 18144 12860 18196 12880
rect 18196 12860 18198 12880
rect 18142 12824 18198 12860
rect 19216 14170 19272 14172
rect 19296 14170 19352 14172
rect 19376 14170 19432 14172
rect 19456 14170 19512 14172
rect 19216 14118 19262 14170
rect 19262 14118 19272 14170
rect 19296 14118 19326 14170
rect 19326 14118 19338 14170
rect 19338 14118 19352 14170
rect 19376 14118 19390 14170
rect 19390 14118 19402 14170
rect 19402 14118 19432 14170
rect 19456 14118 19466 14170
rect 19466 14118 19512 14170
rect 19216 14116 19272 14118
rect 19296 14116 19352 14118
rect 19376 14116 19432 14118
rect 19456 14116 19512 14118
rect 19430 13776 19486 13832
rect 19216 13082 19272 13084
rect 19296 13082 19352 13084
rect 19376 13082 19432 13084
rect 19456 13082 19512 13084
rect 19216 13030 19262 13082
rect 19262 13030 19272 13082
rect 19296 13030 19326 13082
rect 19326 13030 19338 13082
rect 19338 13030 19352 13082
rect 19376 13030 19390 13082
rect 19390 13030 19402 13082
rect 19402 13030 19432 13082
rect 19456 13030 19466 13082
rect 19466 13030 19512 13082
rect 19216 13028 19272 13030
rect 19296 13028 19352 13030
rect 19376 13028 19432 13030
rect 19456 13028 19512 13030
rect 19614 12280 19670 12336
rect 17866 11620 17922 11656
rect 17866 11600 17868 11620
rect 17868 11600 17920 11620
rect 17920 11600 17922 11620
rect 19216 11994 19272 11996
rect 19296 11994 19352 11996
rect 19376 11994 19432 11996
rect 19456 11994 19512 11996
rect 19216 11942 19262 11994
rect 19262 11942 19272 11994
rect 19296 11942 19326 11994
rect 19326 11942 19338 11994
rect 19338 11942 19352 11994
rect 19376 11942 19390 11994
rect 19390 11942 19402 11994
rect 19402 11942 19432 11994
rect 19456 11942 19466 11994
rect 19466 11942 19512 11994
rect 19216 11940 19272 11942
rect 19296 11940 19352 11942
rect 19376 11940 19432 11942
rect 19456 11940 19512 11942
rect 19876 15802 19932 15804
rect 19956 15802 20012 15804
rect 20036 15802 20092 15804
rect 20116 15802 20172 15804
rect 19876 15750 19922 15802
rect 19922 15750 19932 15802
rect 19956 15750 19986 15802
rect 19986 15750 19998 15802
rect 19998 15750 20012 15802
rect 20036 15750 20050 15802
rect 20050 15750 20062 15802
rect 20062 15750 20092 15802
rect 20116 15750 20126 15802
rect 20126 15750 20172 15802
rect 19876 15748 19932 15750
rect 19956 15748 20012 15750
rect 20036 15748 20092 15750
rect 20116 15748 20172 15750
rect 19876 14714 19932 14716
rect 19956 14714 20012 14716
rect 20036 14714 20092 14716
rect 20116 14714 20172 14716
rect 19876 14662 19922 14714
rect 19922 14662 19932 14714
rect 19956 14662 19986 14714
rect 19986 14662 19998 14714
rect 19998 14662 20012 14714
rect 20036 14662 20050 14714
rect 20050 14662 20062 14714
rect 20062 14662 20092 14714
rect 20116 14662 20126 14714
rect 20126 14662 20172 14714
rect 19876 14660 19932 14662
rect 19956 14660 20012 14662
rect 20036 14660 20092 14662
rect 20116 14660 20172 14662
rect 19890 13948 19892 13968
rect 19892 13948 19944 13968
rect 19944 13948 19946 13968
rect 19890 13912 19946 13948
rect 19876 13626 19932 13628
rect 19956 13626 20012 13628
rect 20036 13626 20092 13628
rect 20116 13626 20172 13628
rect 19876 13574 19922 13626
rect 19922 13574 19932 13626
rect 19956 13574 19986 13626
rect 19986 13574 19998 13626
rect 19998 13574 20012 13626
rect 20036 13574 20050 13626
rect 20050 13574 20062 13626
rect 20062 13574 20092 13626
rect 20116 13574 20126 13626
rect 20126 13574 20172 13626
rect 19876 13572 19932 13574
rect 19956 13572 20012 13574
rect 20036 13572 20092 13574
rect 20116 13572 20172 13574
rect 20534 13776 20590 13832
rect 26422 21800 26478 21856
rect 26698 21800 26754 21856
rect 25318 21664 25374 21720
rect 22466 20052 22522 20088
rect 22466 20032 22468 20052
rect 22468 20032 22520 20052
rect 22520 20032 22522 20052
rect 24030 18708 24032 18728
rect 24032 18708 24084 18728
rect 24084 18708 24086 18728
rect 24030 18672 24086 18708
rect 21454 17856 21510 17912
rect 21270 15564 21326 15600
rect 21270 15544 21272 15564
rect 21272 15544 21324 15564
rect 21324 15544 21326 15564
rect 22190 17448 22246 17504
rect 22006 15988 22008 16008
rect 22008 15988 22060 16008
rect 22060 15988 22062 16008
rect 22006 15952 22062 15988
rect 21086 15444 21088 15464
rect 21088 15444 21140 15464
rect 21140 15444 21142 15464
rect 21086 15408 21142 15444
rect 21362 15000 21418 15056
rect 21730 14048 21786 14104
rect 21730 13776 21786 13832
rect 19876 12538 19932 12540
rect 19956 12538 20012 12540
rect 20036 12538 20092 12540
rect 20116 12538 20172 12540
rect 19876 12486 19922 12538
rect 19922 12486 19932 12538
rect 19956 12486 19986 12538
rect 19986 12486 19998 12538
rect 19998 12486 20012 12538
rect 20036 12486 20050 12538
rect 20050 12486 20062 12538
rect 20062 12486 20092 12538
rect 20116 12486 20126 12538
rect 20126 12486 20172 12538
rect 19876 12484 19932 12486
rect 19956 12484 20012 12486
rect 20036 12484 20092 12486
rect 20116 12484 20172 12486
rect 19338 11076 19394 11112
rect 19338 11056 19340 11076
rect 19340 11056 19392 11076
rect 19392 11056 19394 11076
rect 19876 11450 19932 11452
rect 19956 11450 20012 11452
rect 20036 11450 20092 11452
rect 20116 11450 20172 11452
rect 19876 11398 19922 11450
rect 19922 11398 19932 11450
rect 19956 11398 19986 11450
rect 19986 11398 19998 11450
rect 19998 11398 20012 11450
rect 20036 11398 20050 11450
rect 20050 11398 20062 11450
rect 20062 11398 20092 11450
rect 20116 11398 20126 11450
rect 20126 11398 20172 11450
rect 19876 11396 19932 11398
rect 19956 11396 20012 11398
rect 20036 11396 20092 11398
rect 20116 11396 20172 11398
rect 19216 10906 19272 10908
rect 19296 10906 19352 10908
rect 19376 10906 19432 10908
rect 19456 10906 19512 10908
rect 19216 10854 19262 10906
rect 19262 10854 19272 10906
rect 19296 10854 19326 10906
rect 19326 10854 19338 10906
rect 19338 10854 19352 10906
rect 19376 10854 19390 10906
rect 19390 10854 19402 10906
rect 19402 10854 19432 10906
rect 19456 10854 19466 10906
rect 19466 10854 19512 10906
rect 19216 10852 19272 10854
rect 19296 10852 19352 10854
rect 19376 10852 19432 10854
rect 19456 10852 19512 10854
rect 19216 9818 19272 9820
rect 19296 9818 19352 9820
rect 19376 9818 19432 9820
rect 19456 9818 19512 9820
rect 19216 9766 19262 9818
rect 19262 9766 19272 9818
rect 19296 9766 19326 9818
rect 19326 9766 19338 9818
rect 19338 9766 19352 9818
rect 19376 9766 19390 9818
rect 19390 9766 19402 9818
rect 19402 9766 19432 9818
rect 19456 9766 19466 9818
rect 19466 9766 19512 9818
rect 19216 9764 19272 9766
rect 19296 9764 19352 9766
rect 19376 9764 19432 9766
rect 19456 9764 19512 9766
rect 19338 9444 19394 9480
rect 19338 9424 19340 9444
rect 19340 9424 19392 9444
rect 19392 9424 19394 9444
rect 19216 8730 19272 8732
rect 19296 8730 19352 8732
rect 19376 8730 19432 8732
rect 19456 8730 19512 8732
rect 19216 8678 19262 8730
rect 19262 8678 19272 8730
rect 19296 8678 19326 8730
rect 19326 8678 19338 8730
rect 19338 8678 19352 8730
rect 19376 8678 19390 8730
rect 19390 8678 19402 8730
rect 19402 8678 19432 8730
rect 19456 8678 19466 8730
rect 19466 8678 19512 8730
rect 19216 8676 19272 8678
rect 19296 8676 19352 8678
rect 19376 8676 19432 8678
rect 19456 8676 19512 8678
rect 19982 11212 20038 11248
rect 20442 12164 20498 12200
rect 20442 12144 20444 12164
rect 20444 12144 20496 12164
rect 20496 12144 20498 12164
rect 19982 11192 19984 11212
rect 19984 11192 20036 11212
rect 20036 11192 20038 11212
rect 19876 10362 19932 10364
rect 19956 10362 20012 10364
rect 20036 10362 20092 10364
rect 20116 10362 20172 10364
rect 19876 10310 19922 10362
rect 19922 10310 19932 10362
rect 19956 10310 19986 10362
rect 19986 10310 19998 10362
rect 19998 10310 20012 10362
rect 20036 10310 20050 10362
rect 20050 10310 20062 10362
rect 20062 10310 20092 10362
rect 20116 10310 20126 10362
rect 20126 10310 20172 10362
rect 19876 10308 19932 10310
rect 19956 10308 20012 10310
rect 20036 10308 20092 10310
rect 20116 10308 20172 10310
rect 19876 9274 19932 9276
rect 19956 9274 20012 9276
rect 20036 9274 20092 9276
rect 20116 9274 20172 9276
rect 19876 9222 19922 9274
rect 19922 9222 19932 9274
rect 19956 9222 19986 9274
rect 19986 9222 19998 9274
rect 19998 9222 20012 9274
rect 20036 9222 20050 9274
rect 20050 9222 20062 9274
rect 20062 9222 20092 9274
rect 20116 9222 20126 9274
rect 20126 9222 20172 9274
rect 19876 9220 19932 9222
rect 19956 9220 20012 9222
rect 20036 9220 20092 9222
rect 20116 9220 20172 9222
rect 19876 8186 19932 8188
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 19876 8134 19922 8186
rect 19922 8134 19932 8186
rect 19956 8134 19986 8186
rect 19986 8134 19998 8186
rect 19998 8134 20012 8186
rect 20036 8134 20050 8186
rect 20050 8134 20062 8186
rect 20062 8134 20092 8186
rect 20116 8134 20126 8186
rect 20126 8134 20172 8186
rect 19876 8132 19932 8134
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 18142 6180 18198 6216
rect 18142 6160 18144 6180
rect 18144 6160 18196 6180
rect 18196 6160 18198 6180
rect 20534 9444 20590 9480
rect 20534 9424 20536 9444
rect 20536 9424 20588 9444
rect 20588 9424 20590 9444
rect 19216 7642 19272 7644
rect 19296 7642 19352 7644
rect 19376 7642 19432 7644
rect 19456 7642 19512 7644
rect 19216 7590 19262 7642
rect 19262 7590 19272 7642
rect 19296 7590 19326 7642
rect 19326 7590 19338 7642
rect 19338 7590 19352 7642
rect 19376 7590 19390 7642
rect 19390 7590 19402 7642
rect 19402 7590 19432 7642
rect 19456 7590 19466 7642
rect 19466 7590 19512 7642
rect 19216 7588 19272 7590
rect 19296 7588 19352 7590
rect 19376 7588 19432 7590
rect 19456 7588 19512 7590
rect 19154 6976 19210 7032
rect 19246 6860 19302 6896
rect 19876 7098 19932 7100
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 19876 7046 19922 7098
rect 19922 7046 19932 7098
rect 19956 7046 19986 7098
rect 19986 7046 19998 7098
rect 19998 7046 20012 7098
rect 20036 7046 20050 7098
rect 20050 7046 20062 7098
rect 20062 7046 20092 7098
rect 20116 7046 20126 7098
rect 20126 7046 20172 7098
rect 19876 7044 19932 7046
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 19246 6840 19248 6860
rect 19248 6840 19300 6860
rect 19300 6840 19302 6860
rect 18970 6704 19026 6760
rect 19216 6554 19272 6556
rect 19296 6554 19352 6556
rect 19376 6554 19432 6556
rect 19456 6554 19512 6556
rect 19216 6502 19262 6554
rect 19262 6502 19272 6554
rect 19296 6502 19326 6554
rect 19326 6502 19338 6554
rect 19338 6502 19352 6554
rect 19376 6502 19390 6554
rect 19390 6502 19402 6554
rect 19402 6502 19432 6554
rect 19456 6502 19466 6554
rect 19466 6502 19512 6554
rect 19216 6500 19272 6502
rect 19296 6500 19352 6502
rect 19376 6500 19432 6502
rect 19456 6500 19512 6502
rect 19154 6296 19210 6352
rect 19982 6296 20038 6352
rect 18970 6024 19026 6080
rect 18234 4120 18290 4176
rect 19062 5888 19118 5944
rect 18970 5344 19026 5400
rect 19338 6024 19394 6080
rect 19798 6160 19854 6216
rect 19876 6010 19932 6012
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 19876 5958 19922 6010
rect 19922 5958 19932 6010
rect 19956 5958 19986 6010
rect 19986 5958 19998 6010
rect 19998 5958 20012 6010
rect 20036 5958 20050 6010
rect 20050 5958 20062 6010
rect 20062 5958 20092 6010
rect 20116 5958 20126 6010
rect 20126 5958 20172 6010
rect 19876 5956 19932 5958
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 19706 5752 19762 5808
rect 19216 5466 19272 5468
rect 19296 5466 19352 5468
rect 19376 5466 19432 5468
rect 19456 5466 19512 5468
rect 19216 5414 19262 5466
rect 19262 5414 19272 5466
rect 19296 5414 19326 5466
rect 19326 5414 19338 5466
rect 19338 5414 19352 5466
rect 19376 5414 19390 5466
rect 19390 5414 19402 5466
rect 19402 5414 19432 5466
rect 19456 5414 19466 5466
rect 19466 5414 19512 5466
rect 19216 5412 19272 5414
rect 19296 5412 19352 5414
rect 19376 5412 19432 5414
rect 19456 5412 19512 5414
rect 19216 4378 19272 4380
rect 19296 4378 19352 4380
rect 19376 4378 19432 4380
rect 19456 4378 19512 4380
rect 19216 4326 19262 4378
rect 19262 4326 19272 4378
rect 19296 4326 19326 4378
rect 19326 4326 19338 4378
rect 19338 4326 19352 4378
rect 19376 4326 19390 4378
rect 19390 4326 19402 4378
rect 19402 4326 19432 4378
rect 19456 4326 19466 4378
rect 19466 4326 19512 4378
rect 19216 4324 19272 4326
rect 19296 4324 19352 4326
rect 19376 4324 19432 4326
rect 19456 4324 19512 4326
rect 19216 3290 19272 3292
rect 19296 3290 19352 3292
rect 19376 3290 19432 3292
rect 19456 3290 19512 3292
rect 19216 3238 19262 3290
rect 19262 3238 19272 3290
rect 19296 3238 19326 3290
rect 19326 3238 19338 3290
rect 19338 3238 19352 3290
rect 19376 3238 19390 3290
rect 19390 3238 19402 3290
rect 19402 3238 19432 3290
rect 19456 3238 19466 3290
rect 19466 3238 19512 3290
rect 19216 3236 19272 3238
rect 19296 3236 19352 3238
rect 19376 3236 19432 3238
rect 19456 3236 19512 3238
rect 11442 1114 11498 1116
rect 11522 1114 11578 1116
rect 11602 1114 11658 1116
rect 11682 1114 11738 1116
rect 11442 1062 11488 1114
rect 11488 1062 11498 1114
rect 11522 1062 11552 1114
rect 11552 1062 11564 1114
rect 11564 1062 11578 1114
rect 11602 1062 11616 1114
rect 11616 1062 11628 1114
rect 11628 1062 11658 1114
rect 11682 1062 11692 1114
rect 11692 1062 11738 1114
rect 11442 1060 11498 1062
rect 11522 1060 11578 1062
rect 11602 1060 11658 1062
rect 11682 1060 11738 1062
rect 20626 5480 20682 5536
rect 19876 4922 19932 4924
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 19876 4870 19922 4922
rect 19922 4870 19932 4922
rect 19956 4870 19986 4922
rect 19986 4870 19998 4922
rect 19998 4870 20012 4922
rect 20036 4870 20050 4922
rect 20050 4870 20062 4922
rect 20062 4870 20092 4922
rect 20116 4870 20126 4922
rect 20126 4870 20172 4922
rect 19876 4868 19932 4870
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 19876 3834 19932 3836
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 19876 3782 19922 3834
rect 19922 3782 19932 3834
rect 19956 3782 19986 3834
rect 19986 3782 19998 3834
rect 19998 3782 20012 3834
rect 20036 3782 20050 3834
rect 20050 3782 20062 3834
rect 20062 3782 20092 3834
rect 20116 3782 20126 3834
rect 20126 3782 20172 3834
rect 19876 3780 19932 3782
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 21178 5344 21234 5400
rect 21362 5208 21418 5264
rect 22282 14184 22338 14240
rect 23018 15816 23074 15872
rect 22926 15408 22982 15464
rect 23938 15564 23994 15600
rect 23938 15544 23940 15564
rect 23940 15544 23992 15564
rect 23992 15544 23994 15564
rect 24030 15000 24086 15056
rect 24214 15816 24270 15872
rect 22926 13776 22982 13832
rect 23386 13812 23388 13832
rect 23388 13812 23440 13832
rect 23440 13812 23442 13832
rect 23386 13776 23442 13812
rect 25502 21528 25558 21584
rect 26990 21786 27046 21788
rect 27070 21786 27126 21788
rect 27150 21786 27206 21788
rect 27230 21786 27286 21788
rect 26990 21734 27036 21786
rect 27036 21734 27046 21786
rect 27070 21734 27100 21786
rect 27100 21734 27112 21786
rect 27112 21734 27126 21786
rect 27150 21734 27164 21786
rect 27164 21734 27176 21786
rect 27176 21734 27206 21786
rect 27230 21734 27240 21786
rect 27240 21734 27286 21786
rect 26990 21732 27046 21734
rect 27070 21732 27126 21734
rect 27150 21732 27206 21734
rect 27230 21732 27286 21734
rect 28262 21800 28318 21856
rect 25134 19352 25190 19408
rect 27650 21242 27706 21244
rect 27730 21242 27786 21244
rect 27810 21242 27866 21244
rect 27890 21242 27946 21244
rect 27650 21190 27696 21242
rect 27696 21190 27706 21242
rect 27730 21190 27760 21242
rect 27760 21190 27772 21242
rect 27772 21190 27786 21242
rect 27810 21190 27824 21242
rect 27824 21190 27836 21242
rect 27836 21190 27866 21242
rect 27890 21190 27900 21242
rect 27900 21190 27946 21242
rect 27650 21188 27706 21190
rect 27730 21188 27786 21190
rect 27810 21188 27866 21190
rect 27890 21188 27946 21190
rect 26990 20698 27046 20700
rect 27070 20698 27126 20700
rect 27150 20698 27206 20700
rect 27230 20698 27286 20700
rect 26990 20646 27036 20698
rect 27036 20646 27046 20698
rect 27070 20646 27100 20698
rect 27100 20646 27112 20698
rect 27112 20646 27126 20698
rect 27150 20646 27164 20698
rect 27164 20646 27176 20698
rect 27176 20646 27206 20698
rect 27230 20646 27240 20698
rect 27240 20646 27286 20698
rect 26990 20644 27046 20646
rect 27070 20644 27126 20646
rect 27150 20644 27206 20646
rect 27230 20644 27286 20646
rect 26514 20032 26570 20088
rect 25134 18128 25190 18184
rect 24674 17584 24730 17640
rect 25226 17856 25282 17912
rect 24306 14320 24362 14376
rect 24950 17040 25006 17096
rect 25870 18264 25926 18320
rect 25778 17720 25834 17776
rect 27650 20154 27706 20156
rect 27730 20154 27786 20156
rect 27810 20154 27866 20156
rect 27890 20154 27946 20156
rect 27650 20102 27696 20154
rect 27696 20102 27706 20154
rect 27730 20102 27760 20154
rect 27760 20102 27772 20154
rect 27772 20102 27786 20154
rect 27810 20102 27824 20154
rect 27824 20102 27836 20154
rect 27836 20102 27866 20154
rect 27890 20102 27900 20154
rect 27900 20102 27946 20154
rect 27650 20100 27706 20102
rect 27730 20100 27786 20102
rect 27810 20100 27866 20102
rect 27890 20100 27946 20102
rect 26990 19610 27046 19612
rect 27070 19610 27126 19612
rect 27150 19610 27206 19612
rect 27230 19610 27286 19612
rect 26990 19558 27036 19610
rect 27036 19558 27046 19610
rect 27070 19558 27100 19610
rect 27100 19558 27112 19610
rect 27112 19558 27126 19610
rect 27150 19558 27164 19610
rect 27164 19558 27176 19610
rect 27176 19558 27206 19610
rect 27230 19558 27240 19610
rect 27240 19558 27286 19610
rect 26990 19556 27046 19558
rect 27070 19556 27126 19558
rect 27150 19556 27206 19558
rect 27230 19556 27286 19558
rect 26054 17448 26110 17504
rect 25410 15816 25466 15872
rect 24950 13776 25006 13832
rect 25318 14864 25374 14920
rect 25226 14068 25282 14104
rect 25226 14048 25228 14068
rect 25228 14048 25280 14068
rect 25280 14048 25282 14068
rect 22282 12144 22338 12200
rect 22558 12316 22560 12336
rect 22560 12316 22612 12336
rect 22612 12316 22614 12336
rect 22558 12280 22614 12316
rect 22834 12180 22836 12200
rect 22836 12180 22888 12200
rect 22888 12180 22890 12200
rect 22834 12144 22890 12180
rect 22190 9052 22192 9072
rect 22192 9052 22244 9072
rect 22244 9052 22246 9072
rect 22190 9016 22246 9052
rect 22282 8608 22338 8664
rect 22742 10104 22798 10160
rect 23110 12300 23166 12336
rect 23110 12280 23112 12300
rect 23112 12280 23164 12300
rect 23164 12280 23166 12300
rect 22926 8628 22982 8664
rect 22926 8608 22928 8628
rect 22928 8608 22980 8628
rect 22980 8608 22982 8628
rect 23662 9016 23718 9072
rect 24214 9424 24270 9480
rect 25870 15000 25926 15056
rect 26990 18522 27046 18524
rect 27070 18522 27126 18524
rect 27150 18522 27206 18524
rect 27230 18522 27286 18524
rect 26990 18470 27036 18522
rect 27036 18470 27046 18522
rect 27070 18470 27100 18522
rect 27100 18470 27112 18522
rect 27112 18470 27126 18522
rect 27150 18470 27164 18522
rect 27164 18470 27176 18522
rect 27176 18470 27206 18522
rect 27230 18470 27240 18522
rect 27240 18470 27286 18522
rect 26990 18468 27046 18470
rect 27070 18468 27126 18470
rect 27150 18468 27206 18470
rect 27230 18468 27286 18470
rect 27650 19066 27706 19068
rect 27730 19066 27786 19068
rect 27810 19066 27866 19068
rect 27890 19066 27946 19068
rect 27650 19014 27696 19066
rect 27696 19014 27706 19066
rect 27730 19014 27760 19066
rect 27760 19014 27772 19066
rect 27772 19014 27786 19066
rect 27810 19014 27824 19066
rect 27824 19014 27836 19066
rect 27836 19014 27866 19066
rect 27890 19014 27900 19066
rect 27900 19014 27946 19066
rect 27650 19012 27706 19014
rect 27730 19012 27786 19014
rect 27810 19012 27866 19014
rect 27890 19012 27946 19014
rect 28446 19352 28502 19408
rect 29734 19916 29790 19952
rect 29734 19896 29736 19916
rect 29736 19896 29788 19916
rect 29788 19896 29790 19916
rect 30010 19352 30066 19408
rect 27986 18264 28042 18320
rect 27650 17978 27706 17980
rect 27730 17978 27786 17980
rect 27810 17978 27866 17980
rect 27890 17978 27946 17980
rect 27650 17926 27696 17978
rect 27696 17926 27706 17978
rect 27730 17926 27760 17978
rect 27760 17926 27772 17978
rect 27772 17926 27786 17978
rect 27810 17926 27824 17978
rect 27824 17926 27836 17978
rect 27836 17926 27866 17978
rect 27890 17926 27900 17978
rect 27900 17926 27946 17978
rect 27650 17924 27706 17926
rect 27730 17924 27786 17926
rect 27810 17924 27866 17926
rect 27890 17924 27946 17926
rect 26882 17584 26938 17640
rect 26422 14184 26478 14240
rect 26238 12416 26294 12472
rect 22282 6432 22338 6488
rect 22006 6196 22008 6216
rect 22008 6196 22060 6216
rect 22060 6196 22062 6216
rect 22006 6160 22062 6196
rect 21730 5888 21786 5944
rect 22742 5208 22798 5264
rect 22650 4936 22706 4992
rect 19876 2746 19932 2748
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 19876 2694 19922 2746
rect 19922 2694 19932 2746
rect 19956 2694 19986 2746
rect 19986 2694 19998 2746
rect 19998 2694 20012 2746
rect 20036 2694 20050 2746
rect 20050 2694 20062 2746
rect 20062 2694 20092 2746
rect 20116 2694 20126 2746
rect 20126 2694 20172 2746
rect 19876 2692 19932 2694
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 19216 2202 19272 2204
rect 19296 2202 19352 2204
rect 19376 2202 19432 2204
rect 19456 2202 19512 2204
rect 19216 2150 19262 2202
rect 19262 2150 19272 2202
rect 19296 2150 19326 2202
rect 19326 2150 19338 2202
rect 19338 2150 19352 2202
rect 19376 2150 19390 2202
rect 19390 2150 19402 2202
rect 19402 2150 19432 2202
rect 19456 2150 19466 2202
rect 19466 2150 19512 2202
rect 19216 2148 19272 2150
rect 19296 2148 19352 2150
rect 19376 2148 19432 2150
rect 19456 2148 19512 2150
rect 23110 6432 23166 6488
rect 23294 5888 23350 5944
rect 23202 5092 23258 5128
rect 23202 5072 23204 5092
rect 23204 5072 23256 5092
rect 23256 5072 23258 5092
rect 23662 5344 23718 5400
rect 23938 4936 23994 4992
rect 26990 17434 27046 17436
rect 27070 17434 27126 17436
rect 27150 17434 27206 17436
rect 27230 17434 27286 17436
rect 26990 17382 27036 17434
rect 27036 17382 27046 17434
rect 27070 17382 27100 17434
rect 27100 17382 27112 17434
rect 27112 17382 27126 17434
rect 27150 17382 27164 17434
rect 27164 17382 27176 17434
rect 27176 17382 27206 17434
rect 27230 17382 27240 17434
rect 27240 17382 27286 17434
rect 26990 17380 27046 17382
rect 27070 17380 27126 17382
rect 27150 17380 27206 17382
rect 27230 17380 27286 17382
rect 27434 17312 27490 17368
rect 26990 16346 27046 16348
rect 27070 16346 27126 16348
rect 27150 16346 27206 16348
rect 27230 16346 27286 16348
rect 26990 16294 27036 16346
rect 27036 16294 27046 16346
rect 27070 16294 27100 16346
rect 27100 16294 27112 16346
rect 27112 16294 27126 16346
rect 27150 16294 27164 16346
rect 27164 16294 27176 16346
rect 27176 16294 27206 16346
rect 27230 16294 27240 16346
rect 27240 16294 27286 16346
rect 26990 16292 27046 16294
rect 27070 16292 27126 16294
rect 27150 16292 27206 16294
rect 27230 16292 27286 16294
rect 26990 15258 27046 15260
rect 27070 15258 27126 15260
rect 27150 15258 27206 15260
rect 27230 15258 27286 15260
rect 26990 15206 27036 15258
rect 27036 15206 27046 15258
rect 27070 15206 27100 15258
rect 27100 15206 27112 15258
rect 27112 15206 27126 15258
rect 27150 15206 27164 15258
rect 27164 15206 27176 15258
rect 27176 15206 27206 15258
rect 27230 15206 27240 15258
rect 27240 15206 27286 15258
rect 26990 15204 27046 15206
rect 27070 15204 27126 15206
rect 27150 15204 27206 15206
rect 27230 15204 27286 15206
rect 26990 14170 27046 14172
rect 27070 14170 27126 14172
rect 27150 14170 27206 14172
rect 27230 14170 27286 14172
rect 26990 14118 27036 14170
rect 27036 14118 27046 14170
rect 27070 14118 27100 14170
rect 27100 14118 27112 14170
rect 27112 14118 27126 14170
rect 27150 14118 27164 14170
rect 27164 14118 27176 14170
rect 27176 14118 27206 14170
rect 27230 14118 27240 14170
rect 27240 14118 27286 14170
rect 26990 14116 27046 14118
rect 27070 14116 27126 14118
rect 27150 14116 27206 14118
rect 27230 14116 27286 14118
rect 27986 17196 28042 17232
rect 27986 17176 27988 17196
rect 27988 17176 28040 17196
rect 28040 17176 28042 17196
rect 27894 17076 27896 17096
rect 27896 17076 27948 17096
rect 27948 17076 27950 17096
rect 27894 17040 27950 17076
rect 27650 16890 27706 16892
rect 27730 16890 27786 16892
rect 27810 16890 27866 16892
rect 27890 16890 27946 16892
rect 27650 16838 27696 16890
rect 27696 16838 27706 16890
rect 27730 16838 27760 16890
rect 27760 16838 27772 16890
rect 27772 16838 27786 16890
rect 27810 16838 27824 16890
rect 27824 16838 27836 16890
rect 27836 16838 27866 16890
rect 27890 16838 27900 16890
rect 27900 16838 27946 16890
rect 27650 16836 27706 16838
rect 27730 16836 27786 16838
rect 27810 16836 27866 16838
rect 27890 16836 27946 16838
rect 27802 15988 27804 16008
rect 27804 15988 27856 16008
rect 27856 15988 27858 16008
rect 27802 15952 27858 15988
rect 27650 15802 27706 15804
rect 27730 15802 27786 15804
rect 27810 15802 27866 15804
rect 27890 15802 27946 15804
rect 27650 15750 27696 15802
rect 27696 15750 27706 15802
rect 27730 15750 27760 15802
rect 27760 15750 27772 15802
rect 27772 15750 27786 15802
rect 27810 15750 27824 15802
rect 27824 15750 27836 15802
rect 27836 15750 27866 15802
rect 27890 15750 27900 15802
rect 27900 15750 27946 15802
rect 27650 15748 27706 15750
rect 27730 15748 27786 15750
rect 27810 15748 27866 15750
rect 27890 15748 27946 15750
rect 27650 14714 27706 14716
rect 27730 14714 27786 14716
rect 27810 14714 27866 14716
rect 27890 14714 27946 14716
rect 27650 14662 27696 14714
rect 27696 14662 27706 14714
rect 27730 14662 27760 14714
rect 27760 14662 27772 14714
rect 27772 14662 27786 14714
rect 27810 14662 27824 14714
rect 27824 14662 27836 14714
rect 27836 14662 27866 14714
rect 27890 14662 27900 14714
rect 27900 14662 27946 14714
rect 27650 14660 27706 14662
rect 27730 14660 27786 14662
rect 27810 14660 27866 14662
rect 27890 14660 27946 14662
rect 26974 13812 26976 13832
rect 26976 13812 27028 13832
rect 27028 13812 27030 13832
rect 26974 13776 27030 13812
rect 27342 13912 27398 13968
rect 26990 13082 27046 13084
rect 27070 13082 27126 13084
rect 27150 13082 27206 13084
rect 27230 13082 27286 13084
rect 26990 13030 27036 13082
rect 27036 13030 27046 13082
rect 27070 13030 27100 13082
rect 27100 13030 27112 13082
rect 27112 13030 27126 13082
rect 27150 13030 27164 13082
rect 27164 13030 27176 13082
rect 27176 13030 27206 13082
rect 27230 13030 27240 13082
rect 27240 13030 27286 13082
rect 26990 13028 27046 13030
rect 27070 13028 27126 13030
rect 27150 13028 27206 13030
rect 27230 13028 27286 13030
rect 26514 12144 26570 12200
rect 26054 11056 26110 11112
rect 27650 13626 27706 13628
rect 27730 13626 27786 13628
rect 27810 13626 27866 13628
rect 27890 13626 27946 13628
rect 27650 13574 27696 13626
rect 27696 13574 27706 13626
rect 27730 13574 27760 13626
rect 27760 13574 27772 13626
rect 27772 13574 27786 13626
rect 27810 13574 27824 13626
rect 27824 13574 27836 13626
rect 27836 13574 27866 13626
rect 27890 13574 27900 13626
rect 27900 13574 27946 13626
rect 27650 13572 27706 13574
rect 27730 13572 27786 13574
rect 27810 13572 27866 13574
rect 27890 13572 27946 13574
rect 28630 17740 28686 17776
rect 28906 18264 28962 18320
rect 28630 17720 28632 17740
rect 28632 17720 28684 17740
rect 28684 17720 28686 17740
rect 28538 17312 28594 17368
rect 28630 17176 28686 17232
rect 29458 17720 29514 17776
rect 28814 14592 28870 14648
rect 28814 14320 28870 14376
rect 28170 13776 28226 13832
rect 27650 12538 27706 12540
rect 27730 12538 27786 12540
rect 27810 12538 27866 12540
rect 27890 12538 27946 12540
rect 27650 12486 27696 12538
rect 27696 12486 27706 12538
rect 27730 12486 27760 12538
rect 27760 12486 27772 12538
rect 27772 12486 27786 12538
rect 27810 12486 27824 12538
rect 27824 12486 27836 12538
rect 27836 12486 27866 12538
rect 27890 12486 27900 12538
rect 27900 12486 27946 12538
rect 27650 12484 27706 12486
rect 27730 12484 27786 12486
rect 27810 12484 27866 12486
rect 27890 12484 27946 12486
rect 26990 11994 27046 11996
rect 27070 11994 27126 11996
rect 27150 11994 27206 11996
rect 27230 11994 27286 11996
rect 26990 11942 27036 11994
rect 27036 11942 27046 11994
rect 27070 11942 27100 11994
rect 27100 11942 27112 11994
rect 27112 11942 27126 11994
rect 27150 11942 27164 11994
rect 27164 11942 27176 11994
rect 27176 11942 27206 11994
rect 27230 11942 27240 11994
rect 27240 11942 27286 11994
rect 26990 11940 27046 11942
rect 27070 11940 27126 11942
rect 27150 11940 27206 11942
rect 27230 11940 27286 11942
rect 26990 10906 27046 10908
rect 27070 10906 27126 10908
rect 27150 10906 27206 10908
rect 27230 10906 27286 10908
rect 26990 10854 27036 10906
rect 27036 10854 27046 10906
rect 27070 10854 27100 10906
rect 27100 10854 27112 10906
rect 27112 10854 27126 10906
rect 27150 10854 27164 10906
rect 27164 10854 27176 10906
rect 27176 10854 27206 10906
rect 27230 10854 27240 10906
rect 27240 10854 27286 10906
rect 26990 10852 27046 10854
rect 27070 10852 27126 10854
rect 27150 10852 27206 10854
rect 27230 10852 27286 10854
rect 25870 10104 25926 10160
rect 24582 5480 24638 5536
rect 24582 5072 24638 5128
rect 25502 6296 25558 6352
rect 25042 5616 25098 5672
rect 25410 5772 25466 5808
rect 25410 5752 25412 5772
rect 25412 5752 25464 5772
rect 25464 5752 25466 5772
rect 27650 11450 27706 11452
rect 27730 11450 27786 11452
rect 27810 11450 27866 11452
rect 27890 11450 27946 11452
rect 27650 11398 27696 11450
rect 27696 11398 27706 11450
rect 27730 11398 27760 11450
rect 27760 11398 27772 11450
rect 27772 11398 27786 11450
rect 27810 11398 27824 11450
rect 27824 11398 27836 11450
rect 27836 11398 27866 11450
rect 27890 11398 27900 11450
rect 27900 11398 27946 11450
rect 27650 11396 27706 11398
rect 27730 11396 27786 11398
rect 27810 11396 27866 11398
rect 27890 11396 27946 11398
rect 30562 14592 30618 14648
rect 30930 14476 30986 14512
rect 30930 14456 30932 14476
rect 30932 14456 30984 14476
rect 30984 14456 30986 14476
rect 27650 10362 27706 10364
rect 27730 10362 27786 10364
rect 27810 10362 27866 10364
rect 27890 10362 27946 10364
rect 27650 10310 27696 10362
rect 27696 10310 27706 10362
rect 27730 10310 27760 10362
rect 27760 10310 27772 10362
rect 27772 10310 27786 10362
rect 27810 10310 27824 10362
rect 27824 10310 27836 10362
rect 27836 10310 27866 10362
rect 27890 10310 27900 10362
rect 27900 10310 27946 10362
rect 27650 10308 27706 10310
rect 27730 10308 27786 10310
rect 27810 10308 27866 10310
rect 27890 10308 27946 10310
rect 27434 10124 27490 10160
rect 27434 10104 27436 10124
rect 27436 10104 27488 10124
rect 27488 10104 27490 10124
rect 26990 9818 27046 9820
rect 27070 9818 27126 9820
rect 27150 9818 27206 9820
rect 27230 9818 27286 9820
rect 26990 9766 27036 9818
rect 27036 9766 27046 9818
rect 27070 9766 27100 9818
rect 27100 9766 27112 9818
rect 27112 9766 27126 9818
rect 27150 9766 27164 9818
rect 27164 9766 27176 9818
rect 27176 9766 27206 9818
rect 27230 9766 27240 9818
rect 27240 9766 27286 9818
rect 26990 9764 27046 9766
rect 27070 9764 27126 9766
rect 27150 9764 27206 9766
rect 27230 9764 27286 9766
rect 26990 8730 27046 8732
rect 27070 8730 27126 8732
rect 27150 8730 27206 8732
rect 27230 8730 27286 8732
rect 26990 8678 27036 8730
rect 27036 8678 27046 8730
rect 27070 8678 27100 8730
rect 27100 8678 27112 8730
rect 27112 8678 27126 8730
rect 27150 8678 27164 8730
rect 27164 8678 27176 8730
rect 27176 8678 27206 8730
rect 27230 8678 27240 8730
rect 27240 8678 27286 8730
rect 26990 8676 27046 8678
rect 27070 8676 27126 8678
rect 27150 8676 27206 8678
rect 27230 8676 27286 8678
rect 27650 9274 27706 9276
rect 27730 9274 27786 9276
rect 27810 9274 27866 9276
rect 27890 9274 27946 9276
rect 27650 9222 27696 9274
rect 27696 9222 27706 9274
rect 27730 9222 27760 9274
rect 27760 9222 27772 9274
rect 27772 9222 27786 9274
rect 27810 9222 27824 9274
rect 27824 9222 27836 9274
rect 27836 9222 27866 9274
rect 27890 9222 27900 9274
rect 27900 9222 27946 9274
rect 27650 9220 27706 9222
rect 27730 9220 27786 9222
rect 27810 9220 27866 9222
rect 27890 9220 27946 9222
rect 27650 8186 27706 8188
rect 27730 8186 27786 8188
rect 27810 8186 27866 8188
rect 27890 8186 27946 8188
rect 27650 8134 27696 8186
rect 27696 8134 27706 8186
rect 27730 8134 27760 8186
rect 27760 8134 27772 8186
rect 27772 8134 27786 8186
rect 27810 8134 27824 8186
rect 27824 8134 27836 8186
rect 27836 8134 27866 8186
rect 27890 8134 27900 8186
rect 27900 8134 27946 8186
rect 27650 8132 27706 8134
rect 27730 8132 27786 8134
rect 27810 8132 27866 8134
rect 27890 8132 27946 8134
rect 26990 7642 27046 7644
rect 27070 7642 27126 7644
rect 27150 7642 27206 7644
rect 27230 7642 27286 7644
rect 26990 7590 27036 7642
rect 27036 7590 27046 7642
rect 27070 7590 27100 7642
rect 27100 7590 27112 7642
rect 27112 7590 27126 7642
rect 27150 7590 27164 7642
rect 27164 7590 27176 7642
rect 27176 7590 27206 7642
rect 27230 7590 27240 7642
rect 27240 7590 27286 7642
rect 26990 7588 27046 7590
rect 27070 7588 27126 7590
rect 27150 7588 27206 7590
rect 27230 7588 27286 7590
rect 27650 7098 27706 7100
rect 27730 7098 27786 7100
rect 27810 7098 27866 7100
rect 27890 7098 27946 7100
rect 27650 7046 27696 7098
rect 27696 7046 27706 7098
rect 27730 7046 27760 7098
rect 27760 7046 27772 7098
rect 27772 7046 27786 7098
rect 27810 7046 27824 7098
rect 27824 7046 27836 7098
rect 27836 7046 27866 7098
rect 27890 7046 27900 7098
rect 27900 7046 27946 7098
rect 27650 7044 27706 7046
rect 27730 7044 27786 7046
rect 27810 7044 27866 7046
rect 27890 7044 27946 7046
rect 26990 6554 27046 6556
rect 27070 6554 27126 6556
rect 27150 6554 27206 6556
rect 27230 6554 27286 6556
rect 26990 6502 27036 6554
rect 27036 6502 27046 6554
rect 27070 6502 27100 6554
rect 27100 6502 27112 6554
rect 27112 6502 27126 6554
rect 27150 6502 27164 6554
rect 27164 6502 27176 6554
rect 27176 6502 27206 6554
rect 27230 6502 27240 6554
rect 27240 6502 27286 6554
rect 26990 6500 27046 6502
rect 27070 6500 27126 6502
rect 27150 6500 27206 6502
rect 27230 6500 27286 6502
rect 26698 6160 26754 6216
rect 27650 6010 27706 6012
rect 27730 6010 27786 6012
rect 27810 6010 27866 6012
rect 27890 6010 27946 6012
rect 27650 5958 27696 6010
rect 27696 5958 27706 6010
rect 27730 5958 27760 6010
rect 27760 5958 27772 6010
rect 27772 5958 27786 6010
rect 27810 5958 27824 6010
rect 27824 5958 27836 6010
rect 27836 5958 27866 6010
rect 27890 5958 27900 6010
rect 27900 5958 27946 6010
rect 27650 5956 27706 5958
rect 27730 5956 27786 5958
rect 27810 5956 27866 5958
rect 27890 5956 27946 5958
rect 26990 5466 27046 5468
rect 27070 5466 27126 5468
rect 27150 5466 27206 5468
rect 27230 5466 27286 5468
rect 26990 5414 27036 5466
rect 27036 5414 27046 5466
rect 27070 5414 27100 5466
rect 27100 5414 27112 5466
rect 27112 5414 27126 5466
rect 27150 5414 27164 5466
rect 27164 5414 27176 5466
rect 27176 5414 27206 5466
rect 27230 5414 27240 5466
rect 27240 5414 27286 5466
rect 26990 5412 27046 5414
rect 27070 5412 27126 5414
rect 27150 5412 27206 5414
rect 27230 5412 27286 5414
rect 21638 2508 21694 2544
rect 21638 2488 21640 2508
rect 21640 2488 21692 2508
rect 21692 2488 21694 2508
rect 22650 2508 22706 2544
rect 22650 2488 22652 2508
rect 22652 2488 22704 2508
rect 22704 2488 22706 2508
rect 19876 1658 19932 1660
rect 19956 1658 20012 1660
rect 20036 1658 20092 1660
rect 20116 1658 20172 1660
rect 19876 1606 19922 1658
rect 19922 1606 19932 1658
rect 19956 1606 19986 1658
rect 19986 1606 19998 1658
rect 19998 1606 20012 1658
rect 20036 1606 20050 1658
rect 20050 1606 20062 1658
rect 20062 1606 20092 1658
rect 20116 1606 20126 1658
rect 20126 1606 20172 1658
rect 19876 1604 19932 1606
rect 19956 1604 20012 1606
rect 20036 1604 20092 1606
rect 20116 1604 20172 1606
rect 27650 4922 27706 4924
rect 27730 4922 27786 4924
rect 27810 4922 27866 4924
rect 27890 4922 27946 4924
rect 27650 4870 27696 4922
rect 27696 4870 27706 4922
rect 27730 4870 27760 4922
rect 27760 4870 27772 4922
rect 27772 4870 27786 4922
rect 27810 4870 27824 4922
rect 27824 4870 27836 4922
rect 27836 4870 27866 4922
rect 27890 4870 27900 4922
rect 27900 4870 27946 4922
rect 27650 4868 27706 4870
rect 27730 4868 27786 4870
rect 27810 4868 27866 4870
rect 27890 4868 27946 4870
rect 26990 4378 27046 4380
rect 27070 4378 27126 4380
rect 27150 4378 27206 4380
rect 27230 4378 27286 4380
rect 26990 4326 27036 4378
rect 27036 4326 27046 4378
rect 27070 4326 27100 4378
rect 27100 4326 27112 4378
rect 27112 4326 27126 4378
rect 27150 4326 27164 4378
rect 27164 4326 27176 4378
rect 27176 4326 27206 4378
rect 27230 4326 27240 4378
rect 27240 4326 27286 4378
rect 26990 4324 27046 4326
rect 27070 4324 27126 4326
rect 27150 4324 27206 4326
rect 27230 4324 27286 4326
rect 30194 6724 30250 6760
rect 30194 6704 30196 6724
rect 30196 6704 30248 6724
rect 30248 6704 30250 6724
rect 27650 3834 27706 3836
rect 27730 3834 27786 3836
rect 27810 3834 27866 3836
rect 27890 3834 27946 3836
rect 27650 3782 27696 3834
rect 27696 3782 27706 3834
rect 27730 3782 27760 3834
rect 27760 3782 27772 3834
rect 27772 3782 27786 3834
rect 27810 3782 27824 3834
rect 27824 3782 27836 3834
rect 27836 3782 27866 3834
rect 27890 3782 27900 3834
rect 27900 3782 27946 3834
rect 27650 3780 27706 3782
rect 27730 3780 27786 3782
rect 27810 3780 27866 3782
rect 27890 3780 27946 3782
rect 26990 3290 27046 3292
rect 27070 3290 27126 3292
rect 27150 3290 27206 3292
rect 27230 3290 27286 3292
rect 26990 3238 27036 3290
rect 27036 3238 27046 3290
rect 27070 3238 27100 3290
rect 27100 3238 27112 3290
rect 27112 3238 27126 3290
rect 27150 3238 27164 3290
rect 27164 3238 27176 3290
rect 27176 3238 27206 3290
rect 27230 3238 27240 3290
rect 27240 3238 27286 3290
rect 26990 3236 27046 3238
rect 27070 3236 27126 3238
rect 27150 3236 27206 3238
rect 27230 3236 27286 3238
rect 27650 2746 27706 2748
rect 27730 2746 27786 2748
rect 27810 2746 27866 2748
rect 27890 2746 27946 2748
rect 27650 2694 27696 2746
rect 27696 2694 27706 2746
rect 27730 2694 27760 2746
rect 27760 2694 27772 2746
rect 27772 2694 27786 2746
rect 27810 2694 27824 2746
rect 27824 2694 27836 2746
rect 27836 2694 27866 2746
rect 27890 2694 27900 2746
rect 27900 2694 27946 2746
rect 27650 2692 27706 2694
rect 27730 2692 27786 2694
rect 27810 2692 27866 2694
rect 27890 2692 27946 2694
rect 26990 2202 27046 2204
rect 27070 2202 27126 2204
rect 27150 2202 27206 2204
rect 27230 2202 27286 2204
rect 26990 2150 27036 2202
rect 27036 2150 27046 2202
rect 27070 2150 27100 2202
rect 27100 2150 27112 2202
rect 27112 2150 27126 2202
rect 27150 2150 27164 2202
rect 27164 2150 27176 2202
rect 27176 2150 27206 2202
rect 27230 2150 27240 2202
rect 27240 2150 27286 2202
rect 26990 2148 27046 2150
rect 27070 2148 27126 2150
rect 27150 2148 27206 2150
rect 27230 2148 27286 2150
rect 27650 1658 27706 1660
rect 27730 1658 27786 1660
rect 27810 1658 27866 1660
rect 27890 1658 27946 1660
rect 27650 1606 27696 1658
rect 27696 1606 27706 1658
rect 27730 1606 27760 1658
rect 27760 1606 27772 1658
rect 27772 1606 27786 1658
rect 27810 1606 27824 1658
rect 27824 1606 27836 1658
rect 27836 1606 27866 1658
rect 27890 1606 27900 1658
rect 27900 1606 27946 1658
rect 27650 1604 27706 1606
rect 27730 1604 27786 1606
rect 27810 1604 27866 1606
rect 27890 1604 27946 1606
rect 19216 1114 19272 1116
rect 19296 1114 19352 1116
rect 19376 1114 19432 1116
rect 19456 1114 19512 1116
rect 19216 1062 19262 1114
rect 19262 1062 19272 1114
rect 19296 1062 19326 1114
rect 19326 1062 19338 1114
rect 19338 1062 19352 1114
rect 19376 1062 19390 1114
rect 19390 1062 19402 1114
rect 19402 1062 19432 1114
rect 19456 1062 19466 1114
rect 19466 1062 19512 1114
rect 19216 1060 19272 1062
rect 19296 1060 19352 1062
rect 19376 1060 19432 1062
rect 19456 1060 19512 1062
rect 26990 1114 27046 1116
rect 27070 1114 27126 1116
rect 27150 1114 27206 1116
rect 27230 1114 27286 1116
rect 26990 1062 27036 1114
rect 27036 1062 27046 1114
rect 27070 1062 27100 1114
rect 27100 1062 27112 1114
rect 27112 1062 27126 1114
rect 27150 1062 27164 1114
rect 27164 1062 27176 1114
rect 27176 1062 27206 1114
rect 27230 1062 27240 1114
rect 27240 1062 27286 1114
rect 26990 1060 27046 1062
rect 27070 1060 27126 1062
rect 27150 1060 27206 1062
rect 27230 1060 27286 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 12102 570 12158 572
rect 12182 570 12238 572
rect 12262 570 12318 572
rect 12342 570 12398 572
rect 12102 518 12148 570
rect 12148 518 12158 570
rect 12182 518 12212 570
rect 12212 518 12224 570
rect 12224 518 12238 570
rect 12262 518 12276 570
rect 12276 518 12288 570
rect 12288 518 12318 570
rect 12342 518 12352 570
rect 12352 518 12398 570
rect 12102 516 12158 518
rect 12182 516 12238 518
rect 12262 516 12318 518
rect 12342 516 12398 518
rect 19876 570 19932 572
rect 19956 570 20012 572
rect 20036 570 20092 572
rect 20116 570 20172 572
rect 19876 518 19922 570
rect 19922 518 19932 570
rect 19956 518 19986 570
rect 19986 518 19998 570
rect 19998 518 20012 570
rect 20036 518 20050 570
rect 20050 518 20062 570
rect 20062 518 20092 570
rect 20116 518 20126 570
rect 20126 518 20172 570
rect 19876 516 19932 518
rect 19956 516 20012 518
rect 20036 516 20092 518
rect 20116 516 20172 518
rect 27650 570 27706 572
rect 27730 570 27786 572
rect 27810 570 27866 572
rect 27890 570 27946 572
rect 27650 518 27696 570
rect 27696 518 27706 570
rect 27730 518 27760 570
rect 27760 518 27772 570
rect 27772 518 27786 570
rect 27810 518 27824 570
rect 27824 518 27836 570
rect 27836 518 27866 570
rect 27890 518 27900 570
rect 27900 518 27946 570
rect 27650 516 27706 518
rect 27730 516 27786 518
rect 27810 516 27866 518
rect 27890 516 27946 518
<< metal3 >>
rect 11646 21932 11652 21996
rect 11716 21994 11722 21996
rect 11789 21994 11855 21997
rect 12249 21996 12315 21997
rect 24393 21996 24459 21997
rect 11716 21992 11855 21994
rect 11716 21936 11794 21992
rect 11850 21936 11855 21992
rect 11716 21934 11855 21936
rect 11716 21932 11722 21934
rect 11789 21931 11855 21934
rect 12198 21932 12204 21996
rect 12268 21994 12315 21996
rect 24342 21994 24348 21996
rect 12268 21992 12360 21994
rect 12310 21936 12360 21992
rect 12268 21934 12360 21936
rect 24302 21934 24348 21994
rect 24412 21992 24459 21996
rect 24454 21936 24459 21992
rect 12268 21932 12315 21934
rect 24342 21932 24348 21934
rect 24412 21932 24459 21936
rect 27102 21932 27108 21996
rect 27172 21994 27178 21996
rect 27337 21994 27403 21997
rect 27705 21996 27771 21997
rect 27654 21994 27660 21996
rect 27172 21992 27403 21994
rect 27172 21936 27342 21992
rect 27398 21936 27403 21992
rect 27172 21934 27403 21936
rect 27614 21934 27660 21994
rect 27724 21992 27771 21996
rect 27766 21936 27771 21992
rect 27172 21932 27178 21934
rect 12249 21931 12315 21932
rect 24393 21931 24459 21932
rect 27337 21931 27403 21934
rect 27654 21932 27660 21934
rect 27724 21932 27771 21936
rect 27705 21931 27771 21932
rect 7230 21796 7236 21860
rect 7300 21858 7306 21860
rect 8661 21858 8727 21861
rect 7300 21856 8727 21858
rect 7300 21800 8666 21856
rect 8722 21800 8727 21856
rect 7300 21798 8727 21800
rect 7300 21796 7306 21798
rect 8661 21795 8727 21798
rect 21582 21796 21588 21860
rect 21652 21858 21658 21860
rect 22185 21858 22251 21861
rect 23841 21860 23907 21861
rect 23790 21858 23796 21860
rect 21652 21856 22251 21858
rect 21652 21800 22190 21856
rect 22246 21800 22251 21856
rect 21652 21798 22251 21800
rect 23750 21798 23796 21858
rect 23860 21856 23907 21860
rect 23902 21800 23907 21856
rect 21652 21796 21658 21798
rect 22185 21795 22251 21798
rect 23790 21796 23796 21798
rect 23860 21796 23907 21800
rect 25998 21796 26004 21860
rect 26068 21858 26074 21860
rect 26417 21858 26483 21861
rect 26068 21856 26483 21858
rect 26068 21800 26422 21856
rect 26478 21800 26483 21856
rect 26068 21798 26483 21800
rect 26068 21796 26074 21798
rect 23841 21795 23907 21796
rect 26417 21795 26483 21798
rect 26550 21796 26556 21860
rect 26620 21858 26626 21860
rect 26693 21858 26759 21861
rect 28257 21860 28323 21861
rect 28206 21858 28212 21860
rect 26620 21856 26759 21858
rect 26620 21800 26698 21856
rect 26754 21800 26759 21856
rect 26620 21798 26759 21800
rect 28166 21798 28212 21858
rect 28276 21856 28323 21860
rect 28318 21800 28323 21856
rect 26620 21796 26626 21798
rect 26693 21795 26759 21798
rect 28206 21796 28212 21798
rect 28276 21796 28323 21800
rect 28257 21795 28323 21796
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 11432 21792 11748 21793
rect 11432 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11748 21792
rect 11432 21727 11748 21728
rect 19206 21792 19522 21793
rect 19206 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19522 21792
rect 19206 21727 19522 21728
rect 26980 21792 27296 21793
rect 26980 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27296 21792
rect 26980 21727 27296 21728
rect 6085 21724 6151 21725
rect 6085 21722 6132 21724
rect 6040 21720 6132 21722
rect 6040 21664 6090 21720
rect 6040 21662 6132 21664
rect 6085 21660 6132 21662
rect 6196 21660 6202 21724
rect 7782 21660 7788 21724
rect 7852 21722 7858 21724
rect 8017 21722 8083 21725
rect 8385 21724 8451 21725
rect 7852 21720 8083 21722
rect 7852 21664 8022 21720
rect 8078 21664 8083 21720
rect 7852 21662 8083 21664
rect 7852 21660 7858 21662
rect 6085 21659 6151 21660
rect 8017 21659 8083 21662
rect 8334 21660 8340 21724
rect 8404 21722 8451 21724
rect 8404 21720 8496 21722
rect 8446 21664 8496 21720
rect 8404 21662 8496 21664
rect 8404 21660 8451 21662
rect 12750 21660 12756 21724
rect 12820 21722 12826 21724
rect 12985 21722 13051 21725
rect 12820 21720 13051 21722
rect 12820 21664 12990 21720
rect 13046 21664 13051 21720
rect 12820 21662 13051 21664
rect 12820 21660 12826 21662
rect 8385 21659 8451 21660
rect 12985 21659 13051 21662
rect 24894 21660 24900 21724
rect 24964 21722 24970 21724
rect 25313 21722 25379 21725
rect 24964 21720 25379 21722
rect 24964 21664 25318 21720
rect 25374 21664 25379 21720
rect 24964 21662 25379 21664
rect 24964 21660 24970 21662
rect 25313 21659 25379 21662
rect 25497 21588 25563 21589
rect 25446 21586 25452 21588
rect 25406 21526 25452 21586
rect 25516 21584 25563 21588
rect 25558 21528 25563 21584
rect 25446 21524 25452 21526
rect 25516 21524 25563 21528
rect 25497 21523 25563 21524
rect 17166 21388 17172 21452
rect 17236 21450 17242 21452
rect 18045 21450 18111 21453
rect 17236 21448 18111 21450
rect 17236 21392 18050 21448
rect 18106 21392 18111 21448
rect 17236 21390 18111 21392
rect 17236 21388 17242 21390
rect 18045 21387 18111 21390
rect 8937 21314 9003 21317
rect 9438 21314 9444 21316
rect 8937 21312 9444 21314
rect 8937 21256 8942 21312
rect 8998 21256 9444 21312
rect 8937 21254 9444 21256
rect 8937 21251 9003 21254
rect 9438 21252 9444 21254
rect 9508 21252 9514 21316
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 12092 21248 12408 21249
rect 12092 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12408 21248
rect 12092 21183 12408 21184
rect 19866 21248 20182 21249
rect 19866 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20182 21248
rect 19866 21183 20182 21184
rect 27640 21248 27956 21249
rect 27640 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27956 21248
rect 27640 21183 27956 21184
rect 8569 21178 8635 21181
rect 8886 21178 8892 21180
rect 8569 21176 8892 21178
rect 8569 21120 8574 21176
rect 8630 21120 8892 21176
rect 8569 21118 8892 21120
rect 8569 21115 8635 21118
rect 8886 21116 8892 21118
rect 8956 21116 8962 21180
rect 9765 21178 9831 21181
rect 9990 21178 9996 21180
rect 9765 21176 9996 21178
rect 9765 21120 9770 21176
rect 9826 21120 9996 21176
rect 9765 21118 9996 21120
rect 9765 21115 9831 21118
rect 9990 21116 9996 21118
rect 10060 21116 10066 21180
rect 18270 21116 18276 21180
rect 18340 21178 18346 21180
rect 19701 21178 19767 21181
rect 18340 21176 19767 21178
rect 18340 21120 19706 21176
rect 19762 21120 19767 21176
rect 18340 21118 19767 21120
rect 18340 21116 18346 21118
rect 19701 21115 19767 21118
rect 18822 20980 18828 21044
rect 18892 21042 18898 21044
rect 19517 21042 19583 21045
rect 18892 21040 19583 21042
rect 18892 20984 19522 21040
rect 19578 20984 19583 21040
rect 18892 20982 19583 20984
rect 18892 20980 18898 20982
rect 19517 20979 19583 20982
rect 15193 20906 15259 20909
rect 16062 20906 16068 20908
rect 15193 20904 16068 20906
rect 15193 20848 15198 20904
rect 15254 20848 16068 20904
rect 15193 20846 16068 20848
rect 15193 20843 15259 20846
rect 16062 20844 16068 20846
rect 16132 20844 16138 20908
rect 15510 20708 15516 20772
rect 15580 20770 15586 20772
rect 16205 20770 16271 20773
rect 15580 20768 16271 20770
rect 15580 20712 16210 20768
rect 16266 20712 16271 20768
rect 15580 20710 16271 20712
rect 15580 20708 15586 20710
rect 16205 20707 16271 20710
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 11432 20704 11748 20705
rect 11432 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11748 20704
rect 11432 20639 11748 20640
rect 19206 20704 19522 20705
rect 19206 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19522 20704
rect 19206 20639 19522 20640
rect 26980 20704 27296 20705
rect 26980 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27296 20704
rect 26980 20639 27296 20640
rect 11053 20636 11119 20637
rect 13261 20636 13327 20637
rect 11053 20634 11100 20636
rect 11008 20632 11100 20634
rect 11008 20576 11058 20632
rect 11008 20574 11100 20576
rect 11053 20572 11100 20574
rect 11164 20572 11170 20636
rect 13261 20632 13308 20636
rect 13372 20634 13378 20636
rect 13261 20576 13266 20632
rect 13261 20572 13308 20576
rect 13372 20574 13418 20634
rect 13372 20572 13378 20574
rect 14958 20572 14964 20636
rect 15028 20634 15034 20636
rect 15469 20634 15535 20637
rect 15028 20632 15535 20634
rect 15028 20576 15474 20632
rect 15530 20576 15535 20632
rect 15028 20574 15535 20576
rect 15028 20572 15034 20574
rect 11053 20571 11119 20572
rect 13261 20571 13327 20572
rect 15469 20571 15535 20574
rect 16481 20634 16547 20637
rect 16614 20634 16620 20636
rect 16481 20632 16620 20634
rect 16481 20576 16486 20632
rect 16542 20576 16620 20632
rect 16481 20574 16620 20576
rect 16481 20571 16547 20574
rect 16614 20572 16620 20574
rect 16684 20572 16690 20636
rect 9949 20498 10015 20501
rect 14273 20498 14339 20501
rect 18965 20498 19031 20501
rect 9949 20496 19031 20498
rect 9949 20440 9954 20496
rect 10010 20440 14278 20496
rect 14334 20440 18970 20496
rect 19026 20440 19031 20496
rect 9949 20438 19031 20440
rect 9949 20435 10015 20438
rect 14273 20435 14339 20438
rect 18965 20435 19031 20438
rect 20897 20498 20963 20501
rect 21541 20498 21607 20501
rect 20897 20496 21607 20498
rect 20897 20440 20902 20496
rect 20958 20440 21546 20496
rect 21602 20440 21607 20496
rect 20897 20438 21607 20440
rect 20897 20435 20963 20438
rect 21541 20435 21607 20438
rect 6729 20364 6795 20365
rect 6678 20300 6684 20364
rect 6748 20362 6795 20364
rect 15837 20362 15903 20365
rect 18781 20362 18847 20365
rect 6748 20360 6840 20362
rect 6790 20304 6840 20360
rect 6748 20302 6840 20304
rect 15837 20360 18847 20362
rect 15837 20304 15842 20360
rect 15898 20304 18786 20360
rect 18842 20304 18847 20360
rect 15837 20302 18847 20304
rect 6748 20300 6795 20302
rect 6729 20299 6795 20300
rect 15837 20299 15903 20302
rect 18781 20299 18847 20302
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 12092 20160 12408 20161
rect 12092 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12408 20160
rect 12092 20095 12408 20096
rect 19866 20160 20182 20161
rect 19866 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20182 20160
rect 19866 20095 20182 20096
rect 27640 20160 27956 20161
rect 27640 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27956 20160
rect 27640 20095 27956 20096
rect 15561 20090 15627 20093
rect 22461 20090 22527 20093
rect 26509 20090 26575 20093
rect 15561 20088 18154 20090
rect 15561 20032 15566 20088
rect 15622 20032 18154 20088
rect 15561 20030 18154 20032
rect 15561 20027 15627 20030
rect 17718 19892 17724 19956
rect 17788 19954 17794 19956
rect 17953 19954 18019 19957
rect 17788 19952 18019 19954
rect 17788 19896 17958 19952
rect 18014 19896 18019 19952
rect 17788 19894 18019 19896
rect 18094 19954 18154 20030
rect 22461 20088 26575 20090
rect 22461 20032 22466 20088
rect 22522 20032 26514 20088
rect 26570 20032 26575 20088
rect 22461 20030 26575 20032
rect 22461 20027 22527 20030
rect 26509 20027 26575 20030
rect 29729 19954 29795 19957
rect 18094 19952 29795 19954
rect 18094 19896 29734 19952
rect 29790 19896 29795 19952
rect 18094 19894 29795 19896
rect 17788 19892 17794 19894
rect 17953 19891 18019 19894
rect 29729 19891 29795 19894
rect 18045 19818 18111 19821
rect 19333 19818 19399 19821
rect 18045 19816 19399 19818
rect 18045 19760 18050 19816
rect 18106 19760 19338 19816
rect 19394 19760 19399 19816
rect 18045 19758 19399 19760
rect 18045 19755 18111 19758
rect 19333 19755 19399 19758
rect 14825 19682 14891 19685
rect 18873 19682 18939 19685
rect 14825 19680 18939 19682
rect 14825 19624 14830 19680
rect 14886 19624 18878 19680
rect 18934 19624 18939 19680
rect 14825 19622 18939 19624
rect 14825 19619 14891 19622
rect 18873 19619 18939 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 3658 19551 3974 19552
rect 11432 19616 11748 19617
rect 11432 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11748 19616
rect 11432 19551 11748 19552
rect 19206 19616 19522 19617
rect 19206 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19522 19616
rect 19206 19551 19522 19552
rect 26980 19616 27296 19617
rect 26980 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27296 19616
rect 26980 19551 27296 19552
rect 8937 19410 9003 19413
rect 10685 19410 10751 19413
rect 8937 19408 10751 19410
rect 8937 19352 8942 19408
rect 8998 19352 10690 19408
rect 10746 19352 10751 19408
rect 8937 19350 10751 19352
rect 8937 19347 9003 19350
rect 10685 19347 10751 19350
rect 25129 19410 25195 19413
rect 28441 19410 28507 19413
rect 30005 19410 30071 19413
rect 25129 19408 30071 19410
rect 25129 19352 25134 19408
rect 25190 19352 28446 19408
rect 28502 19352 30010 19408
rect 30066 19352 30071 19408
rect 25129 19350 30071 19352
rect 25129 19347 25195 19350
rect 28441 19347 28507 19350
rect 30005 19347 30071 19350
rect 8201 19274 8267 19277
rect 14406 19274 14412 19276
rect 8201 19272 14412 19274
rect 8201 19216 8206 19272
rect 8262 19216 14412 19272
rect 8201 19214 14412 19216
rect 8201 19211 8267 19214
rect 14406 19212 14412 19214
rect 14476 19212 14482 19276
rect 15009 19274 15075 19277
rect 17217 19274 17283 19277
rect 15009 19272 17283 19274
rect 15009 19216 15014 19272
rect 15070 19216 17222 19272
rect 17278 19216 17283 19272
rect 15009 19214 17283 19216
rect 15009 19211 15075 19214
rect 17217 19211 17283 19214
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 12092 19072 12408 19073
rect 12092 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12408 19072
rect 12092 19007 12408 19008
rect 19866 19072 20182 19073
rect 19866 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20182 19072
rect 19866 19007 20182 19008
rect 27640 19072 27956 19073
rect 27640 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27956 19072
rect 27640 19007 27956 19008
rect 7833 18866 7899 18869
rect 13854 18866 13860 18868
rect 7833 18864 13860 18866
rect 7833 18808 7838 18864
rect 7894 18808 13860 18864
rect 7833 18806 13860 18808
rect 7833 18803 7899 18806
rect 13854 18804 13860 18806
rect 13924 18804 13930 18868
rect 8661 18730 8727 18733
rect 24025 18730 24091 18733
rect 8661 18728 24091 18730
rect 8661 18672 8666 18728
rect 8722 18672 24030 18728
rect 24086 18672 24091 18728
rect 8661 18670 24091 18672
rect 8661 18667 8727 18670
rect 24025 18667 24091 18670
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 11432 18528 11748 18529
rect 11432 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11748 18528
rect 11432 18463 11748 18464
rect 19206 18528 19522 18529
rect 19206 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19522 18528
rect 19206 18463 19522 18464
rect 26980 18528 27296 18529
rect 26980 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27296 18528
rect 26980 18463 27296 18464
rect 15193 18322 15259 18325
rect 16113 18322 16179 18325
rect 15193 18320 16179 18322
rect 15193 18264 15198 18320
rect 15254 18264 16118 18320
rect 16174 18264 16179 18320
rect 15193 18262 16179 18264
rect 15193 18259 15259 18262
rect 16113 18259 16179 18262
rect 25865 18322 25931 18325
rect 27981 18322 28047 18325
rect 28901 18322 28967 18325
rect 25865 18320 28967 18322
rect 25865 18264 25870 18320
rect 25926 18264 27986 18320
rect 28042 18264 28906 18320
rect 28962 18264 28967 18320
rect 25865 18262 28967 18264
rect 25865 18259 25931 18262
rect 27981 18259 28047 18262
rect 28901 18259 28967 18262
rect 15009 18186 15075 18189
rect 20294 18186 20300 18188
rect 15009 18184 20300 18186
rect 15009 18128 15014 18184
rect 15070 18128 20300 18184
rect 15009 18126 20300 18128
rect 15009 18123 15075 18126
rect 20294 18124 20300 18126
rect 20364 18186 20370 18188
rect 25129 18186 25195 18189
rect 20364 18184 25195 18186
rect 20364 18128 25134 18184
rect 25190 18128 25195 18184
rect 20364 18126 25195 18128
rect 20364 18124 20370 18126
rect 25129 18123 25195 18126
rect 12893 18050 12959 18053
rect 14733 18050 14799 18053
rect 18321 18050 18387 18053
rect 19241 18050 19307 18053
rect 12893 18048 19307 18050
rect 12893 17992 12898 18048
rect 12954 17992 14738 18048
rect 14794 17992 18326 18048
rect 18382 17992 19246 18048
rect 19302 17992 19307 18048
rect 12893 17990 19307 17992
rect 12893 17987 12959 17990
rect 14733 17987 14799 17990
rect 18321 17987 18387 17990
rect 19241 17987 19307 17990
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 12092 17984 12408 17985
rect 12092 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12408 17984
rect 12092 17919 12408 17920
rect 19866 17984 20182 17985
rect 19866 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20182 17984
rect 19866 17919 20182 17920
rect 27640 17984 27956 17985
rect 27640 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27956 17984
rect 27640 17919 27956 17920
rect 10041 17914 10107 17917
rect 10777 17914 10843 17917
rect 10041 17912 10843 17914
rect 10041 17856 10046 17912
rect 10102 17856 10782 17912
rect 10838 17856 10843 17912
rect 10041 17854 10843 17856
rect 10041 17851 10107 17854
rect 10777 17851 10843 17854
rect 21449 17914 21515 17917
rect 25221 17914 25287 17917
rect 21449 17912 25287 17914
rect 21449 17856 21454 17912
rect 21510 17856 25226 17912
rect 25282 17856 25287 17912
rect 21449 17854 25287 17856
rect 21449 17851 21515 17854
rect 25221 17851 25287 17854
rect 10593 17778 10659 17781
rect 16113 17778 16179 17781
rect 10593 17776 16179 17778
rect 10593 17720 10598 17776
rect 10654 17720 16118 17776
rect 16174 17720 16179 17776
rect 10593 17718 16179 17720
rect 10593 17715 10659 17718
rect 16113 17715 16179 17718
rect 25773 17778 25839 17781
rect 28625 17778 28691 17781
rect 29453 17778 29519 17781
rect 25773 17776 29519 17778
rect 25773 17720 25778 17776
rect 25834 17720 28630 17776
rect 28686 17720 29458 17776
rect 29514 17720 29519 17776
rect 25773 17718 29519 17720
rect 25773 17715 25839 17718
rect 28625 17715 28691 17718
rect 29453 17715 29519 17718
rect 4153 17642 4219 17645
rect 4705 17642 4771 17645
rect 4981 17642 5047 17645
rect 4153 17640 5047 17642
rect 4153 17584 4158 17640
rect 4214 17584 4710 17640
rect 4766 17584 4986 17640
rect 5042 17584 5047 17640
rect 4153 17582 5047 17584
rect 4153 17579 4219 17582
rect 4705 17579 4771 17582
rect 4981 17579 5047 17582
rect 11605 17642 11671 17645
rect 18597 17642 18663 17645
rect 11605 17640 18663 17642
rect 11605 17584 11610 17640
rect 11666 17584 18602 17640
rect 18658 17584 18663 17640
rect 11605 17582 18663 17584
rect 11605 17579 11671 17582
rect 18597 17579 18663 17582
rect 24669 17642 24735 17645
rect 26877 17642 26943 17645
rect 24669 17640 26943 17642
rect 24669 17584 24674 17640
rect 24730 17584 26882 17640
rect 26938 17584 26943 17640
rect 24669 17582 26943 17584
rect 24669 17579 24735 17582
rect 26877 17579 26943 17582
rect 14273 17506 14339 17509
rect 18965 17506 19031 17509
rect 14273 17504 19031 17506
rect 14273 17448 14278 17504
rect 14334 17448 18970 17504
rect 19026 17448 19031 17504
rect 14273 17446 19031 17448
rect 14273 17443 14339 17446
rect 18965 17443 19031 17446
rect 22185 17506 22251 17509
rect 26049 17506 26115 17509
rect 22185 17504 26115 17506
rect 22185 17448 22190 17504
rect 22246 17448 26054 17504
rect 26110 17448 26115 17504
rect 22185 17446 26115 17448
rect 22185 17443 22251 17446
rect 26049 17443 26115 17446
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 11432 17440 11748 17441
rect 11432 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11748 17440
rect 11432 17375 11748 17376
rect 19206 17440 19522 17441
rect 19206 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19522 17440
rect 19206 17375 19522 17376
rect 26980 17440 27296 17441
rect 26980 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27296 17440
rect 26980 17375 27296 17376
rect 27429 17370 27495 17373
rect 28533 17370 28599 17373
rect 27429 17368 28599 17370
rect 27429 17312 27434 17368
rect 27490 17312 28538 17368
rect 28594 17312 28599 17368
rect 27429 17310 28599 17312
rect 27429 17307 27495 17310
rect 28533 17307 28599 17310
rect 10409 17234 10475 17237
rect 20253 17234 20319 17237
rect 10409 17232 20319 17234
rect 10409 17176 10414 17232
rect 10470 17176 20258 17232
rect 20314 17176 20319 17232
rect 10409 17174 20319 17176
rect 10409 17171 10475 17174
rect 20253 17171 20319 17174
rect 27981 17234 28047 17237
rect 28625 17234 28691 17237
rect 27981 17232 28691 17234
rect 27981 17176 27986 17232
rect 28042 17176 28630 17232
rect 28686 17176 28691 17232
rect 27981 17174 28691 17176
rect 27981 17171 28047 17174
rect 28625 17171 28691 17174
rect 6085 17098 6151 17101
rect 6453 17098 6519 17101
rect 11421 17098 11487 17101
rect 6085 17096 11487 17098
rect 6085 17040 6090 17096
rect 6146 17040 6458 17096
rect 6514 17040 11426 17096
rect 11482 17040 11487 17096
rect 6085 17038 11487 17040
rect 6085 17035 6151 17038
rect 6453 17035 6519 17038
rect 11421 17035 11487 17038
rect 24945 17098 25011 17101
rect 27889 17098 27955 17101
rect 24945 17096 27955 17098
rect 24945 17040 24950 17096
rect 25006 17040 27894 17096
rect 27950 17040 27955 17096
rect 24945 17038 27955 17040
rect 24945 17035 25011 17038
rect 27889 17035 27955 17038
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 12092 16896 12408 16897
rect 12092 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12408 16896
rect 12092 16831 12408 16832
rect 19866 16896 20182 16897
rect 19866 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20182 16896
rect 19866 16831 20182 16832
rect 27640 16896 27956 16897
rect 27640 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27956 16896
rect 27640 16831 27956 16832
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 11432 16352 11748 16353
rect 11432 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11748 16352
rect 11432 16287 11748 16288
rect 19206 16352 19522 16353
rect 19206 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19522 16352
rect 19206 16287 19522 16288
rect 26980 16352 27296 16353
rect 26980 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27296 16352
rect 26980 16287 27296 16288
rect 22001 16010 22067 16013
rect 27797 16010 27863 16013
rect 22001 16008 27863 16010
rect 22001 15952 22006 16008
rect 22062 15952 27802 16008
rect 27858 15952 27863 16008
rect 22001 15950 27863 15952
rect 22001 15947 22067 15950
rect 27797 15947 27863 15950
rect 23013 15874 23079 15877
rect 24209 15874 24275 15877
rect 25405 15874 25471 15877
rect 23013 15872 25471 15874
rect 23013 15816 23018 15872
rect 23074 15816 24214 15872
rect 24270 15816 25410 15872
rect 25466 15816 25471 15872
rect 23013 15814 25471 15816
rect 23013 15811 23079 15814
rect 24209 15811 24275 15814
rect 25405 15811 25471 15814
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 12092 15808 12408 15809
rect 12092 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12408 15808
rect 12092 15743 12408 15744
rect 19866 15808 20182 15809
rect 19866 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20182 15808
rect 19866 15743 20182 15744
rect 27640 15808 27956 15809
rect 27640 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27956 15808
rect 27640 15743 27956 15744
rect 21265 15602 21331 15605
rect 23933 15602 23999 15605
rect 21265 15600 23999 15602
rect 21265 15544 21270 15600
rect 21326 15544 23938 15600
rect 23994 15544 23999 15600
rect 21265 15542 23999 15544
rect 21265 15539 21331 15542
rect 23933 15539 23999 15542
rect 16481 15466 16547 15469
rect 18321 15466 18387 15469
rect 16481 15464 18387 15466
rect 16481 15408 16486 15464
rect 16542 15408 18326 15464
rect 18382 15408 18387 15464
rect 16481 15406 18387 15408
rect 16481 15403 16547 15406
rect 18321 15403 18387 15406
rect 21081 15466 21147 15469
rect 22921 15466 22987 15469
rect 21081 15464 22987 15466
rect 21081 15408 21086 15464
rect 21142 15408 22926 15464
rect 22982 15408 22987 15464
rect 21081 15406 22987 15408
rect 21081 15403 21147 15406
rect 22921 15403 22987 15406
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 11432 15264 11748 15265
rect 11432 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11748 15264
rect 11432 15199 11748 15200
rect 19206 15264 19522 15265
rect 19206 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19522 15264
rect 19206 15199 19522 15200
rect 26980 15264 27296 15265
rect 26980 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27296 15264
rect 26980 15199 27296 15200
rect 17217 15058 17283 15061
rect 21357 15058 21423 15061
rect 17217 15056 21423 15058
rect 17217 15000 17222 15056
rect 17278 15000 21362 15056
rect 21418 15000 21423 15056
rect 17217 14998 21423 15000
rect 17217 14995 17283 14998
rect 21357 14995 21423 14998
rect 24025 15058 24091 15061
rect 25865 15058 25931 15061
rect 24025 15056 25931 15058
rect 24025 15000 24030 15056
rect 24086 15000 25870 15056
rect 25926 15000 25931 15056
rect 24025 14998 25931 15000
rect 24025 14995 24091 14998
rect 25865 14995 25931 14998
rect 4981 14922 5047 14925
rect 18781 14922 18847 14925
rect 25313 14922 25379 14925
rect 4981 14920 5090 14922
rect 4981 14864 4986 14920
rect 5042 14864 5090 14920
rect 4981 14859 5090 14864
rect 18781 14920 25379 14922
rect 18781 14864 18786 14920
rect 18842 14864 25318 14920
rect 25374 14864 25379 14920
rect 18781 14862 25379 14864
rect 18781 14859 18847 14862
rect 25313 14859 25379 14862
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 5030 14653 5090 14859
rect 12092 14720 12408 14721
rect 12092 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12408 14720
rect 12092 14655 12408 14656
rect 19866 14720 20182 14721
rect 19866 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20182 14720
rect 19866 14655 20182 14656
rect 27640 14720 27956 14721
rect 27640 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27956 14720
rect 27640 14655 27956 14656
rect 4981 14648 5090 14653
rect 4981 14592 4986 14648
rect 5042 14592 5090 14648
rect 4981 14590 5090 14592
rect 28809 14650 28875 14653
rect 30557 14650 30623 14653
rect 28809 14648 30623 14650
rect 28809 14592 28814 14648
rect 28870 14592 30562 14648
rect 30618 14592 30623 14648
rect 28809 14590 30623 14592
rect 4981 14587 5047 14590
rect 28809 14587 28875 14590
rect 30557 14587 30623 14590
rect 16573 14514 16639 14517
rect 17309 14514 17375 14517
rect 30925 14514 30991 14517
rect 16573 14512 30991 14514
rect 16573 14456 16578 14512
rect 16634 14456 17314 14512
rect 17370 14456 30930 14512
rect 30986 14456 30991 14512
rect 16573 14454 30991 14456
rect 16573 14451 16639 14454
rect 17309 14451 17375 14454
rect 30925 14451 30991 14454
rect 5625 14378 5691 14381
rect 15009 14378 15075 14381
rect 5625 14376 15075 14378
rect 5625 14320 5630 14376
rect 5686 14320 15014 14376
rect 15070 14320 15075 14376
rect 5625 14318 15075 14320
rect 5625 14315 5691 14318
rect 15009 14315 15075 14318
rect 18045 14378 18111 14381
rect 24301 14378 24367 14381
rect 28809 14378 28875 14381
rect 18045 14376 24367 14378
rect 18045 14320 18050 14376
rect 18106 14320 24306 14376
rect 24362 14320 24367 14376
rect 18045 14318 24367 14320
rect 18045 14315 18111 14318
rect 24301 14315 24367 14318
rect 26742 14376 28875 14378
rect 26742 14320 28814 14376
rect 28870 14320 28875 14376
rect 26742 14318 28875 14320
rect 22277 14242 22343 14245
rect 26417 14242 26483 14245
rect 26742 14242 26802 14318
rect 28809 14315 28875 14318
rect 22277 14240 26802 14242
rect 22277 14184 22282 14240
rect 22338 14184 26422 14240
rect 26478 14184 26802 14240
rect 22277 14182 26802 14184
rect 22277 14179 22343 14182
rect 26417 14179 26483 14182
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 11432 14176 11748 14177
rect 11432 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11748 14176
rect 11432 14111 11748 14112
rect 19206 14176 19522 14177
rect 19206 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19522 14176
rect 19206 14111 19522 14112
rect 26980 14176 27296 14177
rect 26980 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27296 14176
rect 26980 14111 27296 14112
rect 21725 14106 21791 14109
rect 25221 14106 25287 14109
rect 21725 14104 25287 14106
rect 21725 14048 21730 14104
rect 21786 14048 25226 14104
rect 25282 14048 25287 14104
rect 21725 14046 25287 14048
rect 21725 14043 21791 14046
rect 25221 14043 25287 14046
rect 9949 13970 10015 13973
rect 13721 13970 13787 13973
rect 9949 13968 13787 13970
rect 9949 13912 9954 13968
rect 10010 13912 13726 13968
rect 13782 13912 13787 13968
rect 9949 13910 13787 13912
rect 9949 13907 10015 13910
rect 13721 13907 13787 13910
rect 19885 13970 19951 13973
rect 27337 13970 27403 13973
rect 19885 13968 27403 13970
rect 19885 13912 19890 13968
rect 19946 13912 27342 13968
rect 27398 13912 27403 13968
rect 19885 13910 27403 13912
rect 19885 13907 19951 13910
rect 27337 13907 27403 13910
rect 9489 13834 9555 13837
rect 13629 13834 13695 13837
rect 9489 13832 13695 13834
rect 9489 13776 9494 13832
rect 9550 13776 13634 13832
rect 13690 13776 13695 13832
rect 9489 13774 13695 13776
rect 9489 13771 9555 13774
rect 13629 13771 13695 13774
rect 19425 13834 19491 13837
rect 20529 13834 20595 13837
rect 21725 13834 21791 13837
rect 19425 13832 21791 13834
rect 19425 13776 19430 13832
rect 19486 13776 20534 13832
rect 20590 13776 21730 13832
rect 21786 13776 21791 13832
rect 19425 13774 21791 13776
rect 19425 13771 19491 13774
rect 20529 13771 20595 13774
rect 21725 13771 21791 13774
rect 22921 13834 22987 13837
rect 23381 13834 23447 13837
rect 24945 13834 25011 13837
rect 26969 13834 27035 13837
rect 28165 13834 28231 13837
rect 22921 13832 28231 13834
rect 22921 13776 22926 13832
rect 22982 13776 23386 13832
rect 23442 13776 24950 13832
rect 25006 13776 26974 13832
rect 27030 13776 28170 13832
rect 28226 13776 28231 13832
rect 22921 13774 28231 13776
rect 22921 13771 22987 13774
rect 23381 13771 23447 13774
rect 24945 13771 25011 13774
rect 26969 13771 27035 13774
rect 28165 13771 28231 13774
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 12092 13632 12408 13633
rect 12092 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12408 13632
rect 12092 13567 12408 13568
rect 19866 13632 20182 13633
rect 19866 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20182 13632
rect 19866 13567 20182 13568
rect 27640 13632 27956 13633
rect 27640 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27956 13632
rect 27640 13567 27956 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 11432 13088 11748 13089
rect 11432 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11748 13088
rect 11432 13023 11748 13024
rect 19206 13088 19522 13089
rect 19206 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19522 13088
rect 19206 13023 19522 13024
rect 26980 13088 27296 13089
rect 26980 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27296 13088
rect 26980 13023 27296 13024
rect 15101 12882 15167 12885
rect 18137 12882 18203 12885
rect 15101 12880 18203 12882
rect 15101 12824 15106 12880
rect 15162 12824 18142 12880
rect 18198 12824 18203 12880
rect 15101 12822 18203 12824
rect 15101 12819 15167 12822
rect 18137 12819 18203 12822
rect 12985 12746 13051 12749
rect 17309 12746 17375 12749
rect 12985 12744 17375 12746
rect 12985 12688 12990 12744
rect 13046 12688 17314 12744
rect 17370 12688 17375 12744
rect 12985 12686 17375 12688
rect 12985 12683 13051 12686
rect 17309 12683 17375 12686
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 12092 12544 12408 12545
rect 12092 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12408 12544
rect 12092 12479 12408 12480
rect 19866 12544 20182 12545
rect 19866 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20182 12544
rect 19866 12479 20182 12480
rect 27640 12544 27956 12545
rect 27640 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27956 12544
rect 27640 12479 27956 12480
rect 26233 12474 26299 12477
rect 26233 12472 26434 12474
rect 26233 12416 26238 12472
rect 26294 12416 26434 12472
rect 26233 12414 26434 12416
rect 26233 12411 26299 12414
rect 10542 12276 10548 12340
rect 10612 12338 10618 12340
rect 15561 12338 15627 12341
rect 10612 12336 15627 12338
rect 10612 12280 15566 12336
rect 15622 12280 15627 12336
rect 10612 12278 15627 12280
rect 10612 12276 10618 12278
rect 15561 12275 15627 12278
rect 19609 12338 19675 12341
rect 22553 12338 22619 12341
rect 23105 12338 23171 12341
rect 19609 12336 23171 12338
rect 19609 12280 19614 12336
rect 19670 12280 22558 12336
rect 22614 12280 23110 12336
rect 23166 12280 23171 12336
rect 19609 12278 23171 12280
rect 19609 12275 19675 12278
rect 22553 12275 22619 12278
rect 23105 12275 23171 12278
rect 20437 12202 20503 12205
rect 22277 12202 22343 12205
rect 22829 12202 22895 12205
rect 20437 12200 22895 12202
rect 20437 12144 20442 12200
rect 20498 12144 22282 12200
rect 22338 12144 22834 12200
rect 22890 12144 22895 12200
rect 20437 12142 22895 12144
rect 26374 12202 26434 12414
rect 26509 12202 26575 12205
rect 26374 12200 26575 12202
rect 26374 12144 26514 12200
rect 26570 12144 26575 12200
rect 26374 12142 26575 12144
rect 20437 12139 20503 12142
rect 22277 12139 22343 12142
rect 22829 12139 22895 12142
rect 26509 12139 26575 12142
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 11432 12000 11748 12001
rect 11432 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11748 12000
rect 11432 11935 11748 11936
rect 19206 12000 19522 12001
rect 19206 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19522 12000
rect 19206 11935 19522 11936
rect 26980 12000 27296 12001
rect 26980 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27296 12000
rect 26980 11935 27296 11936
rect 17861 11658 17927 11661
rect 28758 11658 28764 11660
rect 17861 11656 28764 11658
rect 17861 11600 17866 11656
rect 17922 11600 28764 11656
rect 17861 11598 28764 11600
rect 17861 11595 17927 11598
rect 28758 11596 28764 11598
rect 28828 11596 28834 11660
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 12092 11456 12408 11457
rect 12092 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12408 11456
rect 12092 11391 12408 11392
rect 19866 11456 20182 11457
rect 19866 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20182 11456
rect 19866 11391 20182 11392
rect 27640 11456 27956 11457
rect 27640 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27956 11456
rect 27640 11391 27956 11392
rect 19977 11250 20043 11253
rect 20294 11250 20300 11252
rect 19977 11248 20300 11250
rect 19977 11192 19982 11248
rect 20038 11192 20300 11248
rect 19977 11190 20300 11192
rect 19977 11187 20043 11190
rect 20294 11188 20300 11190
rect 20364 11188 20370 11252
rect 19333 11114 19399 11117
rect 26049 11114 26115 11117
rect 19333 11112 26115 11114
rect 19333 11056 19338 11112
rect 19394 11056 26054 11112
rect 26110 11056 26115 11112
rect 19333 11054 26115 11056
rect 19333 11051 19399 11054
rect 26049 11051 26115 11054
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 11432 10912 11748 10913
rect 11432 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11748 10912
rect 11432 10847 11748 10848
rect 19206 10912 19522 10913
rect 19206 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19522 10912
rect 19206 10847 19522 10848
rect 26980 10912 27296 10913
rect 26980 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27296 10912
rect 26980 10847 27296 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 12092 10368 12408 10369
rect 12092 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12408 10368
rect 12092 10303 12408 10304
rect 19866 10368 20182 10369
rect 19866 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20182 10368
rect 19866 10303 20182 10304
rect 27640 10368 27956 10369
rect 27640 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27956 10368
rect 27640 10303 27956 10304
rect 15009 10162 15075 10165
rect 16941 10162 17007 10165
rect 15009 10160 17007 10162
rect 15009 10104 15014 10160
rect 15070 10104 16946 10160
rect 17002 10104 17007 10160
rect 15009 10102 17007 10104
rect 15009 10099 15075 10102
rect 16941 10099 17007 10102
rect 22737 10162 22803 10165
rect 25865 10162 25931 10165
rect 27429 10162 27495 10165
rect 22737 10160 27495 10162
rect 22737 10104 22742 10160
rect 22798 10104 25870 10160
rect 25926 10104 27434 10160
rect 27490 10104 27495 10160
rect 22737 10102 27495 10104
rect 22737 10099 22803 10102
rect 25865 10099 25931 10102
rect 27429 10099 27495 10102
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 11432 9824 11748 9825
rect 11432 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11748 9824
rect 11432 9759 11748 9760
rect 19206 9824 19522 9825
rect 19206 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19522 9824
rect 19206 9759 19522 9760
rect 26980 9824 27296 9825
rect 26980 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27296 9824
rect 26980 9759 27296 9760
rect 19333 9482 19399 9485
rect 20529 9482 20595 9485
rect 24209 9482 24275 9485
rect 19333 9480 24275 9482
rect 19333 9424 19338 9480
rect 19394 9424 20534 9480
rect 20590 9424 24214 9480
rect 24270 9424 24275 9480
rect 19333 9422 24275 9424
rect 19333 9419 19399 9422
rect 20529 9419 20595 9422
rect 24209 9419 24275 9422
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 12092 9280 12408 9281
rect 12092 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12408 9280
rect 12092 9215 12408 9216
rect 19866 9280 20182 9281
rect 19866 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20182 9280
rect 19866 9215 20182 9216
rect 27640 9280 27956 9281
rect 27640 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27956 9280
rect 27640 9215 27956 9216
rect 22185 9074 22251 9077
rect 23657 9074 23723 9077
rect 22185 9072 23723 9074
rect 22185 9016 22190 9072
rect 22246 9016 23662 9072
rect 23718 9016 23723 9072
rect 22185 9014 23723 9016
rect 22185 9011 22251 9014
rect 23657 9011 23723 9014
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 11432 8736 11748 8737
rect 11432 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11748 8736
rect 11432 8671 11748 8672
rect 19206 8736 19522 8737
rect 19206 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19522 8736
rect 19206 8671 19522 8672
rect 26980 8736 27296 8737
rect 26980 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27296 8736
rect 26980 8671 27296 8672
rect 22277 8666 22343 8669
rect 22921 8666 22987 8669
rect 22277 8664 22987 8666
rect 22277 8608 22282 8664
rect 22338 8608 22926 8664
rect 22982 8608 22987 8664
rect 22277 8606 22987 8608
rect 22277 8603 22343 8606
rect 22921 8603 22987 8606
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 12092 8192 12408 8193
rect 12092 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12408 8192
rect 12092 8127 12408 8128
rect 19866 8192 20182 8193
rect 19866 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20182 8192
rect 19866 8127 20182 8128
rect 27640 8192 27956 8193
rect 27640 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27956 8192
rect 27640 8127 27956 8128
rect 15009 8122 15075 8125
rect 15653 8122 15719 8125
rect 17585 8122 17651 8125
rect 15009 8120 17651 8122
rect 15009 8064 15014 8120
rect 15070 8064 15658 8120
rect 15714 8064 17590 8120
rect 17646 8064 17651 8120
rect 15009 8062 17651 8064
rect 15009 8059 15075 8062
rect 15653 8059 15719 8062
rect 17585 8059 17651 8062
rect 9857 7986 9923 7989
rect 13997 7986 14063 7989
rect 9857 7984 14063 7986
rect 9857 7928 9862 7984
rect 9918 7928 14002 7984
rect 14058 7928 14063 7984
rect 9857 7926 14063 7928
rect 9857 7923 9923 7926
rect 13997 7923 14063 7926
rect 14549 7986 14615 7989
rect 15561 7986 15627 7989
rect 16849 7986 16915 7989
rect 14549 7984 16915 7986
rect 14549 7928 14554 7984
rect 14610 7928 15566 7984
rect 15622 7928 16854 7984
rect 16910 7928 16915 7984
rect 14549 7926 16915 7928
rect 14549 7923 14615 7926
rect 15561 7923 15627 7926
rect 16849 7923 16915 7926
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 11432 7648 11748 7649
rect 11432 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11748 7648
rect 11432 7583 11748 7584
rect 19206 7648 19522 7649
rect 19206 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19522 7648
rect 19206 7583 19522 7584
rect 26980 7648 27296 7649
rect 26980 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27296 7648
rect 26980 7583 27296 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 12092 7104 12408 7105
rect 12092 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12408 7104
rect 12092 7039 12408 7040
rect 19866 7104 20182 7105
rect 19866 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20182 7104
rect 19866 7039 20182 7040
rect 27640 7104 27956 7105
rect 27640 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27956 7104
rect 27640 7039 27956 7040
rect 19006 6972 19012 7036
rect 19076 7034 19082 7036
rect 19149 7034 19215 7037
rect 19076 7032 19215 7034
rect 19076 6976 19154 7032
rect 19210 6976 19215 7032
rect 19076 6974 19215 6976
rect 19076 6972 19082 6974
rect 19149 6971 19215 6974
rect 19241 6898 19307 6901
rect 18830 6896 19307 6898
rect 18830 6840 19246 6896
rect 19302 6840 19307 6896
rect 18830 6838 19307 6840
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 11432 6560 11748 6561
rect 11432 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11748 6560
rect 11432 6495 11748 6496
rect 18830 6354 18890 6838
rect 19241 6835 19307 6838
rect 18965 6762 19031 6765
rect 30189 6762 30255 6765
rect 18965 6760 30255 6762
rect 18965 6704 18970 6760
rect 19026 6704 30194 6760
rect 30250 6704 30255 6760
rect 18965 6702 30255 6704
rect 18965 6699 19031 6702
rect 30189 6699 30255 6702
rect 19206 6560 19522 6561
rect 19206 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19522 6560
rect 19206 6495 19522 6496
rect 26980 6560 27296 6561
rect 26980 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27296 6560
rect 26980 6495 27296 6496
rect 22277 6490 22343 6493
rect 23105 6490 23171 6493
rect 22277 6488 23171 6490
rect 22277 6432 22282 6488
rect 22338 6432 23110 6488
rect 23166 6432 23171 6488
rect 22277 6430 23171 6432
rect 22277 6427 22343 6430
rect 23105 6427 23171 6430
rect 19149 6354 19215 6357
rect 18830 6352 19215 6354
rect 18830 6296 19154 6352
rect 19210 6296 19215 6352
rect 18830 6294 19215 6296
rect 19149 6291 19215 6294
rect 19977 6354 20043 6357
rect 25497 6354 25563 6357
rect 19977 6352 25563 6354
rect 19977 6296 19982 6352
rect 20038 6296 25502 6352
rect 25558 6296 25563 6352
rect 19977 6294 25563 6296
rect 19977 6291 20043 6294
rect 25497 6291 25563 6294
rect 18137 6218 18203 6221
rect 19793 6218 19859 6221
rect 18137 6216 19859 6218
rect 18137 6160 18142 6216
rect 18198 6160 19798 6216
rect 19854 6160 19859 6216
rect 18137 6158 19859 6160
rect 18137 6155 18203 6158
rect 19793 6155 19859 6158
rect 22001 6218 22067 6221
rect 26693 6218 26759 6221
rect 22001 6216 26759 6218
rect 22001 6160 22006 6216
rect 22062 6160 26698 6216
rect 26754 6160 26759 6216
rect 22001 6158 26759 6160
rect 22001 6155 22067 6158
rect 26693 6155 26759 6158
rect 18965 6082 19031 6085
rect 19333 6082 19399 6085
rect 18965 6080 19399 6082
rect 18965 6024 18970 6080
rect 19026 6024 19338 6080
rect 19394 6024 19399 6080
rect 18965 6022 19399 6024
rect 18965 6019 19031 6022
rect 19333 6019 19399 6022
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 12092 6016 12408 6017
rect 12092 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12408 6016
rect 12092 5951 12408 5952
rect 19866 6016 20182 6017
rect 19866 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20182 6016
rect 19866 5951 20182 5952
rect 27640 6016 27956 6017
rect 27640 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27956 6016
rect 27640 5951 27956 5952
rect 19057 5948 19123 5949
rect 19006 5884 19012 5948
rect 19076 5946 19123 5948
rect 21725 5946 21791 5949
rect 23289 5946 23355 5949
rect 19076 5944 19168 5946
rect 19118 5888 19168 5944
rect 19076 5886 19168 5888
rect 21725 5944 23355 5946
rect 21725 5888 21730 5944
rect 21786 5888 23294 5944
rect 23350 5888 23355 5944
rect 21725 5886 23355 5888
rect 19076 5884 19123 5886
rect 19057 5883 19123 5884
rect 21725 5883 21791 5886
rect 23289 5883 23355 5886
rect 19701 5810 19767 5813
rect 25405 5810 25471 5813
rect 19701 5808 25471 5810
rect 19701 5752 19706 5808
rect 19762 5752 25410 5808
rect 25466 5752 25471 5808
rect 19701 5750 25471 5752
rect 19701 5747 19767 5750
rect 25405 5747 25471 5750
rect 15929 5674 15995 5677
rect 25037 5674 25103 5677
rect 15929 5672 25103 5674
rect 15929 5616 15934 5672
rect 15990 5616 25042 5672
rect 25098 5616 25103 5672
rect 15929 5614 25103 5616
rect 15929 5611 15995 5614
rect 25037 5611 25103 5614
rect 20621 5538 20687 5541
rect 24577 5538 24643 5541
rect 20621 5536 24643 5538
rect 20621 5480 20626 5536
rect 20682 5480 24582 5536
rect 24638 5480 24643 5536
rect 20621 5478 24643 5480
rect 20621 5475 20687 5478
rect 24577 5475 24643 5478
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 11432 5472 11748 5473
rect 11432 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11748 5472
rect 11432 5407 11748 5408
rect 19206 5472 19522 5473
rect 19206 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19522 5472
rect 19206 5407 19522 5408
rect 26980 5472 27296 5473
rect 26980 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27296 5472
rect 26980 5407 27296 5408
rect 12525 5402 12591 5405
rect 18965 5402 19031 5405
rect 12525 5400 19031 5402
rect 12525 5344 12530 5400
rect 12586 5344 18970 5400
rect 19026 5344 19031 5400
rect 12525 5342 19031 5344
rect 12525 5339 12591 5342
rect 18965 5339 19031 5342
rect 21173 5402 21239 5405
rect 23657 5402 23723 5405
rect 21173 5400 23723 5402
rect 21173 5344 21178 5400
rect 21234 5344 23662 5400
rect 23718 5344 23723 5400
rect 21173 5342 23723 5344
rect 21173 5339 21239 5342
rect 23657 5339 23723 5342
rect 21357 5266 21423 5269
rect 22737 5266 22803 5269
rect 21357 5264 22803 5266
rect 21357 5208 21362 5264
rect 21418 5208 22742 5264
rect 22798 5208 22803 5264
rect 21357 5206 22803 5208
rect 21357 5203 21423 5206
rect 22737 5203 22803 5206
rect 23197 5130 23263 5133
rect 24577 5130 24643 5133
rect 23197 5128 24643 5130
rect 23197 5072 23202 5128
rect 23258 5072 24582 5128
rect 24638 5072 24643 5128
rect 23197 5070 24643 5072
rect 23197 5067 23263 5070
rect 24577 5067 24643 5070
rect 22645 4994 22711 4997
rect 23933 4994 23999 4997
rect 22645 4992 23999 4994
rect 22645 4936 22650 4992
rect 22706 4936 23938 4992
rect 23994 4936 23999 4992
rect 22645 4934 23999 4936
rect 22645 4931 22711 4934
rect 23933 4931 23999 4934
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 12092 4928 12408 4929
rect 12092 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12408 4928
rect 12092 4863 12408 4864
rect 19866 4928 20182 4929
rect 19866 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20182 4928
rect 19866 4863 20182 4864
rect 27640 4928 27956 4929
rect 27640 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27956 4928
rect 27640 4863 27956 4864
rect 1761 4586 1827 4589
rect 2681 4586 2747 4589
rect 1761 4584 2747 4586
rect 1761 4528 1766 4584
rect 1822 4528 2686 4584
rect 2742 4528 2747 4584
rect 1761 4526 2747 4528
rect 1761 4523 1827 4526
rect 2681 4523 2747 4526
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 11432 4384 11748 4385
rect 11432 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11748 4384
rect 11432 4319 11748 4320
rect 19206 4384 19522 4385
rect 19206 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19522 4384
rect 19206 4319 19522 4320
rect 26980 4384 27296 4385
rect 26980 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27296 4384
rect 26980 4319 27296 4320
rect 14549 4178 14615 4181
rect 18229 4178 18295 4181
rect 14549 4176 18295 4178
rect 14549 4120 14554 4176
rect 14610 4120 18234 4176
rect 18290 4120 18295 4176
rect 14549 4118 18295 4120
rect 14549 4115 14615 4118
rect 18229 4115 18295 4118
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 12092 3840 12408 3841
rect 12092 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12408 3840
rect 12092 3775 12408 3776
rect 19866 3840 20182 3841
rect 19866 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20182 3840
rect 19866 3775 20182 3776
rect 27640 3840 27956 3841
rect 27640 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27956 3840
rect 27640 3775 27956 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 11432 3296 11748 3297
rect 11432 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11748 3296
rect 11432 3231 11748 3232
rect 19206 3296 19522 3297
rect 19206 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19522 3296
rect 19206 3231 19522 3232
rect 26980 3296 27296 3297
rect 26980 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27296 3296
rect 26980 3231 27296 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 12092 2752 12408 2753
rect 12092 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12408 2752
rect 12092 2687 12408 2688
rect 19866 2752 20182 2753
rect 19866 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20182 2752
rect 19866 2687 20182 2688
rect 27640 2752 27956 2753
rect 27640 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27956 2752
rect 27640 2687 27956 2688
rect 21633 2546 21699 2549
rect 22645 2546 22711 2549
rect 21633 2544 22711 2546
rect 21633 2488 21638 2544
rect 21694 2488 22650 2544
rect 22706 2488 22711 2544
rect 21633 2486 22711 2488
rect 21633 2483 21699 2486
rect 22645 2483 22711 2486
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 11432 2208 11748 2209
rect 11432 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11748 2208
rect 11432 2143 11748 2144
rect 19206 2208 19522 2209
rect 19206 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19522 2208
rect 19206 2143 19522 2144
rect 26980 2208 27296 2209
rect 26980 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27296 2208
rect 26980 2143 27296 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 12092 1664 12408 1665
rect 12092 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12408 1664
rect 12092 1599 12408 1600
rect 19866 1664 20182 1665
rect 19866 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20182 1664
rect 19866 1599 20182 1600
rect 27640 1664 27956 1665
rect 27640 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27956 1664
rect 27640 1599 27956 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 11432 1120 11748 1121
rect 11432 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11748 1120
rect 11432 1055 11748 1056
rect 19206 1120 19522 1121
rect 19206 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19522 1120
rect 19206 1055 19522 1056
rect 26980 1120 27296 1121
rect 26980 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27296 1120
rect 26980 1055 27296 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 12092 576 12408 577
rect 12092 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12408 576
rect 12092 511 12408 512
rect 19866 576 20182 577
rect 19866 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20182 576
rect 19866 511 20182 512
rect 27640 576 27956 577
rect 27640 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27956 576
rect 27640 511 27956 512
<< via3 >>
rect 11652 21932 11716 21996
rect 12204 21992 12268 21996
rect 12204 21936 12254 21992
rect 12254 21936 12268 21992
rect 12204 21932 12268 21936
rect 24348 21992 24412 21996
rect 24348 21936 24398 21992
rect 24398 21936 24412 21992
rect 24348 21932 24412 21936
rect 27108 21932 27172 21996
rect 27660 21992 27724 21996
rect 27660 21936 27710 21992
rect 27710 21936 27724 21992
rect 27660 21932 27724 21936
rect 7236 21796 7300 21860
rect 21588 21796 21652 21860
rect 23796 21856 23860 21860
rect 23796 21800 23846 21856
rect 23846 21800 23860 21856
rect 23796 21796 23860 21800
rect 26004 21796 26068 21860
rect 26556 21796 26620 21860
rect 28212 21856 28276 21860
rect 28212 21800 28262 21856
rect 28262 21800 28276 21856
rect 28212 21796 28276 21800
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 11438 21788 11502 21792
rect 11438 21732 11442 21788
rect 11442 21732 11498 21788
rect 11498 21732 11502 21788
rect 11438 21728 11502 21732
rect 11518 21788 11582 21792
rect 11518 21732 11522 21788
rect 11522 21732 11578 21788
rect 11578 21732 11582 21788
rect 11518 21728 11582 21732
rect 11598 21788 11662 21792
rect 11598 21732 11602 21788
rect 11602 21732 11658 21788
rect 11658 21732 11662 21788
rect 11598 21728 11662 21732
rect 11678 21788 11742 21792
rect 11678 21732 11682 21788
rect 11682 21732 11738 21788
rect 11738 21732 11742 21788
rect 11678 21728 11742 21732
rect 19212 21788 19276 21792
rect 19212 21732 19216 21788
rect 19216 21732 19272 21788
rect 19272 21732 19276 21788
rect 19212 21728 19276 21732
rect 19292 21788 19356 21792
rect 19292 21732 19296 21788
rect 19296 21732 19352 21788
rect 19352 21732 19356 21788
rect 19292 21728 19356 21732
rect 19372 21788 19436 21792
rect 19372 21732 19376 21788
rect 19376 21732 19432 21788
rect 19432 21732 19436 21788
rect 19372 21728 19436 21732
rect 19452 21788 19516 21792
rect 19452 21732 19456 21788
rect 19456 21732 19512 21788
rect 19512 21732 19516 21788
rect 19452 21728 19516 21732
rect 26986 21788 27050 21792
rect 26986 21732 26990 21788
rect 26990 21732 27046 21788
rect 27046 21732 27050 21788
rect 26986 21728 27050 21732
rect 27066 21788 27130 21792
rect 27066 21732 27070 21788
rect 27070 21732 27126 21788
rect 27126 21732 27130 21788
rect 27066 21728 27130 21732
rect 27146 21788 27210 21792
rect 27146 21732 27150 21788
rect 27150 21732 27206 21788
rect 27206 21732 27210 21788
rect 27146 21728 27210 21732
rect 27226 21788 27290 21792
rect 27226 21732 27230 21788
rect 27230 21732 27286 21788
rect 27286 21732 27290 21788
rect 27226 21728 27290 21732
rect 6132 21720 6196 21724
rect 6132 21664 6146 21720
rect 6146 21664 6196 21720
rect 6132 21660 6196 21664
rect 7788 21660 7852 21724
rect 8340 21720 8404 21724
rect 8340 21664 8390 21720
rect 8390 21664 8404 21720
rect 8340 21660 8404 21664
rect 12756 21660 12820 21724
rect 24900 21660 24964 21724
rect 25452 21584 25516 21588
rect 25452 21528 25502 21584
rect 25502 21528 25516 21584
rect 25452 21524 25516 21528
rect 17172 21388 17236 21452
rect 9444 21252 9508 21316
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 12098 21244 12162 21248
rect 12098 21188 12102 21244
rect 12102 21188 12158 21244
rect 12158 21188 12162 21244
rect 12098 21184 12162 21188
rect 12178 21244 12242 21248
rect 12178 21188 12182 21244
rect 12182 21188 12238 21244
rect 12238 21188 12242 21244
rect 12178 21184 12242 21188
rect 12258 21244 12322 21248
rect 12258 21188 12262 21244
rect 12262 21188 12318 21244
rect 12318 21188 12322 21244
rect 12258 21184 12322 21188
rect 12338 21244 12402 21248
rect 12338 21188 12342 21244
rect 12342 21188 12398 21244
rect 12398 21188 12402 21244
rect 12338 21184 12402 21188
rect 19872 21244 19936 21248
rect 19872 21188 19876 21244
rect 19876 21188 19932 21244
rect 19932 21188 19936 21244
rect 19872 21184 19936 21188
rect 19952 21244 20016 21248
rect 19952 21188 19956 21244
rect 19956 21188 20012 21244
rect 20012 21188 20016 21244
rect 19952 21184 20016 21188
rect 20032 21244 20096 21248
rect 20032 21188 20036 21244
rect 20036 21188 20092 21244
rect 20092 21188 20096 21244
rect 20032 21184 20096 21188
rect 20112 21244 20176 21248
rect 20112 21188 20116 21244
rect 20116 21188 20172 21244
rect 20172 21188 20176 21244
rect 20112 21184 20176 21188
rect 27646 21244 27710 21248
rect 27646 21188 27650 21244
rect 27650 21188 27706 21244
rect 27706 21188 27710 21244
rect 27646 21184 27710 21188
rect 27726 21244 27790 21248
rect 27726 21188 27730 21244
rect 27730 21188 27786 21244
rect 27786 21188 27790 21244
rect 27726 21184 27790 21188
rect 27806 21244 27870 21248
rect 27806 21188 27810 21244
rect 27810 21188 27866 21244
rect 27866 21188 27870 21244
rect 27806 21184 27870 21188
rect 27886 21244 27950 21248
rect 27886 21188 27890 21244
rect 27890 21188 27946 21244
rect 27946 21188 27950 21244
rect 27886 21184 27950 21188
rect 8892 21116 8956 21180
rect 9996 21116 10060 21180
rect 18276 21116 18340 21180
rect 18828 20980 18892 21044
rect 16068 20844 16132 20908
rect 15516 20708 15580 20772
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 11438 20700 11502 20704
rect 11438 20644 11442 20700
rect 11442 20644 11498 20700
rect 11498 20644 11502 20700
rect 11438 20640 11502 20644
rect 11518 20700 11582 20704
rect 11518 20644 11522 20700
rect 11522 20644 11578 20700
rect 11578 20644 11582 20700
rect 11518 20640 11582 20644
rect 11598 20700 11662 20704
rect 11598 20644 11602 20700
rect 11602 20644 11658 20700
rect 11658 20644 11662 20700
rect 11598 20640 11662 20644
rect 11678 20700 11742 20704
rect 11678 20644 11682 20700
rect 11682 20644 11738 20700
rect 11738 20644 11742 20700
rect 11678 20640 11742 20644
rect 19212 20700 19276 20704
rect 19212 20644 19216 20700
rect 19216 20644 19272 20700
rect 19272 20644 19276 20700
rect 19212 20640 19276 20644
rect 19292 20700 19356 20704
rect 19292 20644 19296 20700
rect 19296 20644 19352 20700
rect 19352 20644 19356 20700
rect 19292 20640 19356 20644
rect 19372 20700 19436 20704
rect 19372 20644 19376 20700
rect 19376 20644 19432 20700
rect 19432 20644 19436 20700
rect 19372 20640 19436 20644
rect 19452 20700 19516 20704
rect 19452 20644 19456 20700
rect 19456 20644 19512 20700
rect 19512 20644 19516 20700
rect 19452 20640 19516 20644
rect 26986 20700 27050 20704
rect 26986 20644 26990 20700
rect 26990 20644 27046 20700
rect 27046 20644 27050 20700
rect 26986 20640 27050 20644
rect 27066 20700 27130 20704
rect 27066 20644 27070 20700
rect 27070 20644 27126 20700
rect 27126 20644 27130 20700
rect 27066 20640 27130 20644
rect 27146 20700 27210 20704
rect 27146 20644 27150 20700
rect 27150 20644 27206 20700
rect 27206 20644 27210 20700
rect 27146 20640 27210 20644
rect 27226 20700 27290 20704
rect 27226 20644 27230 20700
rect 27230 20644 27286 20700
rect 27286 20644 27290 20700
rect 27226 20640 27290 20644
rect 11100 20632 11164 20636
rect 11100 20576 11114 20632
rect 11114 20576 11164 20632
rect 11100 20572 11164 20576
rect 13308 20632 13372 20636
rect 13308 20576 13322 20632
rect 13322 20576 13372 20632
rect 13308 20572 13372 20576
rect 14964 20572 15028 20636
rect 16620 20572 16684 20636
rect 6684 20360 6748 20364
rect 6684 20304 6734 20360
rect 6734 20304 6748 20360
rect 6684 20300 6748 20304
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 12098 20156 12162 20160
rect 12098 20100 12102 20156
rect 12102 20100 12158 20156
rect 12158 20100 12162 20156
rect 12098 20096 12162 20100
rect 12178 20156 12242 20160
rect 12178 20100 12182 20156
rect 12182 20100 12238 20156
rect 12238 20100 12242 20156
rect 12178 20096 12242 20100
rect 12258 20156 12322 20160
rect 12258 20100 12262 20156
rect 12262 20100 12318 20156
rect 12318 20100 12322 20156
rect 12258 20096 12322 20100
rect 12338 20156 12402 20160
rect 12338 20100 12342 20156
rect 12342 20100 12398 20156
rect 12398 20100 12402 20156
rect 12338 20096 12402 20100
rect 19872 20156 19936 20160
rect 19872 20100 19876 20156
rect 19876 20100 19932 20156
rect 19932 20100 19936 20156
rect 19872 20096 19936 20100
rect 19952 20156 20016 20160
rect 19952 20100 19956 20156
rect 19956 20100 20012 20156
rect 20012 20100 20016 20156
rect 19952 20096 20016 20100
rect 20032 20156 20096 20160
rect 20032 20100 20036 20156
rect 20036 20100 20092 20156
rect 20092 20100 20096 20156
rect 20032 20096 20096 20100
rect 20112 20156 20176 20160
rect 20112 20100 20116 20156
rect 20116 20100 20172 20156
rect 20172 20100 20176 20156
rect 20112 20096 20176 20100
rect 27646 20156 27710 20160
rect 27646 20100 27650 20156
rect 27650 20100 27706 20156
rect 27706 20100 27710 20156
rect 27646 20096 27710 20100
rect 27726 20156 27790 20160
rect 27726 20100 27730 20156
rect 27730 20100 27786 20156
rect 27786 20100 27790 20156
rect 27726 20096 27790 20100
rect 27806 20156 27870 20160
rect 27806 20100 27810 20156
rect 27810 20100 27866 20156
rect 27866 20100 27870 20156
rect 27806 20096 27870 20100
rect 27886 20156 27950 20160
rect 27886 20100 27890 20156
rect 27890 20100 27946 20156
rect 27946 20100 27950 20156
rect 27886 20096 27950 20100
rect 17724 19892 17788 19956
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 11438 19612 11502 19616
rect 11438 19556 11442 19612
rect 11442 19556 11498 19612
rect 11498 19556 11502 19612
rect 11438 19552 11502 19556
rect 11518 19612 11582 19616
rect 11518 19556 11522 19612
rect 11522 19556 11578 19612
rect 11578 19556 11582 19612
rect 11518 19552 11582 19556
rect 11598 19612 11662 19616
rect 11598 19556 11602 19612
rect 11602 19556 11658 19612
rect 11658 19556 11662 19612
rect 11598 19552 11662 19556
rect 11678 19612 11742 19616
rect 11678 19556 11682 19612
rect 11682 19556 11738 19612
rect 11738 19556 11742 19612
rect 11678 19552 11742 19556
rect 19212 19612 19276 19616
rect 19212 19556 19216 19612
rect 19216 19556 19272 19612
rect 19272 19556 19276 19612
rect 19212 19552 19276 19556
rect 19292 19612 19356 19616
rect 19292 19556 19296 19612
rect 19296 19556 19352 19612
rect 19352 19556 19356 19612
rect 19292 19552 19356 19556
rect 19372 19612 19436 19616
rect 19372 19556 19376 19612
rect 19376 19556 19432 19612
rect 19432 19556 19436 19612
rect 19372 19552 19436 19556
rect 19452 19612 19516 19616
rect 19452 19556 19456 19612
rect 19456 19556 19512 19612
rect 19512 19556 19516 19612
rect 19452 19552 19516 19556
rect 26986 19612 27050 19616
rect 26986 19556 26990 19612
rect 26990 19556 27046 19612
rect 27046 19556 27050 19612
rect 26986 19552 27050 19556
rect 27066 19612 27130 19616
rect 27066 19556 27070 19612
rect 27070 19556 27126 19612
rect 27126 19556 27130 19612
rect 27066 19552 27130 19556
rect 27146 19612 27210 19616
rect 27146 19556 27150 19612
rect 27150 19556 27206 19612
rect 27206 19556 27210 19612
rect 27146 19552 27210 19556
rect 27226 19612 27290 19616
rect 27226 19556 27230 19612
rect 27230 19556 27286 19612
rect 27286 19556 27290 19612
rect 27226 19552 27290 19556
rect 14412 19212 14476 19276
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 12098 19068 12162 19072
rect 12098 19012 12102 19068
rect 12102 19012 12158 19068
rect 12158 19012 12162 19068
rect 12098 19008 12162 19012
rect 12178 19068 12242 19072
rect 12178 19012 12182 19068
rect 12182 19012 12238 19068
rect 12238 19012 12242 19068
rect 12178 19008 12242 19012
rect 12258 19068 12322 19072
rect 12258 19012 12262 19068
rect 12262 19012 12318 19068
rect 12318 19012 12322 19068
rect 12258 19008 12322 19012
rect 12338 19068 12402 19072
rect 12338 19012 12342 19068
rect 12342 19012 12398 19068
rect 12398 19012 12402 19068
rect 12338 19008 12402 19012
rect 19872 19068 19936 19072
rect 19872 19012 19876 19068
rect 19876 19012 19932 19068
rect 19932 19012 19936 19068
rect 19872 19008 19936 19012
rect 19952 19068 20016 19072
rect 19952 19012 19956 19068
rect 19956 19012 20012 19068
rect 20012 19012 20016 19068
rect 19952 19008 20016 19012
rect 20032 19068 20096 19072
rect 20032 19012 20036 19068
rect 20036 19012 20092 19068
rect 20092 19012 20096 19068
rect 20032 19008 20096 19012
rect 20112 19068 20176 19072
rect 20112 19012 20116 19068
rect 20116 19012 20172 19068
rect 20172 19012 20176 19068
rect 20112 19008 20176 19012
rect 27646 19068 27710 19072
rect 27646 19012 27650 19068
rect 27650 19012 27706 19068
rect 27706 19012 27710 19068
rect 27646 19008 27710 19012
rect 27726 19068 27790 19072
rect 27726 19012 27730 19068
rect 27730 19012 27786 19068
rect 27786 19012 27790 19068
rect 27726 19008 27790 19012
rect 27806 19068 27870 19072
rect 27806 19012 27810 19068
rect 27810 19012 27866 19068
rect 27866 19012 27870 19068
rect 27806 19008 27870 19012
rect 27886 19068 27950 19072
rect 27886 19012 27890 19068
rect 27890 19012 27946 19068
rect 27946 19012 27950 19068
rect 27886 19008 27950 19012
rect 13860 18804 13924 18868
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 11438 18524 11502 18528
rect 11438 18468 11442 18524
rect 11442 18468 11498 18524
rect 11498 18468 11502 18524
rect 11438 18464 11502 18468
rect 11518 18524 11582 18528
rect 11518 18468 11522 18524
rect 11522 18468 11578 18524
rect 11578 18468 11582 18524
rect 11518 18464 11582 18468
rect 11598 18524 11662 18528
rect 11598 18468 11602 18524
rect 11602 18468 11658 18524
rect 11658 18468 11662 18524
rect 11598 18464 11662 18468
rect 11678 18524 11742 18528
rect 11678 18468 11682 18524
rect 11682 18468 11738 18524
rect 11738 18468 11742 18524
rect 11678 18464 11742 18468
rect 19212 18524 19276 18528
rect 19212 18468 19216 18524
rect 19216 18468 19272 18524
rect 19272 18468 19276 18524
rect 19212 18464 19276 18468
rect 19292 18524 19356 18528
rect 19292 18468 19296 18524
rect 19296 18468 19352 18524
rect 19352 18468 19356 18524
rect 19292 18464 19356 18468
rect 19372 18524 19436 18528
rect 19372 18468 19376 18524
rect 19376 18468 19432 18524
rect 19432 18468 19436 18524
rect 19372 18464 19436 18468
rect 19452 18524 19516 18528
rect 19452 18468 19456 18524
rect 19456 18468 19512 18524
rect 19512 18468 19516 18524
rect 19452 18464 19516 18468
rect 26986 18524 27050 18528
rect 26986 18468 26990 18524
rect 26990 18468 27046 18524
rect 27046 18468 27050 18524
rect 26986 18464 27050 18468
rect 27066 18524 27130 18528
rect 27066 18468 27070 18524
rect 27070 18468 27126 18524
rect 27126 18468 27130 18524
rect 27066 18464 27130 18468
rect 27146 18524 27210 18528
rect 27146 18468 27150 18524
rect 27150 18468 27206 18524
rect 27206 18468 27210 18524
rect 27146 18464 27210 18468
rect 27226 18524 27290 18528
rect 27226 18468 27230 18524
rect 27230 18468 27286 18524
rect 27286 18468 27290 18524
rect 27226 18464 27290 18468
rect 20300 18124 20364 18188
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 12098 17980 12162 17984
rect 12098 17924 12102 17980
rect 12102 17924 12158 17980
rect 12158 17924 12162 17980
rect 12098 17920 12162 17924
rect 12178 17980 12242 17984
rect 12178 17924 12182 17980
rect 12182 17924 12238 17980
rect 12238 17924 12242 17980
rect 12178 17920 12242 17924
rect 12258 17980 12322 17984
rect 12258 17924 12262 17980
rect 12262 17924 12318 17980
rect 12318 17924 12322 17980
rect 12258 17920 12322 17924
rect 12338 17980 12402 17984
rect 12338 17924 12342 17980
rect 12342 17924 12398 17980
rect 12398 17924 12402 17980
rect 12338 17920 12402 17924
rect 19872 17980 19936 17984
rect 19872 17924 19876 17980
rect 19876 17924 19932 17980
rect 19932 17924 19936 17980
rect 19872 17920 19936 17924
rect 19952 17980 20016 17984
rect 19952 17924 19956 17980
rect 19956 17924 20012 17980
rect 20012 17924 20016 17980
rect 19952 17920 20016 17924
rect 20032 17980 20096 17984
rect 20032 17924 20036 17980
rect 20036 17924 20092 17980
rect 20092 17924 20096 17980
rect 20032 17920 20096 17924
rect 20112 17980 20176 17984
rect 20112 17924 20116 17980
rect 20116 17924 20172 17980
rect 20172 17924 20176 17980
rect 20112 17920 20176 17924
rect 27646 17980 27710 17984
rect 27646 17924 27650 17980
rect 27650 17924 27706 17980
rect 27706 17924 27710 17980
rect 27646 17920 27710 17924
rect 27726 17980 27790 17984
rect 27726 17924 27730 17980
rect 27730 17924 27786 17980
rect 27786 17924 27790 17980
rect 27726 17920 27790 17924
rect 27806 17980 27870 17984
rect 27806 17924 27810 17980
rect 27810 17924 27866 17980
rect 27866 17924 27870 17980
rect 27806 17920 27870 17924
rect 27886 17980 27950 17984
rect 27886 17924 27890 17980
rect 27890 17924 27946 17980
rect 27946 17924 27950 17980
rect 27886 17920 27950 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 11438 17436 11502 17440
rect 11438 17380 11442 17436
rect 11442 17380 11498 17436
rect 11498 17380 11502 17436
rect 11438 17376 11502 17380
rect 11518 17436 11582 17440
rect 11518 17380 11522 17436
rect 11522 17380 11578 17436
rect 11578 17380 11582 17436
rect 11518 17376 11582 17380
rect 11598 17436 11662 17440
rect 11598 17380 11602 17436
rect 11602 17380 11658 17436
rect 11658 17380 11662 17436
rect 11598 17376 11662 17380
rect 11678 17436 11742 17440
rect 11678 17380 11682 17436
rect 11682 17380 11738 17436
rect 11738 17380 11742 17436
rect 11678 17376 11742 17380
rect 19212 17436 19276 17440
rect 19212 17380 19216 17436
rect 19216 17380 19272 17436
rect 19272 17380 19276 17436
rect 19212 17376 19276 17380
rect 19292 17436 19356 17440
rect 19292 17380 19296 17436
rect 19296 17380 19352 17436
rect 19352 17380 19356 17436
rect 19292 17376 19356 17380
rect 19372 17436 19436 17440
rect 19372 17380 19376 17436
rect 19376 17380 19432 17436
rect 19432 17380 19436 17436
rect 19372 17376 19436 17380
rect 19452 17436 19516 17440
rect 19452 17380 19456 17436
rect 19456 17380 19512 17436
rect 19512 17380 19516 17436
rect 19452 17376 19516 17380
rect 26986 17436 27050 17440
rect 26986 17380 26990 17436
rect 26990 17380 27046 17436
rect 27046 17380 27050 17436
rect 26986 17376 27050 17380
rect 27066 17436 27130 17440
rect 27066 17380 27070 17436
rect 27070 17380 27126 17436
rect 27126 17380 27130 17436
rect 27066 17376 27130 17380
rect 27146 17436 27210 17440
rect 27146 17380 27150 17436
rect 27150 17380 27206 17436
rect 27206 17380 27210 17436
rect 27146 17376 27210 17380
rect 27226 17436 27290 17440
rect 27226 17380 27230 17436
rect 27230 17380 27286 17436
rect 27286 17380 27290 17436
rect 27226 17376 27290 17380
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 12098 16892 12162 16896
rect 12098 16836 12102 16892
rect 12102 16836 12158 16892
rect 12158 16836 12162 16892
rect 12098 16832 12162 16836
rect 12178 16892 12242 16896
rect 12178 16836 12182 16892
rect 12182 16836 12238 16892
rect 12238 16836 12242 16892
rect 12178 16832 12242 16836
rect 12258 16892 12322 16896
rect 12258 16836 12262 16892
rect 12262 16836 12318 16892
rect 12318 16836 12322 16892
rect 12258 16832 12322 16836
rect 12338 16892 12402 16896
rect 12338 16836 12342 16892
rect 12342 16836 12398 16892
rect 12398 16836 12402 16892
rect 12338 16832 12402 16836
rect 19872 16892 19936 16896
rect 19872 16836 19876 16892
rect 19876 16836 19932 16892
rect 19932 16836 19936 16892
rect 19872 16832 19936 16836
rect 19952 16892 20016 16896
rect 19952 16836 19956 16892
rect 19956 16836 20012 16892
rect 20012 16836 20016 16892
rect 19952 16832 20016 16836
rect 20032 16892 20096 16896
rect 20032 16836 20036 16892
rect 20036 16836 20092 16892
rect 20092 16836 20096 16892
rect 20032 16832 20096 16836
rect 20112 16892 20176 16896
rect 20112 16836 20116 16892
rect 20116 16836 20172 16892
rect 20172 16836 20176 16892
rect 20112 16832 20176 16836
rect 27646 16892 27710 16896
rect 27646 16836 27650 16892
rect 27650 16836 27706 16892
rect 27706 16836 27710 16892
rect 27646 16832 27710 16836
rect 27726 16892 27790 16896
rect 27726 16836 27730 16892
rect 27730 16836 27786 16892
rect 27786 16836 27790 16892
rect 27726 16832 27790 16836
rect 27806 16892 27870 16896
rect 27806 16836 27810 16892
rect 27810 16836 27866 16892
rect 27866 16836 27870 16892
rect 27806 16832 27870 16836
rect 27886 16892 27950 16896
rect 27886 16836 27890 16892
rect 27890 16836 27946 16892
rect 27946 16836 27950 16892
rect 27886 16832 27950 16836
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 11438 16348 11502 16352
rect 11438 16292 11442 16348
rect 11442 16292 11498 16348
rect 11498 16292 11502 16348
rect 11438 16288 11502 16292
rect 11518 16348 11582 16352
rect 11518 16292 11522 16348
rect 11522 16292 11578 16348
rect 11578 16292 11582 16348
rect 11518 16288 11582 16292
rect 11598 16348 11662 16352
rect 11598 16292 11602 16348
rect 11602 16292 11658 16348
rect 11658 16292 11662 16348
rect 11598 16288 11662 16292
rect 11678 16348 11742 16352
rect 11678 16292 11682 16348
rect 11682 16292 11738 16348
rect 11738 16292 11742 16348
rect 11678 16288 11742 16292
rect 19212 16348 19276 16352
rect 19212 16292 19216 16348
rect 19216 16292 19272 16348
rect 19272 16292 19276 16348
rect 19212 16288 19276 16292
rect 19292 16348 19356 16352
rect 19292 16292 19296 16348
rect 19296 16292 19352 16348
rect 19352 16292 19356 16348
rect 19292 16288 19356 16292
rect 19372 16348 19436 16352
rect 19372 16292 19376 16348
rect 19376 16292 19432 16348
rect 19432 16292 19436 16348
rect 19372 16288 19436 16292
rect 19452 16348 19516 16352
rect 19452 16292 19456 16348
rect 19456 16292 19512 16348
rect 19512 16292 19516 16348
rect 19452 16288 19516 16292
rect 26986 16348 27050 16352
rect 26986 16292 26990 16348
rect 26990 16292 27046 16348
rect 27046 16292 27050 16348
rect 26986 16288 27050 16292
rect 27066 16348 27130 16352
rect 27066 16292 27070 16348
rect 27070 16292 27126 16348
rect 27126 16292 27130 16348
rect 27066 16288 27130 16292
rect 27146 16348 27210 16352
rect 27146 16292 27150 16348
rect 27150 16292 27206 16348
rect 27206 16292 27210 16348
rect 27146 16288 27210 16292
rect 27226 16348 27290 16352
rect 27226 16292 27230 16348
rect 27230 16292 27286 16348
rect 27286 16292 27290 16348
rect 27226 16288 27290 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 12098 15804 12162 15808
rect 12098 15748 12102 15804
rect 12102 15748 12158 15804
rect 12158 15748 12162 15804
rect 12098 15744 12162 15748
rect 12178 15804 12242 15808
rect 12178 15748 12182 15804
rect 12182 15748 12238 15804
rect 12238 15748 12242 15804
rect 12178 15744 12242 15748
rect 12258 15804 12322 15808
rect 12258 15748 12262 15804
rect 12262 15748 12318 15804
rect 12318 15748 12322 15804
rect 12258 15744 12322 15748
rect 12338 15804 12402 15808
rect 12338 15748 12342 15804
rect 12342 15748 12398 15804
rect 12398 15748 12402 15804
rect 12338 15744 12402 15748
rect 19872 15804 19936 15808
rect 19872 15748 19876 15804
rect 19876 15748 19932 15804
rect 19932 15748 19936 15804
rect 19872 15744 19936 15748
rect 19952 15804 20016 15808
rect 19952 15748 19956 15804
rect 19956 15748 20012 15804
rect 20012 15748 20016 15804
rect 19952 15744 20016 15748
rect 20032 15804 20096 15808
rect 20032 15748 20036 15804
rect 20036 15748 20092 15804
rect 20092 15748 20096 15804
rect 20032 15744 20096 15748
rect 20112 15804 20176 15808
rect 20112 15748 20116 15804
rect 20116 15748 20172 15804
rect 20172 15748 20176 15804
rect 20112 15744 20176 15748
rect 27646 15804 27710 15808
rect 27646 15748 27650 15804
rect 27650 15748 27706 15804
rect 27706 15748 27710 15804
rect 27646 15744 27710 15748
rect 27726 15804 27790 15808
rect 27726 15748 27730 15804
rect 27730 15748 27786 15804
rect 27786 15748 27790 15804
rect 27726 15744 27790 15748
rect 27806 15804 27870 15808
rect 27806 15748 27810 15804
rect 27810 15748 27866 15804
rect 27866 15748 27870 15804
rect 27806 15744 27870 15748
rect 27886 15804 27950 15808
rect 27886 15748 27890 15804
rect 27890 15748 27946 15804
rect 27946 15748 27950 15804
rect 27886 15744 27950 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 11438 15260 11502 15264
rect 11438 15204 11442 15260
rect 11442 15204 11498 15260
rect 11498 15204 11502 15260
rect 11438 15200 11502 15204
rect 11518 15260 11582 15264
rect 11518 15204 11522 15260
rect 11522 15204 11578 15260
rect 11578 15204 11582 15260
rect 11518 15200 11582 15204
rect 11598 15260 11662 15264
rect 11598 15204 11602 15260
rect 11602 15204 11658 15260
rect 11658 15204 11662 15260
rect 11598 15200 11662 15204
rect 11678 15260 11742 15264
rect 11678 15204 11682 15260
rect 11682 15204 11738 15260
rect 11738 15204 11742 15260
rect 11678 15200 11742 15204
rect 19212 15260 19276 15264
rect 19212 15204 19216 15260
rect 19216 15204 19272 15260
rect 19272 15204 19276 15260
rect 19212 15200 19276 15204
rect 19292 15260 19356 15264
rect 19292 15204 19296 15260
rect 19296 15204 19352 15260
rect 19352 15204 19356 15260
rect 19292 15200 19356 15204
rect 19372 15260 19436 15264
rect 19372 15204 19376 15260
rect 19376 15204 19432 15260
rect 19432 15204 19436 15260
rect 19372 15200 19436 15204
rect 19452 15260 19516 15264
rect 19452 15204 19456 15260
rect 19456 15204 19512 15260
rect 19512 15204 19516 15260
rect 19452 15200 19516 15204
rect 26986 15260 27050 15264
rect 26986 15204 26990 15260
rect 26990 15204 27046 15260
rect 27046 15204 27050 15260
rect 26986 15200 27050 15204
rect 27066 15260 27130 15264
rect 27066 15204 27070 15260
rect 27070 15204 27126 15260
rect 27126 15204 27130 15260
rect 27066 15200 27130 15204
rect 27146 15260 27210 15264
rect 27146 15204 27150 15260
rect 27150 15204 27206 15260
rect 27206 15204 27210 15260
rect 27146 15200 27210 15204
rect 27226 15260 27290 15264
rect 27226 15204 27230 15260
rect 27230 15204 27286 15260
rect 27286 15204 27290 15260
rect 27226 15200 27290 15204
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 12098 14716 12162 14720
rect 12098 14660 12102 14716
rect 12102 14660 12158 14716
rect 12158 14660 12162 14716
rect 12098 14656 12162 14660
rect 12178 14716 12242 14720
rect 12178 14660 12182 14716
rect 12182 14660 12238 14716
rect 12238 14660 12242 14716
rect 12178 14656 12242 14660
rect 12258 14716 12322 14720
rect 12258 14660 12262 14716
rect 12262 14660 12318 14716
rect 12318 14660 12322 14716
rect 12258 14656 12322 14660
rect 12338 14716 12402 14720
rect 12338 14660 12342 14716
rect 12342 14660 12398 14716
rect 12398 14660 12402 14716
rect 12338 14656 12402 14660
rect 19872 14716 19936 14720
rect 19872 14660 19876 14716
rect 19876 14660 19932 14716
rect 19932 14660 19936 14716
rect 19872 14656 19936 14660
rect 19952 14716 20016 14720
rect 19952 14660 19956 14716
rect 19956 14660 20012 14716
rect 20012 14660 20016 14716
rect 19952 14656 20016 14660
rect 20032 14716 20096 14720
rect 20032 14660 20036 14716
rect 20036 14660 20092 14716
rect 20092 14660 20096 14716
rect 20032 14656 20096 14660
rect 20112 14716 20176 14720
rect 20112 14660 20116 14716
rect 20116 14660 20172 14716
rect 20172 14660 20176 14716
rect 20112 14656 20176 14660
rect 27646 14716 27710 14720
rect 27646 14660 27650 14716
rect 27650 14660 27706 14716
rect 27706 14660 27710 14716
rect 27646 14656 27710 14660
rect 27726 14716 27790 14720
rect 27726 14660 27730 14716
rect 27730 14660 27786 14716
rect 27786 14660 27790 14716
rect 27726 14656 27790 14660
rect 27806 14716 27870 14720
rect 27806 14660 27810 14716
rect 27810 14660 27866 14716
rect 27866 14660 27870 14716
rect 27806 14656 27870 14660
rect 27886 14716 27950 14720
rect 27886 14660 27890 14716
rect 27890 14660 27946 14716
rect 27946 14660 27950 14716
rect 27886 14656 27950 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 11438 14172 11502 14176
rect 11438 14116 11442 14172
rect 11442 14116 11498 14172
rect 11498 14116 11502 14172
rect 11438 14112 11502 14116
rect 11518 14172 11582 14176
rect 11518 14116 11522 14172
rect 11522 14116 11578 14172
rect 11578 14116 11582 14172
rect 11518 14112 11582 14116
rect 11598 14172 11662 14176
rect 11598 14116 11602 14172
rect 11602 14116 11658 14172
rect 11658 14116 11662 14172
rect 11598 14112 11662 14116
rect 11678 14172 11742 14176
rect 11678 14116 11682 14172
rect 11682 14116 11738 14172
rect 11738 14116 11742 14172
rect 11678 14112 11742 14116
rect 19212 14172 19276 14176
rect 19212 14116 19216 14172
rect 19216 14116 19272 14172
rect 19272 14116 19276 14172
rect 19212 14112 19276 14116
rect 19292 14172 19356 14176
rect 19292 14116 19296 14172
rect 19296 14116 19352 14172
rect 19352 14116 19356 14172
rect 19292 14112 19356 14116
rect 19372 14172 19436 14176
rect 19372 14116 19376 14172
rect 19376 14116 19432 14172
rect 19432 14116 19436 14172
rect 19372 14112 19436 14116
rect 19452 14172 19516 14176
rect 19452 14116 19456 14172
rect 19456 14116 19512 14172
rect 19512 14116 19516 14172
rect 19452 14112 19516 14116
rect 26986 14172 27050 14176
rect 26986 14116 26990 14172
rect 26990 14116 27046 14172
rect 27046 14116 27050 14172
rect 26986 14112 27050 14116
rect 27066 14172 27130 14176
rect 27066 14116 27070 14172
rect 27070 14116 27126 14172
rect 27126 14116 27130 14172
rect 27066 14112 27130 14116
rect 27146 14172 27210 14176
rect 27146 14116 27150 14172
rect 27150 14116 27206 14172
rect 27206 14116 27210 14172
rect 27146 14112 27210 14116
rect 27226 14172 27290 14176
rect 27226 14116 27230 14172
rect 27230 14116 27286 14172
rect 27286 14116 27290 14172
rect 27226 14112 27290 14116
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 12098 13628 12162 13632
rect 12098 13572 12102 13628
rect 12102 13572 12158 13628
rect 12158 13572 12162 13628
rect 12098 13568 12162 13572
rect 12178 13628 12242 13632
rect 12178 13572 12182 13628
rect 12182 13572 12238 13628
rect 12238 13572 12242 13628
rect 12178 13568 12242 13572
rect 12258 13628 12322 13632
rect 12258 13572 12262 13628
rect 12262 13572 12318 13628
rect 12318 13572 12322 13628
rect 12258 13568 12322 13572
rect 12338 13628 12402 13632
rect 12338 13572 12342 13628
rect 12342 13572 12398 13628
rect 12398 13572 12402 13628
rect 12338 13568 12402 13572
rect 19872 13628 19936 13632
rect 19872 13572 19876 13628
rect 19876 13572 19932 13628
rect 19932 13572 19936 13628
rect 19872 13568 19936 13572
rect 19952 13628 20016 13632
rect 19952 13572 19956 13628
rect 19956 13572 20012 13628
rect 20012 13572 20016 13628
rect 19952 13568 20016 13572
rect 20032 13628 20096 13632
rect 20032 13572 20036 13628
rect 20036 13572 20092 13628
rect 20092 13572 20096 13628
rect 20032 13568 20096 13572
rect 20112 13628 20176 13632
rect 20112 13572 20116 13628
rect 20116 13572 20172 13628
rect 20172 13572 20176 13628
rect 20112 13568 20176 13572
rect 27646 13628 27710 13632
rect 27646 13572 27650 13628
rect 27650 13572 27706 13628
rect 27706 13572 27710 13628
rect 27646 13568 27710 13572
rect 27726 13628 27790 13632
rect 27726 13572 27730 13628
rect 27730 13572 27786 13628
rect 27786 13572 27790 13628
rect 27726 13568 27790 13572
rect 27806 13628 27870 13632
rect 27806 13572 27810 13628
rect 27810 13572 27866 13628
rect 27866 13572 27870 13628
rect 27806 13568 27870 13572
rect 27886 13628 27950 13632
rect 27886 13572 27890 13628
rect 27890 13572 27946 13628
rect 27946 13572 27950 13628
rect 27886 13568 27950 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 11438 13084 11502 13088
rect 11438 13028 11442 13084
rect 11442 13028 11498 13084
rect 11498 13028 11502 13084
rect 11438 13024 11502 13028
rect 11518 13084 11582 13088
rect 11518 13028 11522 13084
rect 11522 13028 11578 13084
rect 11578 13028 11582 13084
rect 11518 13024 11582 13028
rect 11598 13084 11662 13088
rect 11598 13028 11602 13084
rect 11602 13028 11658 13084
rect 11658 13028 11662 13084
rect 11598 13024 11662 13028
rect 11678 13084 11742 13088
rect 11678 13028 11682 13084
rect 11682 13028 11738 13084
rect 11738 13028 11742 13084
rect 11678 13024 11742 13028
rect 19212 13084 19276 13088
rect 19212 13028 19216 13084
rect 19216 13028 19272 13084
rect 19272 13028 19276 13084
rect 19212 13024 19276 13028
rect 19292 13084 19356 13088
rect 19292 13028 19296 13084
rect 19296 13028 19352 13084
rect 19352 13028 19356 13084
rect 19292 13024 19356 13028
rect 19372 13084 19436 13088
rect 19372 13028 19376 13084
rect 19376 13028 19432 13084
rect 19432 13028 19436 13084
rect 19372 13024 19436 13028
rect 19452 13084 19516 13088
rect 19452 13028 19456 13084
rect 19456 13028 19512 13084
rect 19512 13028 19516 13084
rect 19452 13024 19516 13028
rect 26986 13084 27050 13088
rect 26986 13028 26990 13084
rect 26990 13028 27046 13084
rect 27046 13028 27050 13084
rect 26986 13024 27050 13028
rect 27066 13084 27130 13088
rect 27066 13028 27070 13084
rect 27070 13028 27126 13084
rect 27126 13028 27130 13084
rect 27066 13024 27130 13028
rect 27146 13084 27210 13088
rect 27146 13028 27150 13084
rect 27150 13028 27206 13084
rect 27206 13028 27210 13084
rect 27146 13024 27210 13028
rect 27226 13084 27290 13088
rect 27226 13028 27230 13084
rect 27230 13028 27286 13084
rect 27286 13028 27290 13084
rect 27226 13024 27290 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 12098 12540 12162 12544
rect 12098 12484 12102 12540
rect 12102 12484 12158 12540
rect 12158 12484 12162 12540
rect 12098 12480 12162 12484
rect 12178 12540 12242 12544
rect 12178 12484 12182 12540
rect 12182 12484 12238 12540
rect 12238 12484 12242 12540
rect 12178 12480 12242 12484
rect 12258 12540 12322 12544
rect 12258 12484 12262 12540
rect 12262 12484 12318 12540
rect 12318 12484 12322 12540
rect 12258 12480 12322 12484
rect 12338 12540 12402 12544
rect 12338 12484 12342 12540
rect 12342 12484 12398 12540
rect 12398 12484 12402 12540
rect 12338 12480 12402 12484
rect 19872 12540 19936 12544
rect 19872 12484 19876 12540
rect 19876 12484 19932 12540
rect 19932 12484 19936 12540
rect 19872 12480 19936 12484
rect 19952 12540 20016 12544
rect 19952 12484 19956 12540
rect 19956 12484 20012 12540
rect 20012 12484 20016 12540
rect 19952 12480 20016 12484
rect 20032 12540 20096 12544
rect 20032 12484 20036 12540
rect 20036 12484 20092 12540
rect 20092 12484 20096 12540
rect 20032 12480 20096 12484
rect 20112 12540 20176 12544
rect 20112 12484 20116 12540
rect 20116 12484 20172 12540
rect 20172 12484 20176 12540
rect 20112 12480 20176 12484
rect 27646 12540 27710 12544
rect 27646 12484 27650 12540
rect 27650 12484 27706 12540
rect 27706 12484 27710 12540
rect 27646 12480 27710 12484
rect 27726 12540 27790 12544
rect 27726 12484 27730 12540
rect 27730 12484 27786 12540
rect 27786 12484 27790 12540
rect 27726 12480 27790 12484
rect 27806 12540 27870 12544
rect 27806 12484 27810 12540
rect 27810 12484 27866 12540
rect 27866 12484 27870 12540
rect 27806 12480 27870 12484
rect 27886 12540 27950 12544
rect 27886 12484 27890 12540
rect 27890 12484 27946 12540
rect 27946 12484 27950 12540
rect 27886 12480 27950 12484
rect 10548 12276 10612 12340
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 11438 11996 11502 12000
rect 11438 11940 11442 11996
rect 11442 11940 11498 11996
rect 11498 11940 11502 11996
rect 11438 11936 11502 11940
rect 11518 11996 11582 12000
rect 11518 11940 11522 11996
rect 11522 11940 11578 11996
rect 11578 11940 11582 11996
rect 11518 11936 11582 11940
rect 11598 11996 11662 12000
rect 11598 11940 11602 11996
rect 11602 11940 11658 11996
rect 11658 11940 11662 11996
rect 11598 11936 11662 11940
rect 11678 11996 11742 12000
rect 11678 11940 11682 11996
rect 11682 11940 11738 11996
rect 11738 11940 11742 11996
rect 11678 11936 11742 11940
rect 19212 11996 19276 12000
rect 19212 11940 19216 11996
rect 19216 11940 19272 11996
rect 19272 11940 19276 11996
rect 19212 11936 19276 11940
rect 19292 11996 19356 12000
rect 19292 11940 19296 11996
rect 19296 11940 19352 11996
rect 19352 11940 19356 11996
rect 19292 11936 19356 11940
rect 19372 11996 19436 12000
rect 19372 11940 19376 11996
rect 19376 11940 19432 11996
rect 19432 11940 19436 11996
rect 19372 11936 19436 11940
rect 19452 11996 19516 12000
rect 19452 11940 19456 11996
rect 19456 11940 19512 11996
rect 19512 11940 19516 11996
rect 19452 11936 19516 11940
rect 26986 11996 27050 12000
rect 26986 11940 26990 11996
rect 26990 11940 27046 11996
rect 27046 11940 27050 11996
rect 26986 11936 27050 11940
rect 27066 11996 27130 12000
rect 27066 11940 27070 11996
rect 27070 11940 27126 11996
rect 27126 11940 27130 11996
rect 27066 11936 27130 11940
rect 27146 11996 27210 12000
rect 27146 11940 27150 11996
rect 27150 11940 27206 11996
rect 27206 11940 27210 11996
rect 27146 11936 27210 11940
rect 27226 11996 27290 12000
rect 27226 11940 27230 11996
rect 27230 11940 27286 11996
rect 27286 11940 27290 11996
rect 27226 11936 27290 11940
rect 28764 11596 28828 11660
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 12098 11452 12162 11456
rect 12098 11396 12102 11452
rect 12102 11396 12158 11452
rect 12158 11396 12162 11452
rect 12098 11392 12162 11396
rect 12178 11452 12242 11456
rect 12178 11396 12182 11452
rect 12182 11396 12238 11452
rect 12238 11396 12242 11452
rect 12178 11392 12242 11396
rect 12258 11452 12322 11456
rect 12258 11396 12262 11452
rect 12262 11396 12318 11452
rect 12318 11396 12322 11452
rect 12258 11392 12322 11396
rect 12338 11452 12402 11456
rect 12338 11396 12342 11452
rect 12342 11396 12398 11452
rect 12398 11396 12402 11452
rect 12338 11392 12402 11396
rect 19872 11452 19936 11456
rect 19872 11396 19876 11452
rect 19876 11396 19932 11452
rect 19932 11396 19936 11452
rect 19872 11392 19936 11396
rect 19952 11452 20016 11456
rect 19952 11396 19956 11452
rect 19956 11396 20012 11452
rect 20012 11396 20016 11452
rect 19952 11392 20016 11396
rect 20032 11452 20096 11456
rect 20032 11396 20036 11452
rect 20036 11396 20092 11452
rect 20092 11396 20096 11452
rect 20032 11392 20096 11396
rect 20112 11452 20176 11456
rect 20112 11396 20116 11452
rect 20116 11396 20172 11452
rect 20172 11396 20176 11452
rect 20112 11392 20176 11396
rect 27646 11452 27710 11456
rect 27646 11396 27650 11452
rect 27650 11396 27706 11452
rect 27706 11396 27710 11452
rect 27646 11392 27710 11396
rect 27726 11452 27790 11456
rect 27726 11396 27730 11452
rect 27730 11396 27786 11452
rect 27786 11396 27790 11452
rect 27726 11392 27790 11396
rect 27806 11452 27870 11456
rect 27806 11396 27810 11452
rect 27810 11396 27866 11452
rect 27866 11396 27870 11452
rect 27806 11392 27870 11396
rect 27886 11452 27950 11456
rect 27886 11396 27890 11452
rect 27890 11396 27946 11452
rect 27946 11396 27950 11452
rect 27886 11392 27950 11396
rect 20300 11188 20364 11252
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 11438 10908 11502 10912
rect 11438 10852 11442 10908
rect 11442 10852 11498 10908
rect 11498 10852 11502 10908
rect 11438 10848 11502 10852
rect 11518 10908 11582 10912
rect 11518 10852 11522 10908
rect 11522 10852 11578 10908
rect 11578 10852 11582 10908
rect 11518 10848 11582 10852
rect 11598 10908 11662 10912
rect 11598 10852 11602 10908
rect 11602 10852 11658 10908
rect 11658 10852 11662 10908
rect 11598 10848 11662 10852
rect 11678 10908 11742 10912
rect 11678 10852 11682 10908
rect 11682 10852 11738 10908
rect 11738 10852 11742 10908
rect 11678 10848 11742 10852
rect 19212 10908 19276 10912
rect 19212 10852 19216 10908
rect 19216 10852 19272 10908
rect 19272 10852 19276 10908
rect 19212 10848 19276 10852
rect 19292 10908 19356 10912
rect 19292 10852 19296 10908
rect 19296 10852 19352 10908
rect 19352 10852 19356 10908
rect 19292 10848 19356 10852
rect 19372 10908 19436 10912
rect 19372 10852 19376 10908
rect 19376 10852 19432 10908
rect 19432 10852 19436 10908
rect 19372 10848 19436 10852
rect 19452 10908 19516 10912
rect 19452 10852 19456 10908
rect 19456 10852 19512 10908
rect 19512 10852 19516 10908
rect 19452 10848 19516 10852
rect 26986 10908 27050 10912
rect 26986 10852 26990 10908
rect 26990 10852 27046 10908
rect 27046 10852 27050 10908
rect 26986 10848 27050 10852
rect 27066 10908 27130 10912
rect 27066 10852 27070 10908
rect 27070 10852 27126 10908
rect 27126 10852 27130 10908
rect 27066 10848 27130 10852
rect 27146 10908 27210 10912
rect 27146 10852 27150 10908
rect 27150 10852 27206 10908
rect 27206 10852 27210 10908
rect 27146 10848 27210 10852
rect 27226 10908 27290 10912
rect 27226 10852 27230 10908
rect 27230 10852 27286 10908
rect 27286 10852 27290 10908
rect 27226 10848 27290 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 12098 10364 12162 10368
rect 12098 10308 12102 10364
rect 12102 10308 12158 10364
rect 12158 10308 12162 10364
rect 12098 10304 12162 10308
rect 12178 10364 12242 10368
rect 12178 10308 12182 10364
rect 12182 10308 12238 10364
rect 12238 10308 12242 10364
rect 12178 10304 12242 10308
rect 12258 10364 12322 10368
rect 12258 10308 12262 10364
rect 12262 10308 12318 10364
rect 12318 10308 12322 10364
rect 12258 10304 12322 10308
rect 12338 10364 12402 10368
rect 12338 10308 12342 10364
rect 12342 10308 12398 10364
rect 12398 10308 12402 10364
rect 12338 10304 12402 10308
rect 19872 10364 19936 10368
rect 19872 10308 19876 10364
rect 19876 10308 19932 10364
rect 19932 10308 19936 10364
rect 19872 10304 19936 10308
rect 19952 10364 20016 10368
rect 19952 10308 19956 10364
rect 19956 10308 20012 10364
rect 20012 10308 20016 10364
rect 19952 10304 20016 10308
rect 20032 10364 20096 10368
rect 20032 10308 20036 10364
rect 20036 10308 20092 10364
rect 20092 10308 20096 10364
rect 20032 10304 20096 10308
rect 20112 10364 20176 10368
rect 20112 10308 20116 10364
rect 20116 10308 20172 10364
rect 20172 10308 20176 10364
rect 20112 10304 20176 10308
rect 27646 10364 27710 10368
rect 27646 10308 27650 10364
rect 27650 10308 27706 10364
rect 27706 10308 27710 10364
rect 27646 10304 27710 10308
rect 27726 10364 27790 10368
rect 27726 10308 27730 10364
rect 27730 10308 27786 10364
rect 27786 10308 27790 10364
rect 27726 10304 27790 10308
rect 27806 10364 27870 10368
rect 27806 10308 27810 10364
rect 27810 10308 27866 10364
rect 27866 10308 27870 10364
rect 27806 10304 27870 10308
rect 27886 10364 27950 10368
rect 27886 10308 27890 10364
rect 27890 10308 27946 10364
rect 27946 10308 27950 10364
rect 27886 10304 27950 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 11438 9820 11502 9824
rect 11438 9764 11442 9820
rect 11442 9764 11498 9820
rect 11498 9764 11502 9820
rect 11438 9760 11502 9764
rect 11518 9820 11582 9824
rect 11518 9764 11522 9820
rect 11522 9764 11578 9820
rect 11578 9764 11582 9820
rect 11518 9760 11582 9764
rect 11598 9820 11662 9824
rect 11598 9764 11602 9820
rect 11602 9764 11658 9820
rect 11658 9764 11662 9820
rect 11598 9760 11662 9764
rect 11678 9820 11742 9824
rect 11678 9764 11682 9820
rect 11682 9764 11738 9820
rect 11738 9764 11742 9820
rect 11678 9760 11742 9764
rect 19212 9820 19276 9824
rect 19212 9764 19216 9820
rect 19216 9764 19272 9820
rect 19272 9764 19276 9820
rect 19212 9760 19276 9764
rect 19292 9820 19356 9824
rect 19292 9764 19296 9820
rect 19296 9764 19352 9820
rect 19352 9764 19356 9820
rect 19292 9760 19356 9764
rect 19372 9820 19436 9824
rect 19372 9764 19376 9820
rect 19376 9764 19432 9820
rect 19432 9764 19436 9820
rect 19372 9760 19436 9764
rect 19452 9820 19516 9824
rect 19452 9764 19456 9820
rect 19456 9764 19512 9820
rect 19512 9764 19516 9820
rect 19452 9760 19516 9764
rect 26986 9820 27050 9824
rect 26986 9764 26990 9820
rect 26990 9764 27046 9820
rect 27046 9764 27050 9820
rect 26986 9760 27050 9764
rect 27066 9820 27130 9824
rect 27066 9764 27070 9820
rect 27070 9764 27126 9820
rect 27126 9764 27130 9820
rect 27066 9760 27130 9764
rect 27146 9820 27210 9824
rect 27146 9764 27150 9820
rect 27150 9764 27206 9820
rect 27206 9764 27210 9820
rect 27146 9760 27210 9764
rect 27226 9820 27290 9824
rect 27226 9764 27230 9820
rect 27230 9764 27286 9820
rect 27286 9764 27290 9820
rect 27226 9760 27290 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 12098 9276 12162 9280
rect 12098 9220 12102 9276
rect 12102 9220 12158 9276
rect 12158 9220 12162 9276
rect 12098 9216 12162 9220
rect 12178 9276 12242 9280
rect 12178 9220 12182 9276
rect 12182 9220 12238 9276
rect 12238 9220 12242 9276
rect 12178 9216 12242 9220
rect 12258 9276 12322 9280
rect 12258 9220 12262 9276
rect 12262 9220 12318 9276
rect 12318 9220 12322 9276
rect 12258 9216 12322 9220
rect 12338 9276 12402 9280
rect 12338 9220 12342 9276
rect 12342 9220 12398 9276
rect 12398 9220 12402 9276
rect 12338 9216 12402 9220
rect 19872 9276 19936 9280
rect 19872 9220 19876 9276
rect 19876 9220 19932 9276
rect 19932 9220 19936 9276
rect 19872 9216 19936 9220
rect 19952 9276 20016 9280
rect 19952 9220 19956 9276
rect 19956 9220 20012 9276
rect 20012 9220 20016 9276
rect 19952 9216 20016 9220
rect 20032 9276 20096 9280
rect 20032 9220 20036 9276
rect 20036 9220 20092 9276
rect 20092 9220 20096 9276
rect 20032 9216 20096 9220
rect 20112 9276 20176 9280
rect 20112 9220 20116 9276
rect 20116 9220 20172 9276
rect 20172 9220 20176 9276
rect 20112 9216 20176 9220
rect 27646 9276 27710 9280
rect 27646 9220 27650 9276
rect 27650 9220 27706 9276
rect 27706 9220 27710 9276
rect 27646 9216 27710 9220
rect 27726 9276 27790 9280
rect 27726 9220 27730 9276
rect 27730 9220 27786 9276
rect 27786 9220 27790 9276
rect 27726 9216 27790 9220
rect 27806 9276 27870 9280
rect 27806 9220 27810 9276
rect 27810 9220 27866 9276
rect 27866 9220 27870 9276
rect 27806 9216 27870 9220
rect 27886 9276 27950 9280
rect 27886 9220 27890 9276
rect 27890 9220 27946 9276
rect 27946 9220 27950 9276
rect 27886 9216 27950 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 11438 8732 11502 8736
rect 11438 8676 11442 8732
rect 11442 8676 11498 8732
rect 11498 8676 11502 8732
rect 11438 8672 11502 8676
rect 11518 8732 11582 8736
rect 11518 8676 11522 8732
rect 11522 8676 11578 8732
rect 11578 8676 11582 8732
rect 11518 8672 11582 8676
rect 11598 8732 11662 8736
rect 11598 8676 11602 8732
rect 11602 8676 11658 8732
rect 11658 8676 11662 8732
rect 11598 8672 11662 8676
rect 11678 8732 11742 8736
rect 11678 8676 11682 8732
rect 11682 8676 11738 8732
rect 11738 8676 11742 8732
rect 11678 8672 11742 8676
rect 19212 8732 19276 8736
rect 19212 8676 19216 8732
rect 19216 8676 19272 8732
rect 19272 8676 19276 8732
rect 19212 8672 19276 8676
rect 19292 8732 19356 8736
rect 19292 8676 19296 8732
rect 19296 8676 19352 8732
rect 19352 8676 19356 8732
rect 19292 8672 19356 8676
rect 19372 8732 19436 8736
rect 19372 8676 19376 8732
rect 19376 8676 19432 8732
rect 19432 8676 19436 8732
rect 19372 8672 19436 8676
rect 19452 8732 19516 8736
rect 19452 8676 19456 8732
rect 19456 8676 19512 8732
rect 19512 8676 19516 8732
rect 19452 8672 19516 8676
rect 26986 8732 27050 8736
rect 26986 8676 26990 8732
rect 26990 8676 27046 8732
rect 27046 8676 27050 8732
rect 26986 8672 27050 8676
rect 27066 8732 27130 8736
rect 27066 8676 27070 8732
rect 27070 8676 27126 8732
rect 27126 8676 27130 8732
rect 27066 8672 27130 8676
rect 27146 8732 27210 8736
rect 27146 8676 27150 8732
rect 27150 8676 27206 8732
rect 27206 8676 27210 8732
rect 27146 8672 27210 8676
rect 27226 8732 27290 8736
rect 27226 8676 27230 8732
rect 27230 8676 27286 8732
rect 27286 8676 27290 8732
rect 27226 8672 27290 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 12098 8188 12162 8192
rect 12098 8132 12102 8188
rect 12102 8132 12158 8188
rect 12158 8132 12162 8188
rect 12098 8128 12162 8132
rect 12178 8188 12242 8192
rect 12178 8132 12182 8188
rect 12182 8132 12238 8188
rect 12238 8132 12242 8188
rect 12178 8128 12242 8132
rect 12258 8188 12322 8192
rect 12258 8132 12262 8188
rect 12262 8132 12318 8188
rect 12318 8132 12322 8188
rect 12258 8128 12322 8132
rect 12338 8188 12402 8192
rect 12338 8132 12342 8188
rect 12342 8132 12398 8188
rect 12398 8132 12402 8188
rect 12338 8128 12402 8132
rect 19872 8188 19936 8192
rect 19872 8132 19876 8188
rect 19876 8132 19932 8188
rect 19932 8132 19936 8188
rect 19872 8128 19936 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 27646 8188 27710 8192
rect 27646 8132 27650 8188
rect 27650 8132 27706 8188
rect 27706 8132 27710 8188
rect 27646 8128 27710 8132
rect 27726 8188 27790 8192
rect 27726 8132 27730 8188
rect 27730 8132 27786 8188
rect 27786 8132 27790 8188
rect 27726 8128 27790 8132
rect 27806 8188 27870 8192
rect 27806 8132 27810 8188
rect 27810 8132 27866 8188
rect 27866 8132 27870 8188
rect 27806 8128 27870 8132
rect 27886 8188 27950 8192
rect 27886 8132 27890 8188
rect 27890 8132 27946 8188
rect 27946 8132 27950 8188
rect 27886 8128 27950 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 11438 7644 11502 7648
rect 11438 7588 11442 7644
rect 11442 7588 11498 7644
rect 11498 7588 11502 7644
rect 11438 7584 11502 7588
rect 11518 7644 11582 7648
rect 11518 7588 11522 7644
rect 11522 7588 11578 7644
rect 11578 7588 11582 7644
rect 11518 7584 11582 7588
rect 11598 7644 11662 7648
rect 11598 7588 11602 7644
rect 11602 7588 11658 7644
rect 11658 7588 11662 7644
rect 11598 7584 11662 7588
rect 11678 7644 11742 7648
rect 11678 7588 11682 7644
rect 11682 7588 11738 7644
rect 11738 7588 11742 7644
rect 11678 7584 11742 7588
rect 19212 7644 19276 7648
rect 19212 7588 19216 7644
rect 19216 7588 19272 7644
rect 19272 7588 19276 7644
rect 19212 7584 19276 7588
rect 19292 7644 19356 7648
rect 19292 7588 19296 7644
rect 19296 7588 19352 7644
rect 19352 7588 19356 7644
rect 19292 7584 19356 7588
rect 19372 7644 19436 7648
rect 19372 7588 19376 7644
rect 19376 7588 19432 7644
rect 19432 7588 19436 7644
rect 19372 7584 19436 7588
rect 19452 7644 19516 7648
rect 19452 7588 19456 7644
rect 19456 7588 19512 7644
rect 19512 7588 19516 7644
rect 19452 7584 19516 7588
rect 26986 7644 27050 7648
rect 26986 7588 26990 7644
rect 26990 7588 27046 7644
rect 27046 7588 27050 7644
rect 26986 7584 27050 7588
rect 27066 7644 27130 7648
rect 27066 7588 27070 7644
rect 27070 7588 27126 7644
rect 27126 7588 27130 7644
rect 27066 7584 27130 7588
rect 27146 7644 27210 7648
rect 27146 7588 27150 7644
rect 27150 7588 27206 7644
rect 27206 7588 27210 7644
rect 27146 7584 27210 7588
rect 27226 7644 27290 7648
rect 27226 7588 27230 7644
rect 27230 7588 27286 7644
rect 27286 7588 27290 7644
rect 27226 7584 27290 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 12098 7100 12162 7104
rect 12098 7044 12102 7100
rect 12102 7044 12158 7100
rect 12158 7044 12162 7100
rect 12098 7040 12162 7044
rect 12178 7100 12242 7104
rect 12178 7044 12182 7100
rect 12182 7044 12238 7100
rect 12238 7044 12242 7100
rect 12178 7040 12242 7044
rect 12258 7100 12322 7104
rect 12258 7044 12262 7100
rect 12262 7044 12318 7100
rect 12318 7044 12322 7100
rect 12258 7040 12322 7044
rect 12338 7100 12402 7104
rect 12338 7044 12342 7100
rect 12342 7044 12398 7100
rect 12398 7044 12402 7100
rect 12338 7040 12402 7044
rect 19872 7100 19936 7104
rect 19872 7044 19876 7100
rect 19876 7044 19932 7100
rect 19932 7044 19936 7100
rect 19872 7040 19936 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 27646 7100 27710 7104
rect 27646 7044 27650 7100
rect 27650 7044 27706 7100
rect 27706 7044 27710 7100
rect 27646 7040 27710 7044
rect 27726 7100 27790 7104
rect 27726 7044 27730 7100
rect 27730 7044 27786 7100
rect 27786 7044 27790 7100
rect 27726 7040 27790 7044
rect 27806 7100 27870 7104
rect 27806 7044 27810 7100
rect 27810 7044 27866 7100
rect 27866 7044 27870 7100
rect 27806 7040 27870 7044
rect 27886 7100 27950 7104
rect 27886 7044 27890 7100
rect 27890 7044 27946 7100
rect 27946 7044 27950 7100
rect 27886 7040 27950 7044
rect 19012 6972 19076 7036
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 11438 6556 11502 6560
rect 11438 6500 11442 6556
rect 11442 6500 11498 6556
rect 11498 6500 11502 6556
rect 11438 6496 11502 6500
rect 11518 6556 11582 6560
rect 11518 6500 11522 6556
rect 11522 6500 11578 6556
rect 11578 6500 11582 6556
rect 11518 6496 11582 6500
rect 11598 6556 11662 6560
rect 11598 6500 11602 6556
rect 11602 6500 11658 6556
rect 11658 6500 11662 6556
rect 11598 6496 11662 6500
rect 11678 6556 11742 6560
rect 11678 6500 11682 6556
rect 11682 6500 11738 6556
rect 11738 6500 11742 6556
rect 11678 6496 11742 6500
rect 19212 6556 19276 6560
rect 19212 6500 19216 6556
rect 19216 6500 19272 6556
rect 19272 6500 19276 6556
rect 19212 6496 19276 6500
rect 19292 6556 19356 6560
rect 19292 6500 19296 6556
rect 19296 6500 19352 6556
rect 19352 6500 19356 6556
rect 19292 6496 19356 6500
rect 19372 6556 19436 6560
rect 19372 6500 19376 6556
rect 19376 6500 19432 6556
rect 19432 6500 19436 6556
rect 19372 6496 19436 6500
rect 19452 6556 19516 6560
rect 19452 6500 19456 6556
rect 19456 6500 19512 6556
rect 19512 6500 19516 6556
rect 19452 6496 19516 6500
rect 26986 6556 27050 6560
rect 26986 6500 26990 6556
rect 26990 6500 27046 6556
rect 27046 6500 27050 6556
rect 26986 6496 27050 6500
rect 27066 6556 27130 6560
rect 27066 6500 27070 6556
rect 27070 6500 27126 6556
rect 27126 6500 27130 6556
rect 27066 6496 27130 6500
rect 27146 6556 27210 6560
rect 27146 6500 27150 6556
rect 27150 6500 27206 6556
rect 27206 6500 27210 6556
rect 27146 6496 27210 6500
rect 27226 6556 27290 6560
rect 27226 6500 27230 6556
rect 27230 6500 27286 6556
rect 27286 6500 27290 6556
rect 27226 6496 27290 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 12098 6012 12162 6016
rect 12098 5956 12102 6012
rect 12102 5956 12158 6012
rect 12158 5956 12162 6012
rect 12098 5952 12162 5956
rect 12178 6012 12242 6016
rect 12178 5956 12182 6012
rect 12182 5956 12238 6012
rect 12238 5956 12242 6012
rect 12178 5952 12242 5956
rect 12258 6012 12322 6016
rect 12258 5956 12262 6012
rect 12262 5956 12318 6012
rect 12318 5956 12322 6012
rect 12258 5952 12322 5956
rect 12338 6012 12402 6016
rect 12338 5956 12342 6012
rect 12342 5956 12398 6012
rect 12398 5956 12402 6012
rect 12338 5952 12402 5956
rect 19872 6012 19936 6016
rect 19872 5956 19876 6012
rect 19876 5956 19932 6012
rect 19932 5956 19936 6012
rect 19872 5952 19936 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 27646 6012 27710 6016
rect 27646 5956 27650 6012
rect 27650 5956 27706 6012
rect 27706 5956 27710 6012
rect 27646 5952 27710 5956
rect 27726 6012 27790 6016
rect 27726 5956 27730 6012
rect 27730 5956 27786 6012
rect 27786 5956 27790 6012
rect 27726 5952 27790 5956
rect 27806 6012 27870 6016
rect 27806 5956 27810 6012
rect 27810 5956 27866 6012
rect 27866 5956 27870 6012
rect 27806 5952 27870 5956
rect 27886 6012 27950 6016
rect 27886 5956 27890 6012
rect 27890 5956 27946 6012
rect 27946 5956 27950 6012
rect 27886 5952 27950 5956
rect 19012 5944 19076 5948
rect 19012 5888 19062 5944
rect 19062 5888 19076 5944
rect 19012 5884 19076 5888
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 11438 5468 11502 5472
rect 11438 5412 11442 5468
rect 11442 5412 11498 5468
rect 11498 5412 11502 5468
rect 11438 5408 11502 5412
rect 11518 5468 11582 5472
rect 11518 5412 11522 5468
rect 11522 5412 11578 5468
rect 11578 5412 11582 5468
rect 11518 5408 11582 5412
rect 11598 5468 11662 5472
rect 11598 5412 11602 5468
rect 11602 5412 11658 5468
rect 11658 5412 11662 5468
rect 11598 5408 11662 5412
rect 11678 5468 11742 5472
rect 11678 5412 11682 5468
rect 11682 5412 11738 5468
rect 11738 5412 11742 5468
rect 11678 5408 11742 5412
rect 19212 5468 19276 5472
rect 19212 5412 19216 5468
rect 19216 5412 19272 5468
rect 19272 5412 19276 5468
rect 19212 5408 19276 5412
rect 19292 5468 19356 5472
rect 19292 5412 19296 5468
rect 19296 5412 19352 5468
rect 19352 5412 19356 5468
rect 19292 5408 19356 5412
rect 19372 5468 19436 5472
rect 19372 5412 19376 5468
rect 19376 5412 19432 5468
rect 19432 5412 19436 5468
rect 19372 5408 19436 5412
rect 19452 5468 19516 5472
rect 19452 5412 19456 5468
rect 19456 5412 19512 5468
rect 19512 5412 19516 5468
rect 19452 5408 19516 5412
rect 26986 5468 27050 5472
rect 26986 5412 26990 5468
rect 26990 5412 27046 5468
rect 27046 5412 27050 5468
rect 26986 5408 27050 5412
rect 27066 5468 27130 5472
rect 27066 5412 27070 5468
rect 27070 5412 27126 5468
rect 27126 5412 27130 5468
rect 27066 5408 27130 5412
rect 27146 5468 27210 5472
rect 27146 5412 27150 5468
rect 27150 5412 27206 5468
rect 27206 5412 27210 5468
rect 27146 5408 27210 5412
rect 27226 5468 27290 5472
rect 27226 5412 27230 5468
rect 27230 5412 27286 5468
rect 27286 5412 27290 5468
rect 27226 5408 27290 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 12098 4924 12162 4928
rect 12098 4868 12102 4924
rect 12102 4868 12158 4924
rect 12158 4868 12162 4924
rect 12098 4864 12162 4868
rect 12178 4924 12242 4928
rect 12178 4868 12182 4924
rect 12182 4868 12238 4924
rect 12238 4868 12242 4924
rect 12178 4864 12242 4868
rect 12258 4924 12322 4928
rect 12258 4868 12262 4924
rect 12262 4868 12318 4924
rect 12318 4868 12322 4924
rect 12258 4864 12322 4868
rect 12338 4924 12402 4928
rect 12338 4868 12342 4924
rect 12342 4868 12398 4924
rect 12398 4868 12402 4924
rect 12338 4864 12402 4868
rect 19872 4924 19936 4928
rect 19872 4868 19876 4924
rect 19876 4868 19932 4924
rect 19932 4868 19936 4924
rect 19872 4864 19936 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 27646 4924 27710 4928
rect 27646 4868 27650 4924
rect 27650 4868 27706 4924
rect 27706 4868 27710 4924
rect 27646 4864 27710 4868
rect 27726 4924 27790 4928
rect 27726 4868 27730 4924
rect 27730 4868 27786 4924
rect 27786 4868 27790 4924
rect 27726 4864 27790 4868
rect 27806 4924 27870 4928
rect 27806 4868 27810 4924
rect 27810 4868 27866 4924
rect 27866 4868 27870 4924
rect 27806 4864 27870 4868
rect 27886 4924 27950 4928
rect 27886 4868 27890 4924
rect 27890 4868 27946 4924
rect 27946 4868 27950 4924
rect 27886 4864 27950 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 11438 4380 11502 4384
rect 11438 4324 11442 4380
rect 11442 4324 11498 4380
rect 11498 4324 11502 4380
rect 11438 4320 11502 4324
rect 11518 4380 11582 4384
rect 11518 4324 11522 4380
rect 11522 4324 11578 4380
rect 11578 4324 11582 4380
rect 11518 4320 11582 4324
rect 11598 4380 11662 4384
rect 11598 4324 11602 4380
rect 11602 4324 11658 4380
rect 11658 4324 11662 4380
rect 11598 4320 11662 4324
rect 11678 4380 11742 4384
rect 11678 4324 11682 4380
rect 11682 4324 11738 4380
rect 11738 4324 11742 4380
rect 11678 4320 11742 4324
rect 19212 4380 19276 4384
rect 19212 4324 19216 4380
rect 19216 4324 19272 4380
rect 19272 4324 19276 4380
rect 19212 4320 19276 4324
rect 19292 4380 19356 4384
rect 19292 4324 19296 4380
rect 19296 4324 19352 4380
rect 19352 4324 19356 4380
rect 19292 4320 19356 4324
rect 19372 4380 19436 4384
rect 19372 4324 19376 4380
rect 19376 4324 19432 4380
rect 19432 4324 19436 4380
rect 19372 4320 19436 4324
rect 19452 4380 19516 4384
rect 19452 4324 19456 4380
rect 19456 4324 19512 4380
rect 19512 4324 19516 4380
rect 19452 4320 19516 4324
rect 26986 4380 27050 4384
rect 26986 4324 26990 4380
rect 26990 4324 27046 4380
rect 27046 4324 27050 4380
rect 26986 4320 27050 4324
rect 27066 4380 27130 4384
rect 27066 4324 27070 4380
rect 27070 4324 27126 4380
rect 27126 4324 27130 4380
rect 27066 4320 27130 4324
rect 27146 4380 27210 4384
rect 27146 4324 27150 4380
rect 27150 4324 27206 4380
rect 27206 4324 27210 4380
rect 27146 4320 27210 4324
rect 27226 4380 27290 4384
rect 27226 4324 27230 4380
rect 27230 4324 27286 4380
rect 27286 4324 27290 4380
rect 27226 4320 27290 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 12098 3836 12162 3840
rect 12098 3780 12102 3836
rect 12102 3780 12158 3836
rect 12158 3780 12162 3836
rect 12098 3776 12162 3780
rect 12178 3836 12242 3840
rect 12178 3780 12182 3836
rect 12182 3780 12238 3836
rect 12238 3780 12242 3836
rect 12178 3776 12242 3780
rect 12258 3836 12322 3840
rect 12258 3780 12262 3836
rect 12262 3780 12318 3836
rect 12318 3780 12322 3836
rect 12258 3776 12322 3780
rect 12338 3836 12402 3840
rect 12338 3780 12342 3836
rect 12342 3780 12398 3836
rect 12398 3780 12402 3836
rect 12338 3776 12402 3780
rect 19872 3836 19936 3840
rect 19872 3780 19876 3836
rect 19876 3780 19932 3836
rect 19932 3780 19936 3836
rect 19872 3776 19936 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 27646 3836 27710 3840
rect 27646 3780 27650 3836
rect 27650 3780 27706 3836
rect 27706 3780 27710 3836
rect 27646 3776 27710 3780
rect 27726 3836 27790 3840
rect 27726 3780 27730 3836
rect 27730 3780 27786 3836
rect 27786 3780 27790 3836
rect 27726 3776 27790 3780
rect 27806 3836 27870 3840
rect 27806 3780 27810 3836
rect 27810 3780 27866 3836
rect 27866 3780 27870 3836
rect 27806 3776 27870 3780
rect 27886 3836 27950 3840
rect 27886 3780 27890 3836
rect 27890 3780 27946 3836
rect 27946 3780 27950 3836
rect 27886 3776 27950 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 11438 3292 11502 3296
rect 11438 3236 11442 3292
rect 11442 3236 11498 3292
rect 11498 3236 11502 3292
rect 11438 3232 11502 3236
rect 11518 3292 11582 3296
rect 11518 3236 11522 3292
rect 11522 3236 11578 3292
rect 11578 3236 11582 3292
rect 11518 3232 11582 3236
rect 11598 3292 11662 3296
rect 11598 3236 11602 3292
rect 11602 3236 11658 3292
rect 11658 3236 11662 3292
rect 11598 3232 11662 3236
rect 11678 3292 11742 3296
rect 11678 3236 11682 3292
rect 11682 3236 11738 3292
rect 11738 3236 11742 3292
rect 11678 3232 11742 3236
rect 19212 3292 19276 3296
rect 19212 3236 19216 3292
rect 19216 3236 19272 3292
rect 19272 3236 19276 3292
rect 19212 3232 19276 3236
rect 19292 3292 19356 3296
rect 19292 3236 19296 3292
rect 19296 3236 19352 3292
rect 19352 3236 19356 3292
rect 19292 3232 19356 3236
rect 19372 3292 19436 3296
rect 19372 3236 19376 3292
rect 19376 3236 19432 3292
rect 19432 3236 19436 3292
rect 19372 3232 19436 3236
rect 19452 3292 19516 3296
rect 19452 3236 19456 3292
rect 19456 3236 19512 3292
rect 19512 3236 19516 3292
rect 19452 3232 19516 3236
rect 26986 3292 27050 3296
rect 26986 3236 26990 3292
rect 26990 3236 27046 3292
rect 27046 3236 27050 3292
rect 26986 3232 27050 3236
rect 27066 3292 27130 3296
rect 27066 3236 27070 3292
rect 27070 3236 27126 3292
rect 27126 3236 27130 3292
rect 27066 3232 27130 3236
rect 27146 3292 27210 3296
rect 27146 3236 27150 3292
rect 27150 3236 27206 3292
rect 27206 3236 27210 3292
rect 27146 3232 27210 3236
rect 27226 3292 27290 3296
rect 27226 3236 27230 3292
rect 27230 3236 27286 3292
rect 27286 3236 27290 3292
rect 27226 3232 27290 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 12098 2748 12162 2752
rect 12098 2692 12102 2748
rect 12102 2692 12158 2748
rect 12158 2692 12162 2748
rect 12098 2688 12162 2692
rect 12178 2748 12242 2752
rect 12178 2692 12182 2748
rect 12182 2692 12238 2748
rect 12238 2692 12242 2748
rect 12178 2688 12242 2692
rect 12258 2748 12322 2752
rect 12258 2692 12262 2748
rect 12262 2692 12318 2748
rect 12318 2692 12322 2748
rect 12258 2688 12322 2692
rect 12338 2748 12402 2752
rect 12338 2692 12342 2748
rect 12342 2692 12398 2748
rect 12398 2692 12402 2748
rect 12338 2688 12402 2692
rect 19872 2748 19936 2752
rect 19872 2692 19876 2748
rect 19876 2692 19932 2748
rect 19932 2692 19936 2748
rect 19872 2688 19936 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 27646 2748 27710 2752
rect 27646 2692 27650 2748
rect 27650 2692 27706 2748
rect 27706 2692 27710 2748
rect 27646 2688 27710 2692
rect 27726 2748 27790 2752
rect 27726 2692 27730 2748
rect 27730 2692 27786 2748
rect 27786 2692 27790 2748
rect 27726 2688 27790 2692
rect 27806 2748 27870 2752
rect 27806 2692 27810 2748
rect 27810 2692 27866 2748
rect 27866 2692 27870 2748
rect 27806 2688 27870 2692
rect 27886 2748 27950 2752
rect 27886 2692 27890 2748
rect 27890 2692 27946 2748
rect 27946 2692 27950 2748
rect 27886 2688 27950 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 11438 2204 11502 2208
rect 11438 2148 11442 2204
rect 11442 2148 11498 2204
rect 11498 2148 11502 2204
rect 11438 2144 11502 2148
rect 11518 2204 11582 2208
rect 11518 2148 11522 2204
rect 11522 2148 11578 2204
rect 11578 2148 11582 2204
rect 11518 2144 11582 2148
rect 11598 2204 11662 2208
rect 11598 2148 11602 2204
rect 11602 2148 11658 2204
rect 11658 2148 11662 2204
rect 11598 2144 11662 2148
rect 11678 2204 11742 2208
rect 11678 2148 11682 2204
rect 11682 2148 11738 2204
rect 11738 2148 11742 2204
rect 11678 2144 11742 2148
rect 19212 2204 19276 2208
rect 19212 2148 19216 2204
rect 19216 2148 19272 2204
rect 19272 2148 19276 2204
rect 19212 2144 19276 2148
rect 19292 2204 19356 2208
rect 19292 2148 19296 2204
rect 19296 2148 19352 2204
rect 19352 2148 19356 2204
rect 19292 2144 19356 2148
rect 19372 2204 19436 2208
rect 19372 2148 19376 2204
rect 19376 2148 19432 2204
rect 19432 2148 19436 2204
rect 19372 2144 19436 2148
rect 19452 2204 19516 2208
rect 19452 2148 19456 2204
rect 19456 2148 19512 2204
rect 19512 2148 19516 2204
rect 19452 2144 19516 2148
rect 26986 2204 27050 2208
rect 26986 2148 26990 2204
rect 26990 2148 27046 2204
rect 27046 2148 27050 2204
rect 26986 2144 27050 2148
rect 27066 2204 27130 2208
rect 27066 2148 27070 2204
rect 27070 2148 27126 2204
rect 27126 2148 27130 2204
rect 27066 2144 27130 2148
rect 27146 2204 27210 2208
rect 27146 2148 27150 2204
rect 27150 2148 27206 2204
rect 27206 2148 27210 2204
rect 27146 2144 27210 2148
rect 27226 2204 27290 2208
rect 27226 2148 27230 2204
rect 27230 2148 27286 2204
rect 27286 2148 27290 2204
rect 27226 2144 27290 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 12098 1660 12162 1664
rect 12098 1604 12102 1660
rect 12102 1604 12158 1660
rect 12158 1604 12162 1660
rect 12098 1600 12162 1604
rect 12178 1660 12242 1664
rect 12178 1604 12182 1660
rect 12182 1604 12238 1660
rect 12238 1604 12242 1660
rect 12178 1600 12242 1604
rect 12258 1660 12322 1664
rect 12258 1604 12262 1660
rect 12262 1604 12318 1660
rect 12318 1604 12322 1660
rect 12258 1600 12322 1604
rect 12338 1660 12402 1664
rect 12338 1604 12342 1660
rect 12342 1604 12398 1660
rect 12398 1604 12402 1660
rect 12338 1600 12402 1604
rect 19872 1660 19936 1664
rect 19872 1604 19876 1660
rect 19876 1604 19932 1660
rect 19932 1604 19936 1660
rect 19872 1600 19936 1604
rect 19952 1660 20016 1664
rect 19952 1604 19956 1660
rect 19956 1604 20012 1660
rect 20012 1604 20016 1660
rect 19952 1600 20016 1604
rect 20032 1660 20096 1664
rect 20032 1604 20036 1660
rect 20036 1604 20092 1660
rect 20092 1604 20096 1660
rect 20032 1600 20096 1604
rect 20112 1660 20176 1664
rect 20112 1604 20116 1660
rect 20116 1604 20172 1660
rect 20172 1604 20176 1660
rect 20112 1600 20176 1604
rect 27646 1660 27710 1664
rect 27646 1604 27650 1660
rect 27650 1604 27706 1660
rect 27706 1604 27710 1660
rect 27646 1600 27710 1604
rect 27726 1660 27790 1664
rect 27726 1604 27730 1660
rect 27730 1604 27786 1660
rect 27786 1604 27790 1660
rect 27726 1600 27790 1604
rect 27806 1660 27870 1664
rect 27806 1604 27810 1660
rect 27810 1604 27866 1660
rect 27866 1604 27870 1660
rect 27806 1600 27870 1604
rect 27886 1660 27950 1664
rect 27886 1604 27890 1660
rect 27890 1604 27946 1660
rect 27946 1604 27950 1660
rect 27886 1600 27950 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 11438 1116 11502 1120
rect 11438 1060 11442 1116
rect 11442 1060 11498 1116
rect 11498 1060 11502 1116
rect 11438 1056 11502 1060
rect 11518 1116 11582 1120
rect 11518 1060 11522 1116
rect 11522 1060 11578 1116
rect 11578 1060 11582 1116
rect 11518 1056 11582 1060
rect 11598 1116 11662 1120
rect 11598 1060 11602 1116
rect 11602 1060 11658 1116
rect 11658 1060 11662 1116
rect 11598 1056 11662 1060
rect 11678 1116 11742 1120
rect 11678 1060 11682 1116
rect 11682 1060 11738 1116
rect 11738 1060 11742 1116
rect 11678 1056 11742 1060
rect 19212 1116 19276 1120
rect 19212 1060 19216 1116
rect 19216 1060 19272 1116
rect 19272 1060 19276 1116
rect 19212 1056 19276 1060
rect 19292 1116 19356 1120
rect 19292 1060 19296 1116
rect 19296 1060 19352 1116
rect 19352 1060 19356 1116
rect 19292 1056 19356 1060
rect 19372 1116 19436 1120
rect 19372 1060 19376 1116
rect 19376 1060 19432 1116
rect 19432 1060 19436 1116
rect 19372 1056 19436 1060
rect 19452 1116 19516 1120
rect 19452 1060 19456 1116
rect 19456 1060 19512 1116
rect 19512 1060 19516 1116
rect 19452 1056 19516 1060
rect 26986 1116 27050 1120
rect 26986 1060 26990 1116
rect 26990 1060 27046 1116
rect 27046 1060 27050 1116
rect 26986 1056 27050 1060
rect 27066 1116 27130 1120
rect 27066 1060 27070 1116
rect 27070 1060 27126 1116
rect 27126 1060 27130 1116
rect 27066 1056 27130 1060
rect 27146 1116 27210 1120
rect 27146 1060 27150 1116
rect 27150 1060 27206 1116
rect 27206 1060 27210 1116
rect 27146 1056 27210 1060
rect 27226 1116 27290 1120
rect 27226 1060 27230 1116
rect 27230 1060 27286 1116
rect 27286 1060 27290 1116
rect 27226 1056 27290 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 12098 572 12162 576
rect 12098 516 12102 572
rect 12102 516 12158 572
rect 12158 516 12162 572
rect 12098 512 12162 516
rect 12178 572 12242 576
rect 12178 516 12182 572
rect 12182 516 12238 572
rect 12238 516 12242 572
rect 12178 512 12242 516
rect 12258 572 12322 576
rect 12258 516 12262 572
rect 12262 516 12318 572
rect 12318 516 12322 572
rect 12258 512 12322 516
rect 12338 572 12402 576
rect 12338 516 12342 572
rect 12342 516 12398 572
rect 12398 516 12402 572
rect 12338 512 12402 516
rect 19872 572 19936 576
rect 19872 516 19876 572
rect 19876 516 19932 572
rect 19932 516 19936 572
rect 19872 512 19936 516
rect 19952 572 20016 576
rect 19952 516 19956 572
rect 19956 516 20012 572
rect 20012 516 20016 572
rect 19952 512 20016 516
rect 20032 572 20096 576
rect 20032 516 20036 572
rect 20036 516 20092 572
rect 20092 516 20096 572
rect 20032 512 20096 516
rect 20112 572 20176 576
rect 20112 516 20116 572
rect 20116 516 20172 572
rect 20172 516 20176 572
rect 20112 512 20176 516
rect 27646 572 27710 576
rect 27646 516 27650 572
rect 27650 516 27706 572
rect 27706 516 27710 572
rect 27646 512 27710 516
rect 27726 572 27790 576
rect 27726 516 27730 572
rect 27730 516 27786 572
rect 27786 516 27790 572
rect 27726 512 27790 516
rect 27806 572 27870 576
rect 27806 516 27810 572
rect 27810 516 27866 572
rect 27866 516 27870 572
rect 27806 512 27870 516
rect 27886 572 27950 576
rect 27886 516 27890 572
rect 27890 516 27946 572
rect 27946 516 27950 572
rect 27886 512 27950 516
<< metal4 >>
rect 3656 21792 3976 21808
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 21248 4636 21808
rect 6134 21725 6194 22304
rect 6131 21724 6197 21725
rect 6131 21660 6132 21724
rect 6196 21660 6197 21724
rect 6131 21659 6197 21660
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 6686 20365 6746 22304
rect 7238 21861 7298 22304
rect 7235 21860 7301 21861
rect 7235 21796 7236 21860
rect 7300 21796 7301 21860
rect 7235 21795 7301 21796
rect 7790 21725 7850 22304
rect 8342 21725 8402 22304
rect 7787 21724 7853 21725
rect 7787 21660 7788 21724
rect 7852 21660 7853 21724
rect 7787 21659 7853 21660
rect 8339 21724 8405 21725
rect 8339 21660 8340 21724
rect 8404 21660 8405 21724
rect 8339 21659 8405 21660
rect 8894 21181 8954 22304
rect 9446 21317 9506 22304
rect 9443 21316 9509 21317
rect 9443 21252 9444 21316
rect 9508 21252 9509 21316
rect 9443 21251 9509 21252
rect 9998 21181 10058 22304
rect 8891 21180 8957 21181
rect 8891 21116 8892 21180
rect 8956 21116 8957 21180
rect 8891 21115 8957 21116
rect 9995 21180 10061 21181
rect 9995 21116 9996 21180
rect 10060 21116 10061 21180
rect 9995 21115 10061 21116
rect 6683 20364 6749 20365
rect 6683 20300 6684 20364
rect 6748 20300 6749 20364
rect 6683 20299 6749 20300
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 10550 12341 10610 22304
rect 11102 20637 11162 22304
rect 11654 21997 11714 22304
rect 12206 21997 12266 22304
rect 11651 21996 11717 21997
rect 11651 21932 11652 21996
rect 11716 21932 11717 21996
rect 11651 21931 11717 21932
rect 12203 21996 12269 21997
rect 12203 21932 12204 21996
rect 12268 21932 12269 21996
rect 12203 21931 12269 21932
rect 11430 21792 11750 21808
rect 11430 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11750 21792
rect 11430 20704 11750 21728
rect 11430 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11750 20704
rect 11099 20636 11165 20637
rect 11099 20572 11100 20636
rect 11164 20572 11165 20636
rect 11099 20571 11165 20572
rect 11430 19616 11750 20640
rect 11430 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11750 19616
rect 11430 18528 11750 19552
rect 11430 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11750 18528
rect 11430 17440 11750 18464
rect 11430 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11750 17440
rect 11430 16352 11750 17376
rect 11430 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11750 16352
rect 11430 15264 11750 16288
rect 11430 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11750 15264
rect 11430 14176 11750 15200
rect 11430 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11750 14176
rect 11430 13088 11750 14112
rect 11430 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11750 13088
rect 10547 12340 10613 12341
rect 10547 12276 10548 12340
rect 10612 12276 10613 12340
rect 10547 12275 10613 12276
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 11430 12000 11750 13024
rect 11430 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11750 12000
rect 11430 10912 11750 11936
rect 11430 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11750 10912
rect 11430 9824 11750 10848
rect 11430 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11750 9824
rect 11430 8736 11750 9760
rect 11430 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11750 8736
rect 11430 7648 11750 8672
rect 11430 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11750 7648
rect 11430 6560 11750 7584
rect 11430 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11750 6560
rect 11430 5472 11750 6496
rect 11430 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11750 5472
rect 11430 4384 11750 5408
rect 11430 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11750 4384
rect 11430 3296 11750 4320
rect 11430 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11750 3296
rect 11430 2208 11750 3232
rect 11430 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11750 2208
rect 11430 1120 11750 2144
rect 11430 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11750 1120
rect 11430 496 11750 1056
rect 12090 21248 12410 21808
rect 12758 21725 12818 22304
rect 12755 21724 12821 21725
rect 12755 21660 12756 21724
rect 12820 21660 12821 21724
rect 12755 21659 12821 21660
rect 12090 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12410 21248
rect 12090 20160 12410 21184
rect 13310 20637 13370 22304
rect 13307 20636 13373 20637
rect 13307 20572 13308 20636
rect 13372 20572 13373 20636
rect 13307 20571 13373 20572
rect 12090 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12410 20160
rect 12090 19072 12410 20096
rect 12090 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12410 19072
rect 12090 17984 12410 19008
rect 13862 18869 13922 22304
rect 14414 19277 14474 22304
rect 14966 20637 15026 22304
rect 15518 20773 15578 22304
rect 16070 20909 16130 22304
rect 16067 20908 16133 20909
rect 16067 20844 16068 20908
rect 16132 20844 16133 20908
rect 16067 20843 16133 20844
rect 15515 20772 15581 20773
rect 15515 20708 15516 20772
rect 15580 20708 15581 20772
rect 15515 20707 15581 20708
rect 16622 20637 16682 22304
rect 17174 21453 17234 22304
rect 17171 21452 17237 21453
rect 17171 21388 17172 21452
rect 17236 21388 17237 21452
rect 17171 21387 17237 21388
rect 14963 20636 15029 20637
rect 14963 20572 14964 20636
rect 15028 20572 15029 20636
rect 14963 20571 15029 20572
rect 16619 20636 16685 20637
rect 16619 20572 16620 20636
rect 16684 20572 16685 20636
rect 16619 20571 16685 20572
rect 17726 19957 17786 22304
rect 18278 21181 18338 22304
rect 18275 21180 18341 21181
rect 18275 21116 18276 21180
rect 18340 21116 18341 21180
rect 18275 21115 18341 21116
rect 18830 21045 18890 22304
rect 19382 22104 19442 22304
rect 19934 22104 19994 22304
rect 20486 22104 20546 22304
rect 21038 22104 21098 22304
rect 21590 21861 21650 22304
rect 22142 22104 22202 22304
rect 22694 22104 22754 22304
rect 23246 22104 23306 22304
rect 23798 21861 23858 22304
rect 24350 21997 24410 22304
rect 24347 21996 24413 21997
rect 24347 21932 24348 21996
rect 24412 21932 24413 21996
rect 24347 21931 24413 21932
rect 21587 21860 21653 21861
rect 19204 21792 19524 21808
rect 19204 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19524 21792
rect 18827 21044 18893 21045
rect 18827 20980 18828 21044
rect 18892 20980 18893 21044
rect 18827 20979 18893 20980
rect 19204 20704 19524 21728
rect 19204 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19524 20704
rect 17723 19956 17789 19957
rect 17723 19892 17724 19956
rect 17788 19892 17789 19956
rect 17723 19891 17789 19892
rect 19204 19616 19524 20640
rect 19204 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19524 19616
rect 14411 19276 14477 19277
rect 14411 19212 14412 19276
rect 14476 19212 14477 19276
rect 14411 19211 14477 19212
rect 13859 18868 13925 18869
rect 13859 18804 13860 18868
rect 13924 18804 13925 18868
rect 13859 18803 13925 18804
rect 12090 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12410 17984
rect 12090 16896 12410 17920
rect 12090 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12410 16896
rect 12090 15808 12410 16832
rect 12090 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12410 15808
rect 12090 14720 12410 15744
rect 12090 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12410 14720
rect 12090 13632 12410 14656
rect 12090 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12410 13632
rect 12090 12544 12410 13568
rect 12090 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12410 12544
rect 12090 11456 12410 12480
rect 12090 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12410 11456
rect 12090 10368 12410 11392
rect 12090 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12410 10368
rect 12090 9280 12410 10304
rect 12090 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12410 9280
rect 12090 8192 12410 9216
rect 12090 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12410 8192
rect 12090 7104 12410 8128
rect 12090 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12410 7104
rect 12090 6016 12410 7040
rect 19204 18528 19524 19552
rect 19204 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19524 18528
rect 19204 17440 19524 18464
rect 19204 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19524 17440
rect 19204 16352 19524 17376
rect 19204 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19524 16352
rect 19204 15264 19524 16288
rect 19204 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19524 15264
rect 19204 14176 19524 15200
rect 19204 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19524 14176
rect 19204 13088 19524 14112
rect 19204 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19524 13088
rect 19204 12000 19524 13024
rect 19204 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19524 12000
rect 19204 10912 19524 11936
rect 19204 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19524 10912
rect 19204 9824 19524 10848
rect 19204 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19524 9824
rect 19204 8736 19524 9760
rect 19204 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19524 8736
rect 19204 7648 19524 8672
rect 19204 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19524 7648
rect 19011 7036 19077 7037
rect 19011 6972 19012 7036
rect 19076 6972 19077 7036
rect 19011 6971 19077 6972
rect 12090 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12410 6016
rect 12090 4928 12410 5952
rect 19014 5949 19074 6971
rect 19204 6560 19524 7584
rect 19204 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19524 6560
rect 19011 5948 19077 5949
rect 19011 5884 19012 5948
rect 19076 5884 19077 5948
rect 19011 5883 19077 5884
rect 12090 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12410 4928
rect 12090 3840 12410 4864
rect 12090 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12410 3840
rect 12090 2752 12410 3776
rect 12090 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12410 2752
rect 12090 1664 12410 2688
rect 12090 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12410 1664
rect 12090 576 12410 1600
rect 12090 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12410 576
rect 12090 496 12410 512
rect 19204 5472 19524 6496
rect 19204 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19524 5472
rect 19204 4384 19524 5408
rect 19204 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19524 4384
rect 19204 3296 19524 4320
rect 19204 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19524 3296
rect 19204 2208 19524 3232
rect 19204 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19524 2208
rect 19204 1120 19524 2144
rect 19204 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19524 1120
rect 19204 496 19524 1056
rect 19864 21248 20184 21808
rect 21587 21796 21588 21860
rect 21652 21796 21653 21860
rect 21587 21795 21653 21796
rect 23795 21860 23861 21861
rect 23795 21796 23796 21860
rect 23860 21796 23861 21860
rect 23795 21795 23861 21796
rect 24902 21725 24962 22304
rect 24899 21724 24965 21725
rect 24899 21660 24900 21724
rect 24964 21660 24965 21724
rect 24899 21659 24965 21660
rect 25454 21589 25514 22304
rect 26006 21861 26066 22304
rect 26558 21861 26618 22304
rect 27110 21997 27170 22304
rect 27662 21997 27722 22304
rect 27107 21996 27173 21997
rect 27107 21932 27108 21996
rect 27172 21932 27173 21996
rect 27107 21931 27173 21932
rect 27659 21996 27725 21997
rect 27659 21932 27660 21996
rect 27724 21932 27725 21996
rect 27659 21931 27725 21932
rect 28214 21861 28274 22304
rect 26003 21860 26069 21861
rect 26003 21796 26004 21860
rect 26068 21796 26069 21860
rect 26003 21795 26069 21796
rect 26555 21860 26621 21861
rect 26555 21796 26556 21860
rect 26620 21796 26621 21860
rect 28211 21860 28277 21861
rect 26555 21795 26621 21796
rect 26978 21792 27298 21808
rect 26978 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27298 21792
rect 25451 21588 25517 21589
rect 25451 21524 25452 21588
rect 25516 21524 25517 21588
rect 25451 21523 25517 21524
rect 19864 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20184 21248
rect 19864 20160 20184 21184
rect 19864 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20184 20160
rect 19864 19072 20184 20096
rect 19864 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20184 19072
rect 19864 17984 20184 19008
rect 26978 20704 27298 21728
rect 26978 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27298 20704
rect 26978 19616 27298 20640
rect 26978 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27298 19616
rect 26978 18528 27298 19552
rect 26978 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27298 18528
rect 20299 18188 20365 18189
rect 20299 18124 20300 18188
rect 20364 18124 20365 18188
rect 20299 18123 20365 18124
rect 19864 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20184 17984
rect 19864 16896 20184 17920
rect 19864 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20184 16896
rect 19864 15808 20184 16832
rect 19864 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20184 15808
rect 19864 14720 20184 15744
rect 19864 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20184 14720
rect 19864 13632 20184 14656
rect 19864 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20184 13632
rect 19864 12544 20184 13568
rect 19864 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20184 12544
rect 19864 11456 20184 12480
rect 19864 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20184 11456
rect 19864 10368 20184 11392
rect 20302 11253 20362 18123
rect 26978 17440 27298 18464
rect 26978 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27298 17440
rect 26978 16352 27298 17376
rect 26978 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27298 16352
rect 26978 15264 27298 16288
rect 26978 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27298 15264
rect 26978 14176 27298 15200
rect 26978 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27298 14176
rect 26978 13088 27298 14112
rect 26978 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27298 13088
rect 26978 12000 27298 13024
rect 26978 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27298 12000
rect 20299 11252 20365 11253
rect 20299 11188 20300 11252
rect 20364 11188 20365 11252
rect 20299 11187 20365 11188
rect 19864 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20184 10368
rect 19864 9280 20184 10304
rect 19864 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20184 9280
rect 19864 8192 20184 9216
rect 19864 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20184 8192
rect 19864 7104 20184 8128
rect 19864 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20184 7104
rect 19864 6016 20184 7040
rect 19864 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20184 6016
rect 19864 4928 20184 5952
rect 19864 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20184 4928
rect 19864 3840 20184 4864
rect 19864 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20184 3840
rect 19864 2752 20184 3776
rect 19864 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20184 2752
rect 19864 1664 20184 2688
rect 19864 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20184 1664
rect 19864 576 20184 1600
rect 19864 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20184 576
rect 19864 496 20184 512
rect 26978 10912 27298 11936
rect 26978 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27298 10912
rect 26978 9824 27298 10848
rect 26978 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27298 9824
rect 26978 8736 27298 9760
rect 26978 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27298 8736
rect 26978 7648 27298 8672
rect 26978 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27298 7648
rect 26978 6560 27298 7584
rect 26978 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27298 6560
rect 26978 5472 27298 6496
rect 26978 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27298 5472
rect 26978 4384 27298 5408
rect 26978 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27298 4384
rect 26978 3296 27298 4320
rect 26978 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27298 3296
rect 26978 2208 27298 3232
rect 26978 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27298 2208
rect 26978 1120 27298 2144
rect 26978 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27298 1120
rect 26978 496 27298 1056
rect 27638 21248 27958 21808
rect 28211 21796 28212 21860
rect 28276 21796 28277 21860
rect 28211 21795 28277 21796
rect 27638 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27958 21248
rect 27638 20160 27958 21184
rect 27638 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27958 20160
rect 27638 19072 27958 20096
rect 27638 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27958 19072
rect 27638 17984 27958 19008
rect 27638 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27958 17984
rect 27638 16896 27958 17920
rect 27638 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27958 16896
rect 27638 15808 27958 16832
rect 27638 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27958 15808
rect 27638 14720 27958 15744
rect 27638 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27958 14720
rect 27638 13632 27958 14656
rect 27638 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27958 13632
rect 27638 12544 27958 13568
rect 27638 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27958 12544
rect 27638 11456 27958 12480
rect 28766 11661 28826 22304
rect 29318 22104 29378 22304
rect 28763 11660 28829 11661
rect 28763 11596 28764 11660
rect 28828 11596 28829 11660
rect 28763 11595 28829 11596
rect 27638 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27958 11456
rect 27638 10368 27958 11392
rect 27638 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27958 10368
rect 27638 9280 27958 10304
rect 27638 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27958 9280
rect 27638 8192 27958 9216
rect 27638 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27958 8192
rect 27638 7104 27958 8128
rect 27638 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27958 7104
rect 27638 6016 27958 7040
rect 27638 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27958 6016
rect 27638 4928 27958 5952
rect 27638 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27958 4928
rect 27638 3840 27958 4864
rect 27638 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27958 3840
rect 27638 2752 27958 3776
rect 27638 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27958 2752
rect 27638 1664 27958 2688
rect 27638 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27958 1664
rect 27638 576 27958 1600
rect 27638 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27958 576
rect 27638 496 27958 512
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1
transform -1 0 6716 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1
transform 1 0 18676 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1
transform 1 0 18676 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1
transform -1 0 21988 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1
transform 1 0 22172 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1
transform -1 0 18676 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1
transform -1 0 24104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1
transform -1 0 24104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1
transform -1 0 25576 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1
transform 1 0 24196 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1
transform -1 0 26496 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1
transform -1 0 29900 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1
transform -1 0 5612 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1
transform 1 0 6072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1
transform 1 0 5060 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1
transform -1 0 3496 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1
transform 1 0 4416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1
transform 1 0 10672 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1
transform 1 0 29900 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1
transform -1 0 20148 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1
transform 1 0 12144 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1
transform 1 0 21988 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1
transform -1 0 27048 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1
transform -1 0 25208 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781__1
timestamp 1
transform 1 0 5336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781__2
timestamp 1
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0782_
timestamp 1
transform -1 0 8004 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _0783_
timestamp 1
transform 1 0 6808 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _0784_
timestamp 1
transform -1 0 13800 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__mux4_1  _0785_
timestamp 1
transform 1 0 4876 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0786_
timestamp 1
transform 1 0 4968 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _0787_
timestamp 1
transform -1 0 8280 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0788_
timestamp 1
transform -1 0 8924 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0789_
timestamp 1
transform -1 0 11224 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0790_
timestamp 1
transform 1 0 7268 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1
transform 1 0 9200 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_2  _0792_
timestamp 1
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0793_
timestamp 1
transform 1 0 25760 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0794_
timestamp 1
transform -1 0 26220 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0795_
timestamp 1
transform 1 0 20976 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0796_
timestamp 1
transform 1 0 22908 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0797_
timestamp 1
transform 1 0 26220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0798_
timestamp 1
transform -1 0 26128 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0799_
timestamp 1
transform 1 0 15916 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0800_
timestamp 1
transform 1 0 20148 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0801_
timestamp 1
transform -1 0 25668 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0802_
timestamp 1
transform 1 0 23920 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0803_
timestamp 1
transform 1 0 26956 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0804_
timestamp 1
transform 1 0 21528 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0805_
timestamp 1
transform 1 0 22080 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0806_
timestamp 1
transform -1 0 23460 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0807_
timestamp 1
transform 1 0 24380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0808_
timestamp 1
transform -1 0 26956 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0809_
timestamp 1
transform -1 0 26956 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0810_
timestamp 1
transform 1 0 19412 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0811_
timestamp 1
transform 1 0 22632 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0812_
timestamp 1
transform -1 0 23276 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0813_
timestamp 1
transform -1 0 25116 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0814_
timestamp 1
transform 1 0 16928 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0815_
timestamp 1
transform 1 0 18676 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _0816_
timestamp 1
transform 1 0 23552 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 1
transform -1 0 19780 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0818_
timestamp 1
transform 1 0 23276 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0819_
timestamp 1
transform -1 0 22908 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0820_
timestamp 1
transform -1 0 27140 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0821_
timestamp 1
transform 1 0 22540 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0822_
timestamp 1
transform 1 0 21804 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0823_
timestamp 1
transform -1 0 24748 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0824_
timestamp 1
transform -1 0 23920 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0825_
timestamp 1
transform -1 0 23736 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0826_
timestamp 1
transform -1 0 17388 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0827_
timestamp 1
transform -1 0 18400 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0828_
timestamp 1
transform -1 0 24656 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0829_
timestamp 1
transform -1 0 25576 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0830_
timestamp 1
transform -1 0 24380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1
transform -1 0 22448 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0832_
timestamp 1
transform -1 0 21896 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0833_
timestamp 1
transform 1 0 22448 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0834_
timestamp 1
transform -1 0 26680 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0835_
timestamp 1
transform -1 0 23552 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0836_
timestamp 1
transform 1 0 14996 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0837_
timestamp 1
transform 1 0 15180 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0838_
timestamp 1
transform -1 0 15272 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0839_
timestamp 1
transform 1 0 16468 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0840_
timestamp 1
transform 1 0 16192 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0841_
timestamp 1
transform 1 0 17112 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0842_
timestamp 1
transform 1 0 16284 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0843_
timestamp 1
transform 1 0 14168 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0844_
timestamp 1
transform 1 0 15180 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1
transform 1 0 14260 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1
transform -1 0 15180 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0847_
timestamp 1
transform 1 0 20056 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0848_
timestamp 1
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0849_
timestamp 1
transform 1 0 19044 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0850_
timestamp 1
transform 1 0 20332 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0851_
timestamp 1
transform 1 0 19872 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0852_
timestamp 1
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1
transform -1 0 14352 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0854_
timestamp 1
transform 1 0 15180 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0855_
timestamp 1
transform 1 0 12972 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _0856_
timestamp 1
transform -1 0 12972 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0857_
timestamp 1
transform 1 0 19688 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0858_
timestamp 1
transform -1 0 22632 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0859_
timestamp 1
transform 1 0 21252 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0860_
timestamp 1
transform -1 0 23368 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0861_
timestamp 1
transform -1 0 23644 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0862_
timestamp 1
transform -1 0 27876 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0863_
timestamp 1
transform -1 0 28336 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0864_
timestamp 1
transform 1 0 23828 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0865_
timestamp 1
transform -1 0 27140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0866_
timestamp 1
transform -1 0 28336 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0867_
timestamp 1
transform 1 0 25300 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0868_
timestamp 1
transform -1 0 25484 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0869_
timestamp 1
transform 1 0 25576 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 1
transform 1 0 25944 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0871_
timestamp 1
transform 1 0 19136 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0872_
timestamp 1
transform -1 0 19688 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1
transform 1 0 17848 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0874_
timestamp 1
transform -1 0 24932 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0875_
timestamp 1
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0876_
timestamp 1
transform -1 0 26220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0877_
timestamp 1
transform -1 0 27232 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0878_
timestamp 1
transform 1 0 15364 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0879_
timestamp 1
transform -1 0 25576 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0880_
timestamp 1
transform 1 0 19412 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0881_
timestamp 1
transform 1 0 28888 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1
transform -1 0 30728 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0883_
timestamp 1
transform -1 0 30268 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0884_
timestamp 1
transform -1 0 29992 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1
transform 1 0 29256 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0886_
timestamp 1
transform 1 0 29532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0887_
timestamp 1
transform -1 0 18216 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0888_
timestamp 1
transform 1 0 19136 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0889_
timestamp 1
transform 1 0 17940 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0890_
timestamp 1
transform 1 0 18216 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0891_
timestamp 1
transform 1 0 18676 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0892_
timestamp 1
transform 1 0 20056 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0893_
timestamp 1
transform -1 0 19504 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0894_
timestamp 1
transform 1 0 15732 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0895_
timestamp 1
transform 1 0 17296 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0896_
timestamp 1
transform -1 0 19136 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0897_
timestamp 1
transform -1 0 19136 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0898_
timestamp 1
transform 1 0 17480 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0899_
timestamp 1
transform -1 0 16468 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0900_
timestamp 1
transform 1 0 16100 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _0901_
timestamp 1
transform -1 0 8464 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_2  _0902_
timestamp 1
transform -1 0 13156 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0903_
timestamp 1
transform -1 0 18216 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0904_
timestamp 1
transform 1 0 22448 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0905_
timestamp 1
transform -1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0906_
timestamp 1
transform 1 0 21344 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0907_
timestamp 1
transform 1 0 17664 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0908_
timestamp 1
transform -1 0 18584 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _0909_
timestamp 1
transform 1 0 17296 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1
transform 1 0 18676 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 1
transform 1 0 16284 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0912_
timestamp 1
transform -1 0 20884 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _0913_
timestamp 1
transform 1 0 21344 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0914_
timestamp 1
transform 1 0 20056 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0915_
timestamp 1
transform 1 0 17756 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0916_
timestamp 1
transform 1 0 18400 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_2  _0917_
timestamp 1
transform -1 0 12604 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _0918_
timestamp 1
transform -1 0 11592 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0919_
timestamp 1
transform -1 0 11960 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0920_
timestamp 1
transform -1 0 12512 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1
transform -1 0 12052 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0922_
timestamp 1
transform 1 0 11040 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0923_
timestamp 1
transform -1 0 13432 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0924_
timestamp 1
transform -1 0 12880 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0925_
timestamp 1
transform 1 0 11868 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1
transform -1 0 12788 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0927_
timestamp 1
transform 1 0 10396 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0928_
timestamp 1
transform 1 0 11224 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0929_
timestamp 1
transform -1 0 15180 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1
transform 1 0 13616 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0931_
timestamp 1
transform -1 0 11960 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0932_
timestamp 1
transform -1 0 12972 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0933_
timestamp 1
transform 1 0 10028 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0934_
timestamp 1
transform -1 0 12880 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0935_
timestamp 1
transform 1 0 11132 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0936_
timestamp 1
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1
transform -1 0 14812 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0938_
timestamp 1
transform 1 0 13524 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0939_
timestamp 1
transform 1 0 13524 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0940_
timestamp 1
transform -1 0 14536 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 1
transform -1 0 13524 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0942_
timestamp 1
transform 1 0 12880 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0944_
timestamp 1
transform 1 0 12604 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0945_
timestamp 1
transform 1 0 19228 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0946_
timestamp 1
transform -1 0 23000 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1
transform -1 0 23460 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0948_
timestamp 1
transform 1 0 22264 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0949_
timestamp 1
transform 1 0 22172 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0950_
timestamp 1
transform -1 0 28704 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0951_
timestamp 1
transform 1 0 28336 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0952_
timestamp 1
transform -1 0 24380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0953_
timestamp 1
transform -1 0 29716 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0954_
timestamp 1
transform 1 0 28796 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0955_
timestamp 1
transform 1 0 18676 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1
transform 1 0 18308 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0957_
timestamp 1
transform 1 0 30176 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1
transform 1 0 28428 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0959_
timestamp 1
transform -1 0 29348 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0960_
timestamp 1
transform -1 0 30176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0961_
timestamp 1
transform -1 0 14904 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _0962_
timestamp 1
transform -1 0 13984 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0964_
timestamp 1
transform 1 0 8372 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0965_
timestamp 1
transform -1 0 8004 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0966_
timestamp 1
transform 1 0 9200 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0967_
timestamp 1
transform -1 0 9384 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0968_
timestamp 1
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0969_
timestamp 1
transform 1 0 7820 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0970_
timestamp 1
transform 1 0 8464 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0971_
timestamp 1
transform 1 0 7820 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0972_
timestamp 1
transform -1 0 27416 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0973_
timestamp 1
transform 1 0 24932 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0974_
timestamp 1
transform -1 0 26220 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 1
transform 1 0 22724 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0976_
timestamp 1
transform -1 0 22724 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0977_
timestamp 1
transform -1 0 22172 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1
transform 1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0979_
timestamp 1
transform 1 0 20424 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0980_
timestamp 1
transform -1 0 19136 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0981_
timestamp 1
transform -1 0 18676 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0983_
timestamp 1
transform -1 0 17480 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 1
transform -1 0 16744 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0985_
timestamp 1
transform 1 0 15364 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0986_
timestamp 1
transform -1 0 16008 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0987_
timestamp 1
transform 1 0 16468 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0988_
timestamp 1
transform 1 0 17664 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 1
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0990_
timestamp 1
transform 1 0 18768 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0991_
timestamp 1
transform 1 0 19412 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0992_
timestamp 1
transform 1 0 21252 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0993_
timestamp 1
transform -1 0 24932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0994_
timestamp 1
transform 1 0 22724 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0995_
timestamp 1
transform 1 0 27784 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0996_
timestamp 1
transform -1 0 28520 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0997_
timestamp 1
transform 1 0 27232 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0998_
timestamp 1
transform -1 0 27048 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0999_
timestamp 1
transform -1 0 27232 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1000_
timestamp 1
transform 1 0 26312 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1001_
timestamp 1
transform -1 0 26404 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1002_
timestamp 1
transform -1 0 23920 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1003_
timestamp 1
transform -1 0 23552 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1
transform -1 0 24380 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1005_
timestamp 1
transform 1 0 22632 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1
transform -1 0 26128 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1007_
timestamp 1
transform 1 0 25300 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1
transform 1 0 27232 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1009_
timestamp 1
transform 1 0 26772 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1
transform -1 0 27876 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1011_
timestamp 1
transform 1 0 26404 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1
transform 1 0 27968 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1013_
timestamp 1
transform 1 0 27968 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1014_
timestamp 1
transform -1 0 28060 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1015_
timestamp 1
transform 1 0 28244 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1
transform 1 0 28060 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1017_
timestamp 1
transform 1 0 28520 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1
transform 1 0 29164 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1019_
timestamp 1
transform 1 0 28244 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1020_
timestamp 1
transform -1 0 13156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1021_
timestamp 1
transform -1 0 10028 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1022_
timestamp 1
transform -1 0 7636 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1023_
timestamp 1
transform -1 0 8280 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1024_
timestamp 1
transform -1 0 6348 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1025_
timestamp 1
transform -1 0 6256 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1026_
timestamp 1
transform -1 0 3864 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1027_
timestamp 1
transform -1 0 4968 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1028_
timestamp 1
transform -1 0 3128 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1029_
timestamp 1
transform -1 0 6992 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1
transform -1 0 14352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1031_
timestamp 1
transform 1 0 5152 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1032_
timestamp 1
transform -1 0 3680 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1033_
timestamp 1
transform -1 0 4508 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1034_
timestamp 1
transform -1 0 3036 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1035_
timestamp 1
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1036_
timestamp 1
transform -1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1037_
timestamp 1
transform -1 0 2024 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1038_
timestamp 1
transform 1 0 4048 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1039_
timestamp 1
transform -1 0 4600 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1040_
timestamp 1
transform -1 0 3128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1041_
timestamp 1
transform -1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1042_
timestamp 1
transform -1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1
transform 1 0 2116 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1044_
timestamp 1
transform -1 0 6624 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1045_
timestamp 1
transform -1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1046_
timestamp 1
transform -1 0 6164 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1047_
timestamp 1
transform 1 0 5428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1048_
timestamp 1
transform -1 0 7176 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1
transform -1 0 6992 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1050_
timestamp 1
transform -1 0 8924 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1051_
timestamp 1
transform 1 0 8280 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1052_
timestamp 1
transform 1 0 11408 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1053_
timestamp 1
transform -1 0 9292 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1054_
timestamp 1
transform 1 0 10948 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1055_
timestamp 1
transform 1 0 9568 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1056_
timestamp 1
transform 1 0 13524 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 1
transform 1 0 12420 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1058_
timestamp 1
transform -1 0 15180 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1059_
timestamp 1
transform -1 0 12696 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1060_
timestamp 1
transform 1 0 12052 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1061_
timestamp 1
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1062_
timestamp 1
transform 1 0 18400 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1063_
timestamp 1
transform -1 0 21896 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1064_
timestamp 1
transform -1 0 21344 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1
transform 1 0 19872 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1066_
timestamp 1
transform 1 0 4508 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1067_
timestamp 1
transform -1 0 4324 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1
transform -1 0 6900 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1069_
timestamp 1
transform 1 0 4232 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1070_
timestamp 1
transform -1 0 6440 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1071_
timestamp 1
transform 1 0 5060 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1072_
timestamp 1
transform 1 0 13616 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1073_
timestamp 1
transform -1 0 14536 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1074_
timestamp 1
transform 1 0 9476 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1075_
timestamp 1
transform -1 0 10672 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1
transform 1 0 13156 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1077_
timestamp 1
transform -1 0 14352 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1
transform -1 0 13708 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1
transform -1 0 13432 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1080_
timestamp 1
transform 1 0 18768 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1081_
timestamp 1
transform -1 0 19596 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1082_
timestamp 1
transform 1 0 26036 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1083_
timestamp 1
transform -1 0 27140 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1084_
timestamp 1
transform 1 0 29072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1085_
timestamp 1
transform -1 0 29348 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1086_
timestamp 1
transform 1 0 14444 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1087_
timestamp 1
transform -1 0 14904 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1088_
timestamp 1
transform -1 0 10856 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1089_
timestamp 1
transform 1 0 11132 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1090_
timestamp 1
transform 1 0 10212 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1091_
timestamp 1
transform 1 0 10120 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1092_
timestamp 1
transform 1 0 7084 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1093_
timestamp 1
transform -1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1094_
timestamp 1
transform 1 0 9108 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp 1
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1
transform 1 0 10856 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1097_
timestamp 1
transform -1 0 12052 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1
transform 1 0 7820 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1
transform -1 0 9936 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1
transform 1 0 8740 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1
transform 1 0 7084 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1103_
timestamp 1
transform 1 0 7544 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1
transform -1 0 9568 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1105_
timestamp 1
transform 1 0 8372 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1
transform 1 0 12512 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1107_
timestamp 1
transform -1 0 12512 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1108_
timestamp 1
transform 1 0 10948 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1109_
timestamp 1
transform 1 0 11224 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1110_
timestamp 1
transform 1 0 8556 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1111_
timestamp 1
transform 1 0 9016 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1
transform -1 0 10396 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1113_
timestamp 1
transform 1 0 9016 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1114_
timestamp 1
transform 1 0 11776 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1115_
timestamp 1
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1
transform 1 0 11408 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1
transform 1 0 12604 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1
transform 1 0 13432 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1119_
timestamp 1
transform 1 0 11868 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1120_
timestamp 1
transform -1 0 8648 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1
transform 1 0 10304 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1
transform -1 0 11408 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1
transform 1 0 9844 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1124_
timestamp 1
transform 1 0 3128 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1125_
timestamp 1
transform 1 0 3588 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1126_
timestamp 1
transform -1 0 3956 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1127_
timestamp 1
transform -1 0 4048 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1128_
timestamp 1
transform -1 0 4508 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _1129_
timestamp 1
transform 1 0 2944 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1130_
timestamp 1
transform -1 0 4416 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 1
transform -1 0 3128 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1132_
timestamp 1
transform -1 0 4508 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1133_
timestamp 1
transform -1 0 3680 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1134_
timestamp 1
transform 1 0 4600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1135_
timestamp 1
transform 1 0 3772 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1136_
timestamp 1
transform 1 0 3404 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1137_
timestamp 1
transform -1 0 2944 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1138_
timestamp 1
transform 1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1139_
timestamp 1
transform -1 0 2392 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1140_
timestamp 1
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1141_
timestamp 1
transform -1 0 2484 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1142_
timestamp 1
transform 1 0 3864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp 1
transform -1 0 3496 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1144_
timestamp 1
transform -1 0 2576 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1145_
timestamp 1
transform 1 0 3680 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1146_
timestamp 1
transform -1 0 3128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1147_
timestamp 1
transform -1 0 16376 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1148_
timestamp 1
transform 1 0 17204 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1149_
timestamp 1
transform -1 0 9568 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1150_
timestamp 1
transform -1 0 28520 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1151_
timestamp 1
transform 1 0 17848 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1152_
timestamp 1
transform 1 0 8924 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1153_
timestamp 1
transform 1 0 19044 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1154_
timestamp 1
transform -1 0 19964 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1155_
timestamp 1
transform 1 0 15180 0 1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__o22ai_1  _1156_
timestamp 1
transform 1 0 17756 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _1157_
timestamp 1
transform 1 0 17388 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1158_
timestamp 1
transform 1 0 17112 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1159_
timestamp 1
transform 1 0 15180 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1160_
timestamp 1
transform 1 0 16100 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1161_
timestamp 1
transform 1 0 15364 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1
transform 1 0 16652 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _1163_
timestamp 1
transform -1 0 17204 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1164_
timestamp 1
transform -1 0 17112 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1165_
timestamp 1
transform -1 0 16008 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1166_
timestamp 1
transform -1 0 16928 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1167_
timestamp 1
transform -1 0 16652 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1
transform -1 0 16836 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1169_
timestamp 1
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1170_
timestamp 1
transform 1 0 16468 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1171_
timestamp 1
transform 1 0 13984 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1172_
timestamp 1
transform -1 0 15088 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1173_
timestamp 1
transform 1 0 14352 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1174_
timestamp 1
transform -1 0 13432 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1175_
timestamp 1
transform -1 0 13984 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1176_
timestamp 1
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1177_
timestamp 1
transform 1 0 14076 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1178_
timestamp 1
transform 1 0 13708 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1179_
timestamp 1
transform 1 0 13524 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1
transform 1 0 12144 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1181_
timestamp 1
transform 1 0 6808 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1182_
timestamp 1
transform 1 0 2300 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1183_
timestamp 1
transform 1 0 7176 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1184_
timestamp 1
transform 1 0 5888 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1
transform 1 0 5796 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1186_
timestamp 1
transform -1 0 6624 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1
transform 1 0 6532 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1188_
timestamp 1
transform 1 0 6992 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1
transform 1 0 5244 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1190_
timestamp 1
transform -1 0 6532 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1191_
timestamp 1
transform -1 0 6164 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1192_
timestamp 1
transform -1 0 4692 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1
transform -1 0 3956 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1
transform 1 0 3956 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1195_
timestamp 1
transform 1 0 4692 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1196_
timestamp 1
transform -1 0 3404 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1197_
timestamp 1
transform 1 0 2024 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1198_
timestamp 1
transform 1 0 2484 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1199_
timestamp 1
transform -1 0 3036 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1200_
timestamp 1
transform 1 0 2300 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1201_
timestamp 1
transform -1 0 15548 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1
transform -1 0 5704 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1203_
timestamp 1
transform 1 0 4508 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1204_
timestamp 1
transform -1 0 5428 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1205_
timestamp 1
transform 1 0 3864 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1206_
timestamp 1
transform 1 0 3956 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1207_
timestamp 1
transform -1 0 4692 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1208_
timestamp 1
transform 1 0 5060 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1209_
timestamp 1
transform 1 0 4692 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1210_
timestamp 1
transform -1 0 6256 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1211_
timestamp 1
transform 1 0 5244 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1212_
timestamp 1
transform 1 0 5796 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1213_
timestamp 1
transform -1 0 6256 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1214_
timestamp 1
transform 1 0 5152 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1215_
timestamp 1
transform 1 0 5796 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1216_
timestamp 1
transform -1 0 6256 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1217_
timestamp 1
transform 1 0 4508 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1218_
timestamp 1
transform 1 0 6256 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1219_
timestamp 1
transform -1 0 5704 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1220_
timestamp 1
transform -1 0 5428 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1221_
timestamp 1
transform -1 0 5520 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1222_
timestamp 1
transform 1 0 10580 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1223_
timestamp 1
transform -1 0 10764 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1224_
timestamp 1
transform 1 0 11408 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1225_
timestamp 1
transform 1 0 5796 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1226_
timestamp 1
transform -1 0 6072 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1227_
timestamp 1
transform 1 0 4600 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1228_
timestamp 1
transform 1 0 3956 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1229_
timestamp 1
transform 1 0 2392 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1230_
timestamp 1
transform 1 0 5060 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1231_
timestamp 1
transform 1 0 6072 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1232_
timestamp 1
transform 1 0 4232 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1
transform 1 0 2116 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1234_
timestamp 1
transform -1 0 5612 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 1
transform 1 0 6532 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1236_
timestamp 1
transform -1 0 5520 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1237_
timestamp 1
transform 1 0 4508 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1238_
timestamp 1
transform 1 0 3036 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1239_
timestamp 1
transform 1 0 4048 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1240_
timestamp 1
transform 1 0 3312 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1241_
timestamp 1
transform -1 0 4048 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1242_
timestamp 1
transform -1 0 7268 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1243_
timestamp 1
transform -1 0 26128 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1244_
timestamp 1
transform -1 0 19228 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1245_
timestamp 1
transform 1 0 21436 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1246_
timestamp 1
transform -1 0 22908 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1247_
timestamp 1
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1248_
timestamp 1
transform -1 0 19228 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1249_
timestamp 1
transform 1 0 15456 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1250_
timestamp 1
transform 1 0 16008 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1251_
timestamp 1
transform -1 0 17664 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1252_
timestamp 1
transform 1 0 9476 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1253_
timestamp 1
transform 1 0 10948 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1254_
timestamp 1
transform -1 0 10120 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1255_
timestamp 1
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1256_
timestamp 1
transform -1 0 10856 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__or3b_1  _1257_
timestamp 1
transform 1 0 10120 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1258_
timestamp 1
transform -1 0 8648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1259_
timestamp 1
transform 1 0 9108 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1261_
timestamp 1
transform -1 0 25576 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1262_
timestamp 1
transform -1 0 27048 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1263_
timestamp 1
transform 1 0 25576 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1264_
timestamp 1
transform 1 0 29900 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1265_
timestamp 1
transform -1 0 29532 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1266_
timestamp 1
transform 1 0 27416 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1267_
timestamp 1
transform -1 0 26128 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1268_
timestamp 1
transform 1 0 18676 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1269_
timestamp 1
transform 1 0 19044 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1270_
timestamp 1
transform -1 0 19688 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1271_
timestamp 1
transform -1 0 19044 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1272_
timestamp 1
transform -1 0 19320 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1273_
timestamp 1
transform -1 0 20240 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1
transform 1 0 17480 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1275_
timestamp 1
transform 1 0 20516 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1276_
timestamp 1
transform -1 0 22448 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1277_
timestamp 1
transform -1 0 23736 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1278_
timestamp 1
transform 1 0 22724 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1279_
timestamp 1
transform -1 0 24288 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1280_
timestamp 1
transform 1 0 23828 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1281_
timestamp 1
transform 1 0 23000 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1282_
timestamp 1
transform 1 0 25668 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1283_
timestamp 1
transform 1 0 25392 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1284_
timestamp 1
transform 1 0 25300 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1285_
timestamp 1
transform 1 0 25024 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1286_
timestamp 1
transform -1 0 25392 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1287_
timestamp 1
transform -1 0 27784 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1288_
timestamp 1
transform 1 0 26864 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1289_
timestamp 1
transform 1 0 26496 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1290_
timestamp 1
transform -1 0 27140 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1291_
timestamp 1
transform -1 0 27416 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1292_
timestamp 1
transform 1 0 27508 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1293_
timestamp 1
transform -1 0 30636 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1294_
timestamp 1
transform -1 0 29900 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1295_
timestamp 1
transform 1 0 29992 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1296_
timestamp 1
transform -1 0 29624 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1297_
timestamp 1
transform 1 0 27784 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1298_
timestamp 1
transform -1 0 29716 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1299_
timestamp 1
transform -1 0 29992 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1300_
timestamp 1
transform -1 0 31280 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1301_
timestamp 1
transform -1 0 28888 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1302_
timestamp 1
transform 1 0 27784 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1303_
timestamp 1
transform -1 0 30452 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1304_
timestamp 1
transform 1 0 29900 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1305_
timestamp 1
transform 1 0 28244 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1306_
timestamp 1
transform -1 0 28428 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1307_
timestamp 1
transform 1 0 27968 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1308_
timestamp 1
transform 1 0 28336 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1309_
timestamp 1
transform 1 0 28980 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1310_
timestamp 1
transform -1 0 28152 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1
transform -1 0 29716 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1
transform 1 0 27784 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1313_
timestamp 1
transform -1 0 30820 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1314_
timestamp 1
transform -1 0 30084 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1315_
timestamp 1
transform -1 0 31096 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1316_
timestamp 1
transform 1 0 29808 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1317_
timestamp 1
transform 1 0 28428 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1318_
timestamp 1
transform -1 0 29072 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1319_
timestamp 1
transform 1 0 28980 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1320_
timestamp 1
transform -1 0 28888 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1321_
timestamp 1
transform -1 0 29348 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1
transform -1 0 27508 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1
transform -1 0 26220 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1324_
timestamp 1
transform -1 0 25760 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1325_
timestamp 1
transform 1 0 27416 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1326_
timestamp 1
transform 1 0 26220 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1327_
timestamp 1
transform 1 0 24012 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1328_
timestamp 1
transform 1 0 27232 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1329_
timestamp 1
transform -1 0 25668 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1330_
timestamp 1
transform 1 0 25668 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1331_
timestamp 1
transform 1 0 24012 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1
transform 1 0 23368 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1333_
timestamp 1
transform -1 0 24564 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1334_
timestamp 1
transform -1 0 25300 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1335_
timestamp 1
transform 1 0 25300 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1336_
timestamp 1
transform -1 0 24932 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1
transform 1 0 20700 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1338_
timestamp 1
transform -1 0 23828 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1339_
timestamp 1
transform -1 0 23092 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1340_
timestamp 1
transform 1 0 22724 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1341_
timestamp 1
transform -1 0 23000 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1
transform -1 0 21988 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1343_
timestamp 1
transform -1 0 21712 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1344_
timestamp 1
transform 1 0 21712 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1345_
timestamp 1
transform -1 0 21160 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 1
transform 1 0 15548 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1347_
timestamp 1
transform -1 0 16100 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _1348_
timestamp 1
transform -1 0 19688 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1349_
timestamp 1
transform -1 0 19136 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1350_
timestamp 1
transform 1 0 18400 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1351_
timestamp 1
transform -1 0 17572 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1352_
timestamp 1
transform -1 0 18952 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 1
transform 1 0 18492 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1
transform -1 0 18584 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1355_
timestamp 1
transform 1 0 21344 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1356_
timestamp 1
transform 1 0 22908 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1357_
timestamp 1
transform 1 0 21252 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1
transform -1 0 21160 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1359_
timestamp 1
transform 1 0 21988 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1360_
timestamp 1
transform -1 0 21160 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1361_
timestamp 1
transform -1 0 22172 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1362_
timestamp 1
transform -1 0 25944 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1363_
timestamp 1
transform -1 0 9108 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1364_
timestamp 1
transform 1 0 9936 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1365_
timestamp 1
transform 1 0 5796 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1366_
timestamp 1
transform -1 0 6808 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1367__3
timestamp 1
transform -1 0 11316 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1368__4
timestamp 1
transform -1 0 21620 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1369__5
timestamp 1
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1370__6
timestamp 1
transform 1 0 19596 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1371__7
timestamp 1
transform -1 0 17204 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1372__8
timestamp 1
transform -1 0 16744 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1373__9
timestamp 1
transform 1 0 19964 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1374__10
timestamp 1
transform 1 0 23828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1375__11
timestamp 1
transform -1 0 26312 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1376__12
timestamp 1
transform 1 0 23460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1377__13
timestamp 1
transform -1 0 26772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1378__14
timestamp 1
transform 1 0 28612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1379__15
timestamp 1
transform 1 0 28980 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1380__16
timestamp 1
transform 1 0 31096 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1381__17
timestamp 1
transform -1 0 30084 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1382__18
timestamp 1
transform 1 0 28980 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1383__19
timestamp 1
transform 1 0 28612 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1384__20
timestamp 1
transform -1 0 28060 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1385__21
timestamp 1
transform -1 0 25208 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1386__22
timestamp 1
transform -1 0 24288 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1387__23
timestamp 1
transform 1 0 17112 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1388__24
timestamp 1
transform 1 0 8648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1389__25
timestamp 1
transform -1 0 14996 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1390__26
timestamp 1
transform 1 0 5152 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1391__27
timestamp 1
transform 1 0 1288 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1392__28
timestamp 1
transform -1 0 1932 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1393__29
timestamp 1
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1394__30
timestamp 1
transform -1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1395__31
timestamp 1
transform 1 0 1288 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1396__32
timestamp 1
transform -1 0 2300 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1397__33
timestamp 1
transform -1 0 4232 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1398__34
timestamp 1
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1399__35
timestamp 1
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1400__36
timestamp 1
transform 1 0 1288 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1401__37
timestamp 1
transform 1 0 7176 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1402__38
timestamp 1
transform 1 0 11868 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1403__39
timestamp 1
transform -1 0 12972 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1404__40
timestamp 1
transform 1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1405__41
timestamp 1
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1406__42
timestamp 1
transform -1 0 2668 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1407__43
timestamp 1
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1408__44
timestamp 1
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1409__45
timestamp 1
transform -1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1410__46
timestamp 1
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1411__47
timestamp 1
transform -1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1412__48
timestamp 1
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1413__49
timestamp 1
transform -1 0 6072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1414__50
timestamp 1
transform 1 0 8464 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1415__51
timestamp 1
transform 1 0 8004 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1416__52
timestamp 1
transform -1 0 12880 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1417__53
timestamp 1
transform -1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1418__54
timestamp 1
transform 1 0 12972 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1419__55
timestamp 1
transform -1 0 9016 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1420__56
timestamp 1
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1421__57
timestamp 1
transform -1 0 12236 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1422__58
timestamp 1
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1423__59
timestamp 1
transform -1 0 7084 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1424__60
timestamp 1
transform -1 0 10304 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1425__61
timestamp 1
transform -1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1426__62
timestamp 1
transform -1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1427__63
timestamp 1
transform -1 0 8740 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1428__64
timestamp 1
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1429__65
timestamp 1
transform -1 0 10120 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1430__66
timestamp 1
transform -1 0 16376 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1431__67
timestamp 1
transform -1 0 29716 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1432__68
timestamp 1
transform -1 0 28704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1433__69
timestamp 1
transform -1 0 19872 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1434__70
timestamp 1
transform -1 0 14076 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1435__71
timestamp 1
transform -1 0 14444 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1436__72
timestamp 1
transform -1 0 11316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1437__73
timestamp 1
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1438__74
timestamp 1
transform 1 0 22356 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1439__75
timestamp 1
transform -1 0 14628 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1440__76
timestamp 1
transform 1 0 12052 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1441__77
timestamp 1
transform -1 0 13432 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1442__78
timestamp 1
transform -1 0 12052 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1443__79
timestamp 1
transform 1 0 9016 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1444__80
timestamp 1
transform 1 0 8924 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1445__81
timestamp 1
transform -1 0 7268 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1446__82
timestamp 1
transform -1 0 4600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1447__83
timestamp 1
transform 1 0 4600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1448__84
timestamp 1
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1449__85
timestamp 1
transform -1 0 2116 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1450__86
timestamp 1
transform -1 0 5244 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1451__87
timestamp 1
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1452__88
timestamp 1
transform 1 0 3220 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1453__89
timestamp 1
transform -1 0 4232 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1454__90
timestamp 1
transform 1 0 2024 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1455__91
timestamp 1
transform -1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1456__92
timestamp 1
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1457__93
timestamp 1
transform -1 0 29348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1458__94
timestamp 1
transform 1 0 28612 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1459__95
timestamp 1
transform -1 0 26772 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1460__96
timestamp 1
transform -1 0 28152 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1461__97
timestamp 1
transform 1 0 25208 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1462__98
timestamp 1
transform -1 0 22816 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1463__99
timestamp 1
transform 1 0 24932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1464__100
timestamp 1
transform 1 0 24380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1465__101
timestamp 1
transform 1 0 20516 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1466__102
timestamp 1
transform -1 0 20424 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1467__103
timestamp 1
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1468__104
timestamp 1
transform -1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1469__105
timestamp 1
transform 1 0 16192 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1470__106
timestamp 1
transform 1 0 14996 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1471__107
timestamp 1
transform 1 0 9936 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1472__108
timestamp 1
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1473__109
timestamp 1
transform -1 0 8188 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1474__110
timestamp 1
transform 1 0 6532 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1475__111
timestamp 1
transform 1 0 30728 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1476__112
timestamp 1
transform 1 0 28060 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1477__113
timestamp 1
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1478__114
timestamp 1
transform -1 0 29624 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1479__115
timestamp 1
transform -1 0 24656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1480__116
timestamp 1
transform 1 0 28152 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1481__117
timestamp 1
transform 1 0 21988 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1482__118
timestamp 1
transform -1 0 23736 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1483__119
timestamp 1
transform -1 0 13800 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1484__120
timestamp 1
transform 1 0 13156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1485__121
timestamp 1
transform -1 0 10488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1486__122
timestamp 1
transform 1 0 10580 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1487__123
timestamp 1
transform -1 0 13800 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1488__124
timestamp 1
transform -1 0 11224 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1489__125
timestamp 1
transform -1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1490__126
timestamp 1
transform -1 0 10028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1491__127
timestamp 1
transform 1 0 17020 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1492__128
timestamp 1
transform 1 0 14996 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1493__129
timestamp 1
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1494__130
timestamp 1
transform -1 0 26772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1495__131
timestamp 1
transform 1 0 24656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1496__132
timestamp 1
transform -1 0 28612 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1497__133
timestamp 1
transform -1 0 25668 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1498__134
timestamp 1
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1499__135
timestamp 1
transform 1 0 23828 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1500__136
timestamp 1
transform -1 0 22080 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1501__137
timestamp 1
transform 1 0 13340 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1502__138
timestamp 1
transform 1 0 13616 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1503__139
timestamp 1
transform 1 0 20332 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1504__140
timestamp 1
transform 1 0 18768 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1505__141
timestamp 1
transform -1 0 21252 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1506__142
timestamp 1
transform -1 0 17112 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1507__143
timestamp 1
transform 1 0 16192 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1508__144
timestamp 1
transform 1 0 14444 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1509_
timestamp 1
transform 1 0 5612 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1510_
timestamp 1
transform -1 0 11040 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1511_
timestamp 1
transform 1 0 21252 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1512_
timestamp 1
transform 1 0 21160 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1513_
timestamp 1
transform -1 0 20424 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1514_
timestamp 1
transform 1 0 16836 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1515_
timestamp 1
transform 1 0 16100 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1516_
timestamp 1
transform 1 0 21252 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1517_
timestamp 1
transform -1 0 23644 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1518_
timestamp 1
transform -1 0 26036 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1519_
timestamp 1
transform 1 0 23828 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1520_
timestamp 1
transform 1 0 26404 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1521_
timestamp 1
transform 1 0 29256 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1522_
timestamp 1
transform 1 0 29348 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1
transform -1 0 30544 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1
transform -1 0 29900 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1
transform 1 0 29348 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1
transform 1 0 29256 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1
transform 1 0 27324 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1
transform 1 0 24840 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1
transform 1 0 23828 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1530_
timestamp 1
transform 1 0 17204 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1
transform 1 0 9108 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1
transform 1 0 14628 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1
transform -1 0 22724 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1534_
timestamp 1
transform 1 0 28980 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1535_
timestamp 1
transform 1 0 28428 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1536_
timestamp 1
transform 1 0 26956 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1537_
timestamp 1
transform 1 0 28980 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1538_
timestamp 1
transform 1 0 25852 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1539_
timestamp 1
transform 1 0 24656 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1540_
timestamp 1
transform 1 0 24380 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1541_
timestamp 1
transform 1 0 23644 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1542_
timestamp 1
transform 1 0 5796 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1543_
timestamp 1
transform 1 0 1564 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1544_
timestamp 1
transform 1 0 1564 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1545_
timestamp 1
transform 1 0 1656 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1546_
timestamp 1
transform 1 0 1380 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1547_
timestamp 1
transform 1 0 1564 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1548_
timestamp 1
transform 1 0 1932 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1549_
timestamp 1
transform 1 0 3220 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1550_
timestamp 1
transform 1 0 5612 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1551_
timestamp 1
transform 1 0 5796 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1552_
timestamp 1
transform 1 0 1472 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1553_
timestamp 1
transform -1 0 7176 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1554_
timestamp 1
transform 1 0 12236 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1555_
timestamp 1
transform 1 0 12604 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1556_
timestamp 1
transform 1 0 14720 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1557_
timestamp 1
transform 1 0 14904 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1558_
timestamp 1
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1559_
timestamp 1
transform 1 0 1656 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1560_
timestamp 1
transform 1 0 1656 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1561_
timestamp 1
transform 1 0 1840 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1562_
timestamp 1
transform 1 0 1656 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1563_
timestamp 1
transform 1 0 1932 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1564_
timestamp 1
transform 1 0 3588 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1565_
timestamp 1
transform -1 0 5888 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1566_
timestamp 1
transform 1 0 8648 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1567_
timestamp 1
transform 1 0 8372 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1568_
timestamp 1
transform 1 0 11960 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1569_
timestamp 1
transform -1 0 13248 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1570_
timestamp 1
transform -1 0 13708 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1571_
timestamp 1
transform 1 0 9200 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1572_
timestamp 1
transform 1 0 8740 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1573_
timestamp 1
transform -1 0 11224 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1574_
timestamp 1
transform 1 0 8188 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1575_
timestamp 1
transform 1 0 6716 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1576_
timestamp 1
transform -1 0 10028 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1577_
timestamp 1
transform -1 0 8832 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1578_
timestamp 1
transform -1 0 12788 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1579_
timestamp 1
transform 1 0 8372 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1580_
timestamp 1
transform 1 0 7636 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1
transform 1 0 10120 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1
transform -1 0 16008 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1
transform 1 0 29348 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1
transform -1 0 28060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1
transform 1 0 19228 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1
transform 1 0 13708 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1
transform 1 0 14076 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1
transform 1 0 10948 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1
transform 1 0 14076 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1
transform -1 0 22356 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1
transform 1 0 14076 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1
transform 1 0 12604 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1
transform 1 0 12880 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1
transform -1 0 11408 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1
transform 1 0 9292 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1
transform -1 0 9844 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1
transform 1 0 6164 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1
transform 1 0 4232 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1
transform 1 0 4876 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1
transform 1 0 1656 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1
transform 1 0 1748 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1
transform 1 0 1656 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1
transform 1 0 3496 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1
transform 1 0 3680 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1
transform 1 0 3404 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1607_
timestamp 1
transform -1 0 30544 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1
transform -1 0 30268 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1
transform 1 0 28980 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1
transform 1 0 28980 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1
transform 1 0 26404 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1
transform 1 0 27508 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1
transform -1 0 26312 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1
transform 1 0 23276 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1
transform -1 0 25300 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1
transform -1 0 23736 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1
transform 1 0 20792 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1618_
timestamp 1
transform 1 0 19596 0 -1 1632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1
transform 1 0 19320 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1
transform 1 0 17112 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1
transform 1 0 16192 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1
transform 1 0 15272 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1623_
timestamp 1
transform -1 0 9936 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1
transform -1 0 8740 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1
transform 1 0 7820 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1
transform -1 0 30820 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1
transform 1 0 28704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1
transform 1 0 18676 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1
transform 1 0 29256 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1
transform 1 0 23828 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1
transform 1 0 28980 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1
transform 1 0 22264 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1
transform 1 0 22908 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1
transform 1 0 12880 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1
transform 1 0 13524 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1
transform 1 0 10488 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1
transform 1 0 13156 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1
transform 1 0 10948 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1
transform 1 0 11500 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1
transform 1 0 10580 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1
transform 1 0 17756 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1
transform 1 0 15272 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1
transform 1 0 18860 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1
transform 1 0 26404 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1
transform 1 0 24932 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1
transform -1 0 27876 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1
transform 1 0 23644 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1
transform -1 0 27968 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1
transform -1 0 23552 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1
transform 1 0 21712 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1
transform 1 0 13432 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1
transform 1 0 13708 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1
transform 1 0 20608 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1
transform 1 0 19504 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1
transform 1 0 19688 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1
transform 1 0 16744 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1
transform 1 0 16100 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1
transform 1 0 14720 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1667_
timestamp 1
transform 1 0 9568 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1668_
timestamp 1
transform 1 0 8740 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1669_
timestamp 1
transform 1 0 8372 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1670_
timestamp 1
transform -1 0 8188 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1671_
timestamp 1
transform -1 0 6348 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1672_
timestamp 1
transform 1 0 8004 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1673_
timestamp 1
transform 1 0 7452 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1674_
timestamp 1
transform 1 0 11132 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1675_
timestamp 1
transform -1 0 10580 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1676_
timestamp 1
transform -1 0 16008 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 17940 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1
transform -1 0 7176 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1
transform 1 0 6256 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1
transform -1 0 13432 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1
transform 1 0 5796 0 -1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1
transform -1 0 6716 0 1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1
transform -1 0 12788 0 -1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1
transform 1 0 12788 0 -1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1
transform 1 0 21252 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1
transform 1 0 21252 0 -1 9248
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1
transform 1 0 26404 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1
transform 1 0 26496 0 1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1
transform 1 0 19872 0 1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1
transform -1 0 22264 0 -1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1
transform 1 0 26036 0 1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1
transform 1 0 26404 0 -1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_6  clkload0
timestamp 1
transform -1 0 7820 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  clkload1
timestamp 1
transform 1 0 12604 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  clkload2
timestamp 1
transform 1 0 12604 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_8  clkload3
timestamp 1
transform -1 0 5704 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  clkload4
timestamp 1
transform 1 0 4416 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_8  clkload5
timestamp 1
transform 1 0 11776 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_4  clkload6
timestamp 1
transform 1 0 11132 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  clkload7
timestamp 1
transform 1 0 20792 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_8  clkload8
timestamp 1
transform 1 0 20332 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload9
timestamp 1
transform -1 0 26312 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  clkload10
timestamp 1
transform -1 0 27968 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  clkload11
timestamp 1
transform 1 0 19688 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_12  clkload12
timestamp 1
transform 1 0 21068 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  clkload13
timestamp 1
transform 1 0 26404 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_16  clkload14
timestamp 1
transform -1 0 27232 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1
transform -1 0 17112 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout12
timestamp 1
transform 1 0 23828 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 1
transform 1 0 21988 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1
transform 1 0 22724 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout16
timestamp 1
transform -1 0 14444 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1
transform -1 0 5060 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 1
transform 1 0 24288 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1
transform 1 0 24288 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1
transform -1 0 24012 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1
transform -1 0 17296 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1
transform 1 0 23920 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1
transform 1 0 18216 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1
transform 1 0 22356 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1
transform -1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1
transform -1 0 17756 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1
transform 1 0 20148 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1
transform 1 0 28060 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1
transform 1 0 16284 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1
transform 1 0 15548 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1
transform 1 0 17112 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1
transform -1 0 10764 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1
transform -1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1
transform 1 0 16100 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1
transform -1 0 14904 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout40
timestamp 1
transform 1 0 16744 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1
transform -1 0 19688 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1
transform -1 0 19688 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1
transform -1 0 20516 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1
transform 1 0 27140 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1
transform -1 0 16652 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1
transform -1 0 26772 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1
transform 1 0 13800 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1
transform 1 0 14904 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 1
transform -1 0 14444 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1
transform 1 0 2760 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 1
transform -1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 1
transform 1 0 15456 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 1
transform -1 0 10028 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 1
transform -1 0 11592 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 1
transform 1 0 16652 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 1
transform -1 0 15640 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp 1
transform -1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp 1
transform -1 0 26312 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 1
transform 1 0 27692 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1
transform 1 0 30820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp 1
transform -1 0 22172 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp 1
transform -1 0 29900 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp 1
transform -1 0 30268 0 -1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1
transform 1 0 5796 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_65
timestamp 1
transform 1 0 6532 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77
timestamp 1
transform 1 0 7636 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1
transform 1 0 8188 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_94
timestamp 1636968456
transform 1 0 9200 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_106
timestamp 1
transform 1 0 10304 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636968456
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636968456
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_202
timestamp 1
transform 1 0 19136 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_220
timestamp 1
transform 1 0 20792 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636968456
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636968456
transform 1 0 30084 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333
timestamp 1
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_39
timestamp 1
transform 1 0 4140 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_91
timestamp 1
transform 1 0 8924 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1
transform 1 0 16100 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_194
timestamp 1
transform 1 0 18400 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_205
timestamp 1
transform 1 0 19412 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_237
timestamp 1
transform 1 0 22356 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_263
timestamp 1
transform 1 0 24748 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_288
timestamp 1
transform 1 0 27048 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_292
timestamp 1
transform 1 0 27416 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_309
timestamp 1636968456
transform 1 0 28980 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_321
timestamp 1636968456
transform 1 0 30084 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_333
timestamp 1
transform 1 0 31188 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_71
timestamp 1
transform 1 0 7084 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1
transform 1 0 8096 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_101
timestamp 1
transform 1 0 9844 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_159
timestamp 1
transform 1 0 15180 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_219
timestamp 1
transform 1 0 20700 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_228
timestamp 1
transform 1 0 21528 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_236
timestamp 1
transform 1 0 22264 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1
transform 1 0 23552 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_300
timestamp 1
transform 1 0 28152 0 1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636968456
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636968456
transform 1 0 30084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 1
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_27
timestamp 1
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_33
timestamp 1636968456
transform 1 0 3588 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_45
timestamp 1
transform 1 0 4692 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1
transform 1 0 5796 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_71
timestamp 1
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_94
timestamp 1
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_120
timestamp 1
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_128
timestamp 1
transform 1 0 12328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_153
timestamp 1
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_160
timestamp 1
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 1
transform 1 0 16100 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_197
timestamp 1
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_201
timestamp 1
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_208
timestamp 1636968456
transform 1 0 19688 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_220
timestamp 1
transform 1 0 20792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_248
timestamp 1
transform 1 0 23368 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_271
timestamp 1
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 1
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_281
timestamp 1
transform 1 0 26404 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_297
timestamp 1636968456
transform 1 0 27876 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_309
timestamp 1636968456
transform 1 0 28980 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_321
timestamp 1636968456
transform 1 0 30084 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_333
timestamp 1
transform 1 0 31188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3
timestamp 1
transform 1 0 828 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 1
transform 1 0 3220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_45
timestamp 1
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_49
timestamp 1
transform 1 0 5060 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_53
timestamp 1
transform 1 0 5428 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_66
timestamp 1
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_73
timestamp 1
transform 1 0 7268 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_89
timestamp 1
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_116
timestamp 1636968456
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_128
timestamp 1
transform 1 0 12328 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_132
timestamp 1
transform 1 0 12696 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_151
timestamp 1636968456
transform 1 0 14444 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_163
timestamp 1636968456
transform 1 0 15548 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_175
timestamp 1636968456
transform 1 0 16652 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_187
timestamp 1
transform 1 0 17756 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_200
timestamp 1636968456
transform 1 0 18952 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_212
timestamp 1
transform 1 0 20056 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_216
timestamp 1
transform 1 0 20424 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_256
timestamp 1636968456
transform 1 0 24104 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_268
timestamp 1636968456
transform 1 0 25208 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_295
timestamp 1
transform 1 0 27692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_325
timestamp 1
transform 1 0 30452 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_333
timestamp 1
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1
transform 1 0 828 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_11
timestamp 1
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_29
timestamp 1
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_36
timestamp 1
transform 1 0 3864 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636968456
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636968456
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_93
timestamp 1
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_97
timestamp 1
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636968456
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1636968456
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_137
timestamp 1
transform 1 0 13156 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_145
timestamp 1
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_150
timestamp 1636968456
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_162
timestamp 1
transform 1 0 15456 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_175
timestamp 1636968456
transform 1 0 16652 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_187
timestamp 1
transform 1 0 17756 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_197
timestamp 1636968456
transform 1 0 18676 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_209
timestamp 1636968456
transform 1 0 19780 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_221
timestamp 1
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_225
timestamp 1
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_244
timestamp 1636968456
transform 1 0 23000 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_256
timestamp 1
transform 1 0 24104 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_264
timestamp 1
transform 1 0 24840 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 1
transform 1 0 26404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_288
timestamp 1
transform 1 0 27048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_296
timestamp 1
transform 1 0 27784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_303
timestamp 1
transform 1 0 28428 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_309
timestamp 1
transform 1 0 28980 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_313
timestamp 1636968456
transform 1 0 29348 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_325
timestamp 1
transform 1 0 30452 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_333
timestamp 1
transform 1 0 31188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1
transform 1 0 828 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_11
timestamp 1
transform 1 0 1564 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_44
timestamp 1
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_69
timestamp 1
transform 1 0 6900 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_77
timestamp 1
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_103
timestamp 1
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_124
timestamp 1636968456
transform 1 0 11960 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_136
timestamp 1
transform 1 0 13064 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_205
timestamp 1636968456
transform 1 0 19412 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_217
timestamp 1636968456
transform 1 0 20516 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_229
timestamp 1
transform 1 0 21620 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_233
timestamp 1
transform 1 0 21988 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_241
timestamp 1
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_256
timestamp 1636968456
transform 1 0 24104 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_268
timestamp 1636968456
transform 1 0 25208 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_280
timestamp 1
transform 1 0 26312 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_288
timestamp 1
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_295
timestamp 1
transform 1 0 27692 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_325
timestamp 1
transform 1 0 30452 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 1
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1
transform 1 0 828 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_11
timestamp 1
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636968456
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_69
timestamp 1
transform 1 0 6900 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_77
timestamp 1
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_95
timestamp 1636968456
transform 1 0 9292 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_107
timestamp 1
transform 1 0 10396 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_155
timestamp 1
transform 1 0 14812 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_159
timestamp 1
transform 1 0 15180 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_176
timestamp 1
transform 1 0 16744 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_191
timestamp 1
transform 1 0 18124 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_213
timestamp 1
transform 1 0 20148 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp 1
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_225
timestamp 1
transform 1 0 21252 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_233
timestamp 1
transform 1 0 21988 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_247
timestamp 1
transform 1 0 23276 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_257
timestamp 1
transform 1 0 24196 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_263
timestamp 1
transform 1 0 24748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 1
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_292
timestamp 1
transform 1 0 27416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_304
timestamp 1
transform 1 0 28520 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_323
timestamp 1636968456
transform 1 0 30268 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 1
transform 1 0 828 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_68
timestamp 1636968456
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_96
timestamp 1636968456
transform 1 0 9384 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_108
timestamp 1
transform 1 0 10488 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_112
timestamp 1
transform 1 0 10856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_133
timestamp 1
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_152
timestamp 1636968456
transform 1 0 14536 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_164
timestamp 1
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_172
timestamp 1636968456
transform 1 0 16376 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_184
timestamp 1636968456
transform 1 0 17480 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_200
timestamp 1636968456
transform 1 0 18952 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_212
timestamp 1
transform 1 0 20056 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_220
timestamp 1
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_234
timestamp 1
transform 1 0 22080 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_238
timestamp 1
transform 1 0 22448 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_279
timestamp 1636968456
transform 1 0 26220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_291
timestamp 1
transform 1 0 27324 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_295
timestamp 1
transform 1 0 27692 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_332
timestamp 1
transform 1 0 31096 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_15
timestamp 1
transform 1 0 1932 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_70
timestamp 1
transform 1 0 6992 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_78
timestamp 1
transform 1 0 7728 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_84
timestamp 1
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_102
timestamp 1
transform 1 0 9936 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_120
timestamp 1
transform 1 0 11592 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_128
timestamp 1
transform 1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_144
timestamp 1636968456
transform 1 0 13800 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_156
timestamp 1636968456
transform 1 0 14904 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636968456
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1636968456
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_193
timestamp 1
transform 1 0 18308 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_209
timestamp 1636968456
transform 1 0 19780 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_262
timestamp 1
transform 1 0 24656 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_268
timestamp 1
transform 1 0 25208 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_272
timestamp 1
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636968456
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_293
timestamp 1
transform 1 0 27508 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_316
timestamp 1636968456
transform 1 0 29624 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_328
timestamp 1
transform 1 0 30728 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_334
timestamp 1
transform 1 0 31280 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636968456
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_48
timestamp 1636968456
transform 1 0 4968 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_60
timestamp 1
transform 1 0 6072 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_105
timestamp 1636968456
transform 1 0 10212 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_117
timestamp 1
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_124
timestamp 1
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_146
timestamp 1636968456
transform 1 0 13984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_158
timestamp 1
transform 1 0 15088 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_166
timestamp 1
transform 1 0 15824 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_174
timestamp 1
transform 1 0 16560 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_185
timestamp 1
transform 1 0 17572 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_219
timestamp 1636968456
transform 1 0 20700 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_249
timestamp 1
transform 1 0 23460 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_256
timestamp 1636968456
transform 1 0 24104 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_268
timestamp 1
transform 1 0 25208 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_276
timestamp 1
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1636968456
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_309
timestamp 1
transform 1 0 28980 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_323
timestamp 1636968456
transform 1 0 30268 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636968456
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636968456
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_27
timestamp 1
transform 1 0 3036 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_40
timestamp 1
transform 1 0 4232 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 1
transform 1 0 5060 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_61
timestamp 1
transform 1 0 6164 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_97
timestamp 1
transform 1 0 9476 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_105
timestamp 1
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_129
timestamp 1
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_156
timestamp 1
transform 1 0 14904 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_160
timestamp 1
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1636968456
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_181
timestamp 1
transform 1 0 17204 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_193
timestamp 1
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_211
timestamp 1
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_219
timestamp 1
transform 1 0 20700 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_236
timestamp 1
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_263
timestamp 1
transform 1 0 24748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_272
timestamp 1
transform 1 0 25576 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1636968456
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_305
timestamp 1
transform 1 0 28612 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_328
timestamp 1
transform 1 0 30728 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_334
timestamp 1
transform 1 0 31280 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636968456
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636968456
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636968456
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636968456
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1636968456
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_96
timestamp 1
transform 1 0 9384 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_167
timestamp 1636968456
transform 1 0 15916 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_179
timestamp 1
transform 1 0 17020 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_203
timestamp 1
transform 1 0 19228 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_211
timestamp 1
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_236
timestamp 1636968456
transform 1 0 22264 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_248
timestamp 1
transform 1 0 23368 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1
transform 1 0 23828 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_257
timestamp 1
transform 1 0 24196 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_268
timestamp 1
transform 1 0 25208 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_290
timestamp 1
transform 1 0 27232 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_298
timestamp 1
transform 1 0 27968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_325
timestamp 1
transform 1 0 30452 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 1
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636968456
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_27
timestamp 1
transform 1 0 3036 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 1
transform 1 0 5060 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1636968456
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_69
timestamp 1
transform 1 0 6900 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_75
timestamp 1
transform 1 0 7452 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_84
timestamp 1636968456
transform 1 0 8280 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_96
timestamp 1
transform 1 0 9384 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_100
timestamp 1
transform 1 0 9752 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_104
timestamp 1
transform 1 0 10120 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_108
timestamp 1
transform 1 0 10488 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_130
timestamp 1
transform 1 0 12512 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_136
timestamp 1
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_158
timestamp 1
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_175
timestamp 1
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_194
timestamp 1
transform 1 0 18400 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_205
timestamp 1
transform 1 0 19412 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_213
timestamp 1
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_236
timestamp 1
transform 1 0 22264 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_259
timestamp 1636968456
transform 1 0 24380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_271
timestamp 1
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_292
timestamp 1
transform 1 0 27416 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_330
timestamp 1
transform 1 0 30912 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_334
timestamp 1
transform 1 0 31280 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_15
timestamp 1
transform 1 0 1932 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_21
timestamp 1
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_34
timestamp 1
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_66
timestamp 1636968456
transform 1 0 6624 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp 1
transform 1 0 7728 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_89
timestamp 1636968456
transform 1 0 8740 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_101
timestamp 1636968456
transform 1 0 9844 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_113
timestamp 1636968456
transform 1 0 10948 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_125
timestamp 1636968456
transform 1 0 12052 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_144
timestamp 1
transform 1 0 13800 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_150
timestamp 1
transform 1 0 14352 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_170
timestamp 1
transform 1 0 16192 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_192
timestamp 1
transform 1 0 18216 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_213
timestamp 1
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_234
timestamp 1
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1636968456
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_265
timestamp 1
transform 1 0 24932 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_271
timestamp 1
transform 1 0 25484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_278
timestamp 1
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_298
timestamp 1
transform 1 0 27968 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_317
timestamp 1636968456
transform 1 0 29716 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_329
timestamp 1
transform 1 0 30820 0 1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_38
timestamp 1
transform 1 0 4048 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_63
timestamp 1
transform 1 0 6348 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_71
timestamp 1
transform 1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_98
timestamp 1636968456
transform 1 0 9568 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp 1
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_140
timestamp 1636968456
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_152
timestamp 1
transform 1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_164
timestamp 1
transform 1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_169
timestamp 1
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_177
timestamp 1
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_183
timestamp 1
transform 1 0 17388 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_191
timestamp 1
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_203
timestamp 1
transform 1 0 19228 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_209
timestamp 1
transform 1 0 19780 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_244
timestamp 1
transform 1 0 23000 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_250
timestamp 1
transform 1 0 23552 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_262
timestamp 1636968456
transform 1 0 24656 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_274
timestamp 1
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_281
timestamp 1
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_298
timestamp 1
transform 1 0 27968 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_306
timestamp 1
transform 1 0 28704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_328
timestamp 1
transform 1 0 30728 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_334
timestamp 1
transform 1 0 31280 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_3
timestamp 1
transform 1 0 828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_69
timestamp 1
transform 1 0 6900 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_134
timestamp 1
transform 1 0 12880 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1
transform 1 0 13524 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_148
timestamp 1
transform 1 0 14168 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_159
timestamp 1
transform 1 0 15180 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_167
timestamp 1
transform 1 0 15916 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_174
timestamp 1636968456
transform 1 0 16560 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_186
timestamp 1
transform 1 0 17664 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_197
timestamp 1
transform 1 0 18676 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_208
timestamp 1
transform 1 0 19688 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_220
timestamp 1636968456
transform 1 0 20792 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_232
timestamp 1
transform 1 0 21896 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_277
timestamp 1
transform 1 0 26036 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_309
timestamp 1
transform 1 0 28980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_316
timestamp 1
transform 1 0 29624 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_322
timestamp 1636968456
transform 1 0 30176 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_334
timestamp 1
transform 1 0 31280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1
transform 1 0 828 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_11
timestamp 1
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_20
timestamp 1
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_26
timestamp 1
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_47
timestamp 1
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_64
timestamp 1
transform 1 0 6440 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_72
timestamp 1
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_98
timestamp 1
transform 1 0 9568 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1
transform 1 0 10948 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1636968456
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_153
timestamp 1
transform 1 0 14628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1
transform 1 0 16100 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_186
timestamp 1636968456
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_198
timestamp 1
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_206
timestamp 1
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_233
timestamp 1
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_240
timestamp 1
transform 1 0 22632 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_248
timestamp 1
transform 1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_267
timestamp 1
transform 1 0 25116 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_275
timestamp 1
transform 1 0 25852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_302
timestamp 1
transform 1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1
transform 1 0 30820 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636968456
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_15
timestamp 1
transform 1 0 1932 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_21
timestamp 1
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_32
timestamp 1
transform 1 0 3496 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_40
timestamp 1
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_45
timestamp 1
transform 1 0 4692 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_53
timestamp 1
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_62
timestamp 1636968456
transform 1 0 6256 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_74
timestamp 1
transform 1 0 7360 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_78
timestamp 1
transform 1 0 7728 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_96
timestamp 1
transform 1 0 9384 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_104
timestamp 1
transform 1 0 10120 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_110
timestamp 1
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_136
timestamp 1
transform 1 0 13064 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_144
timestamp 1
transform 1 0 13800 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_185
timestamp 1
transform 1 0 17572 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_197
timestamp 1
transform 1 0 18676 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_225
timestamp 1636968456
transform 1 0 21252 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_237
timestamp 1636968456
transform 1 0 22356 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1
transform 1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_261
timestamp 1
transform 1 0 24564 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_273
timestamp 1
transform 1 0 25668 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_288
timestamp 1636968456
transform 1 0 27048 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_300
timestamp 1
transform 1 0 28152 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_309
timestamp 1
transform 1 0 28980 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_313
timestamp 1
transform 1 0 29348 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_322
timestamp 1
transform 1 0 30176 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_331
timestamp 1
transform 1 0 31004 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1
transform 1 0 828 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_11
timestamp 1
transform 1 0 1564 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_43
timestamp 1
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_48
timestamp 1
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_64
timestamp 1636968456
transform 1 0 6440 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_76
timestamp 1636968456
transform 1 0 7544 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_88
timestamp 1
transform 1 0 8648 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_102
timestamp 1
transform 1 0 9936 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636968456
transform 1 0 10948 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636968456
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1636968456
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1636968456
transform 1 0 14260 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_161
timestamp 1
transform 1 0 15364 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1
transform 1 0 16100 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_175
timestamp 1636968456
transform 1 0 16652 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_187
timestamp 1636968456
transform 1 0 17756 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_199
timestamp 1
transform 1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 1
transform 1 0 20608 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_225
timestamp 1
transform 1 0 21252 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_250
timestamp 1636968456
transform 1 0 23552 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_262
timestamp 1
transform 1 0 24656 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_268
timestamp 1
transform 1 0 25208 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_297
timestamp 1
transform 1 0 27876 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1
transform 1 0 30820 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 1
transform 1 0 828 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_32
timestamp 1
transform 1 0 3496 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_59
timestamp 1636968456
transform 1 0 5980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_71
timestamp 1
transform 1 0 7084 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_75
timestamp 1
transform 1 0 7452 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_106
timestamp 1
transform 1 0 10304 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_114
timestamp 1
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_124
timestamp 1
transform 1 0 11960 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_130
timestamp 1
transform 1 0 12512 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1636968456
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_153
timestamp 1
transform 1 0 14628 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_159
timestamp 1
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_189
timestamp 1
transform 1 0 17940 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_197
timestamp 1
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_219
timestamp 1
transform 1 0 20700 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_256
timestamp 1
transform 1 0 24104 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_281
timestamp 1
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 1
transform 1 0 28704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_309
timestamp 1
transform 1 0 28980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_313
timestamp 1
transform 1 0 29348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_317
timestamp 1
transform 1 0 29716 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_327
timestamp 1
transform 1 0 30636 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636968456
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_22
timestamp 1
transform 1 0 2576 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_40
timestamp 1
transform 1 0 4232 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_48
timestamp 1
transform 1 0 4968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_62
timestamp 1
transform 1 0 6256 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_66
timestamp 1
transform 1 0 6624 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_103
timestamp 1
transform 1 0 10028 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_120
timestamp 1
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_144
timestamp 1
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_156
timestamp 1
transform 1 0 14904 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_185
timestamp 1
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1
transform 1 0 20516 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_225
timestamp 1
transform 1 0 21252 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_231
timestamp 1
transform 1 0 21804 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_248
timestamp 1636968456
transform 1 0 23368 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_260
timestamp 1
transform 1 0 24472 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_271
timestamp 1
transform 1 0 25484 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_299
timestamp 1636968456
transform 1 0 28060 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_311
timestamp 1
transform 1 0 29164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1
transform 1 0 30820 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 1
transform 1 0 828 0 1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_45
timestamp 1636968456
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_57
timestamp 1
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_65
timestamp 1
transform 1 0 6532 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_93
timestamp 1
transform 1 0 9108 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_105
timestamp 1
transform 1 0 10212 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_113
timestamp 1
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_120
timestamp 1
transform 1 0 11592 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_124
timestamp 1
transform 1 0 11960 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_128
timestamp 1
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 1
transform 1 0 12972 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_146
timestamp 1
transform 1 0 13984 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_173
timestamp 1
transform 1 0 16468 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_202
timestamp 1636968456
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_214
timestamp 1636968456
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_226
timestamp 1636968456
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_238
timestamp 1636968456
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1
transform 1 0 23552 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1636968456
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_265
timestamp 1
transform 1 0 24932 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_273
timestamp 1
transform 1 0 25668 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_285
timestamp 1636968456
transform 1 0 26772 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_297
timestamp 1
transform 1 0 27876 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_328
timestamp 1
transform 1 0 30728 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_334
timestamp 1
transform 1 0 31280 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636968456
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_15
timestamp 1
transform 1 0 1932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_42
timestamp 1
transform 1 0 4416 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_50
timestamp 1
transform 1 0 5152 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_74
timestamp 1
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_83
timestamp 1
transform 1 0 8188 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_87
timestamp 1
transform 1 0 8556 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_98
timestamp 1
transform 1 0 9568 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_129
timestamp 1
transform 1 0 12420 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_154
timestamp 1
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_158
timestamp 1
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_162
timestamp 1
transform 1 0 15456 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1
transform 1 0 16100 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_176
timestamp 1
transform 1 0 16744 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_182
timestamp 1
transform 1 0 17296 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_200
timestamp 1636968456
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_212
timestamp 1636968456
transform 1 0 20056 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_233
timestamp 1636968456
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_245
timestamp 1
transform 1 0 23092 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1
transform 1 0 26128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_281
timestamp 1
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_289
timestamp 1
transform 1 0 27140 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_307
timestamp 1
transform 1 0 28796 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_316
timestamp 1
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_333
timestamp 1
transform 1 0 31188 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636968456
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_15
timestamp 1
transform 1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_19
timestamp 1
transform 1 0 2300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_23
timestamp 1
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 1
transform 1 0 3220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_42
timestamp 1
transform 1 0 4416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_53
timestamp 1
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636968456
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_111
timestamp 1
transform 1 0 10764 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_117
timestamp 1636968456
transform 1 0 11316 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_129
timestamp 1
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_147
timestamp 1
transform 1 0 14076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_155
timestamp 1
transform 1 0 14812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_163
timestamp 1
transform 1 0 15548 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_174
timestamp 1
transform 1 0 16560 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1636968456
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_209
timestamp 1
transform 1 0 19780 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_240
timestamp 1
transform 1 0 22632 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_278
timestamp 1
transform 1 0 26128 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_292
timestamp 1
transform 1 0 27416 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1
transform 1 0 28704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_309
timestamp 1
transform 1 0 28980 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_327
timestamp 1
transform 1 0 30636 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1
transform 1 0 828 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_9
timestamp 1
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_31
timestamp 1636968456
transform 1 0 3404 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_43
timestamp 1
transform 1 0 4508 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_67
timestamp 1
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_86
timestamp 1
transform 1 0 8464 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_121
timestamp 1
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_133
timestamp 1
transform 1 0 12788 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_137
timestamp 1
transform 1 0 13156 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_169
timestamp 1
transform 1 0 16100 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_175
timestamp 1
transform 1 0 16652 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_179
timestamp 1
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_192
timestamp 1
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_199
timestamp 1
transform 1 0 18860 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_207
timestamp 1
transform 1 0 19596 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_281
timestamp 1
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_299
timestamp 1
transform 1 0 28060 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_308
timestamp 1
transform 1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_334
timestamp 1
transform 1 0 31280 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1
transform 1 0 828 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_7
timestamp 1
transform 1 0 1196 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_53
timestamp 1
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_75
timestamp 1
transform 1 0 7452 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 1
transform 1 0 8372 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_127
timestamp 1
transform 1 0 12236 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_131
timestamp 1
transform 1 0 12604 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1
transform 1 0 13524 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_167
timestamp 1
transform 1 0 15916 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_180
timestamp 1
transform 1 0 17112 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_205
timestamp 1
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_217
timestamp 1
transform 1 0 20516 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_231
timestamp 1636968456
transform 1 0 21804 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_243
timestamp 1
transform 1 0 22908 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_260
timestamp 1
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_294
timestamp 1
transform 1 0 27600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_325
timestamp 1
transform 1 0 30452 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_333
timestamp 1
transform 1 0 31188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1
transform 1 0 828 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_7
timestamp 1
transform 1 0 1196 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_36
timestamp 1
transform 1 0 3864 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_77
timestamp 1636968456
transform 1 0 7636 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_121
timestamp 1
transform 1 0 11684 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_143
timestamp 1
transform 1 0 13708 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_159
timestamp 1
transform 1 0 15180 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_169
timestamp 1
transform 1 0 16100 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_214
timestamp 1
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1636968456
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_249
timestamp 1
transform 1 0 23460 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_253
timestamp 1
transform 1 0 23828 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_262
timestamp 1
transform 1 0 24656 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_268
timestamp 1636968456
transform 1 0 25208 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1636968456
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_293
timestamp 1
transform 1 0 27508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_328
timestamp 1
transform 1 0 30728 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_334
timestamp 1
transform 1 0 31280 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1
transform 1 0 828 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_29
timestamp 1
transform 1 0 3220 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_37
timestamp 1
transform 1 0 3956 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_75
timestamp 1
transform 1 0 7452 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_100
timestamp 1
transform 1 0 9752 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_111
timestamp 1
transform 1 0 10764 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_149
timestamp 1636968456
transform 1 0 14260 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_161
timestamp 1636968456
transform 1 0 15364 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_173
timestamp 1
transform 1 0 16468 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_179
timestamp 1
transform 1 0 17020 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_276
timestamp 1
transform 1 0 25944 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1636968456
transform 1 0 30084 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_333
timestamp 1
transform 1 0 31188 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1636968456
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_15
timestamp 1
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_41
timestamp 1
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1636968456
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_81
timestamp 1
transform 1 0 8004 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_89
timestamp 1
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_121
timestamp 1
transform 1 0 11684 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_144
timestamp 1
transform 1 0 13800 0 -1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_172
timestamp 1636968456
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_201
timestamp 1
transform 1 0 19044 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_294
timestamp 1
transform 1 0 27600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_301
timestamp 1
transform 1 0 28244 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_326
timestamp 1
transform 1 0 30544 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_334
timestamp 1
transform 1 0 31280 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_3
timestamp 1
transform 1 0 828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_25
timestamp 1
transform 1 0 2852 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1
transform 1 0 3220 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_39
timestamp 1
transform 1 0 4140 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_66
timestamp 1636968456
transform 1 0 6624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_78
timestamp 1
transform 1 0 7728 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_120
timestamp 1
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_179
timestamp 1
transform 1 0 17020 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_187
timestamp 1
transform 1 0 17756 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_193
timestamp 1
transform 1 0 18308 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_208
timestamp 1
transform 1 0 19688 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_256
timestamp 1
transform 1 0 24104 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636968456
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_15
timestamp 1
transform 1 0 1932 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_19
timestamp 1
transform 1 0 2300 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_73
timestamp 1
transform 1 0 7268 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_81
timestamp 1
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_122
timestamp 1
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_145
timestamp 1
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_180
timestamp 1636968456
transform 1 0 17112 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_192
timestamp 1
transform 1 0 18216 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_198
timestamp 1
transform 1 0 18768 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_210
timestamp 1
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_218
timestamp 1
transform 1 0 20608 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_253
timestamp 1
transform 1 0 23828 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_263
timestamp 1
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_299
timestamp 1
transform 1 0 28060 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_310
timestamp 1
transform 1 0 29072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1
transform 1 0 30820 0 -1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1636968456
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_15
timestamp 1
transform 1 0 1932 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_23
timestamp 1
transform 1 0 2668 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_29
timestamp 1
transform 1 0 3220 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_68
timestamp 1636968456
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_80
timestamp 1
transform 1 0 7912 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_85
timestamp 1
transform 1 0 8372 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_120
timestamp 1
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_130
timestamp 1
transform 1 0 12512 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_149
timestamp 1
transform 1 0 14260 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_155
timestamp 1
transform 1 0 14812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_160
timestamp 1
transform 1 0 15272 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_182
timestamp 1636968456
transform 1 0 17296 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_197
timestamp 1
transform 1 0 18676 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_201
timestamp 1
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_219
timestamp 1
transform 1 0 20700 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_244
timestamp 1
transform 1 0 23000 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_248
timestamp 1
transform 1 0 23368 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_269
timestamp 1
transform 1 0 25300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_287
timestamp 1
transform 1 0 26956 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_295
timestamp 1
transform 1 0 27692 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_326
timestamp 1
transform 1 0 30544 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_334
timestamp 1
transform 1 0 31280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1
transform 1 0 828 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_35
timestamp 1
transform 1 0 3772 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_61
timestamp 1636968456
transform 1 0 6164 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_73
timestamp 1636968456
transform 1 0 7268 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_85
timestamp 1
transform 1 0 8372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1
transform 1 0 10764 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_134
timestamp 1636968456
transform 1 0 12880 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_146
timestamp 1
transform 1 0 13984 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_154
timestamp 1
transform 1 0 14720 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_158
timestamp 1
transform 1 0 15088 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_162
timestamp 1
transform 1 0 15456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_177
timestamp 1636968456
transform 1 0 16836 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_189
timestamp 1
transform 1 0 17940 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_200
timestamp 1
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_208
timestamp 1636968456
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 1
transform 1 0 20792 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_241
timestamp 1636968456
transform 1 0 22724 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_253
timestamp 1
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_276
timestamp 1
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_297
timestamp 1
transform 1 0 27876 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_333
timestamp 1
transform 1 0 31188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_3
timestamp 1
transform 1 0 828 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_11
timestamp 1
transform 1 0 1564 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_15
timestamp 1
transform 1 0 1932 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_45
timestamp 1636968456
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_57
timestamp 1636968456
transform 1 0 5796 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_69
timestamp 1
transform 1 0 6900 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_81
timestamp 1
transform 1 0 8004 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_113
timestamp 1636968456
transform 1 0 10948 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_125
timestamp 1636968456
transform 1 0 12052 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1
transform 1 0 13156 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_141
timestamp 1
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_152
timestamp 1
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_182
timestamp 1
transform 1 0 17296 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_216
timestamp 1
transform 1 0 20424 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_224
timestamp 1
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_229
timestamp 1636968456
transform 1 0 21620 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_241
timestamp 1
transform 1 0 22724 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1
transform 1 0 23460 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_253
timestamp 1
transform 1 0 23828 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_260
timestamp 1636968456
transform 1 0 24472 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_272
timestamp 1
transform 1 0 25576 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_278
timestamp 1
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_285
timestamp 1636968456
transform 1 0 26772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_304
timestamp 1
transform 1 0 28520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_328
timestamp 1
transform 1 0 30728 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_334
timestamp 1
transform 1 0 31280 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1636968456
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_15
timestamp 1
transform 1 0 1932 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_31
timestamp 1
transform 1 0 3404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_38
timestamp 1
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_42
timestamp 1
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_49
timestamp 1
transform 1 0 5060 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_67
timestamp 1636968456
transform 1 0 6716 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_79
timestamp 1636968456
transform 1 0 7820 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_91
timestamp 1
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1
transform 1 0 10580 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_121
timestamp 1
transform 1 0 11684 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_146
timestamp 1
transform 1 0 13984 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_159
timestamp 1
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_178
timestamp 1636968456
transform 1 0 16928 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_190
timestamp 1
transform 1 0 18032 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_194
timestamp 1
transform 1 0 18400 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_210
timestamp 1
transform 1 0 19872 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_218
timestamp 1
transform 1 0 20608 0 -1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_239
timestamp 1636968456
transform 1 0 22540 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_251
timestamp 1636968456
transform 1 0 23644 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_263
timestamp 1
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1
transform 1 0 26220 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_288
timestamp 1
transform 1 0 27048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_301
timestamp 1
transform 1 0 28244 0 -1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_323
timestamp 1636968456
transform 1 0 30268 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_3
timestamp 1
transform 1 0 828 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_7
timestamp 1
transform 1 0 1196 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_45
timestamp 1
transform 1 0 4692 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_54
timestamp 1
transform 1 0 5520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_85
timestamp 1
transform 1 0 8372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_117
timestamp 1
transform 1 0 11316 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_158
timestamp 1
transform 1 0 15088 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_185
timestamp 1
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_192
timestamp 1
transform 1 0 18216 0 1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_202
timestamp 1636968456
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_214
timestamp 1
transform 1 0 20240 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_249
timestamp 1
transform 1 0 23460 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_253
timestamp 1
transform 1 0 23828 0 1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_291
timestamp 1636968456
transform 1 0 27324 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_303
timestamp 1
transform 1 0 28428 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1
transform 1 0 28796 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_325
timestamp 1
transform 1 0 30452 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_333
timestamp 1
transform 1 0 31188 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1636968456
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_40
timestamp 1
transform 1 0 4232 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_44
timestamp 1
transform 1 0 4600 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_48
timestamp 1
transform 1 0 4968 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_73
timestamp 1
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_102
timestamp 1
transform 1 0 9936 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1
transform 1 0 10580 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 1
transform 1 0 10948 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_121
timestamp 1
transform 1 0 11684 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_129
timestamp 1
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_159
timestamp 1
transform 1 0 15180 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1
transform 1 0 15916 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_169
timestamp 1
transform 1 0 16100 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_211
timestamp 1
transform 1 0 19964 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_219
timestamp 1
transform 1 0 20700 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_244
timestamp 1
transform 1 0 23000 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_250
timestamp 1
transform 1 0 23552 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_270
timestamp 1
transform 1 0 25392 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_274
timestamp 1
transform 1 0 25760 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 1
transform 1 0 26404 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_324
timestamp 1
transform 1 0 30360 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_332
timestamp 1
transform 1 0 31096 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636968456
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_15
timestamp 1
transform 1 0 1932 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_19
timestamp 1
transform 1 0 2300 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_23
timestamp 1
transform 1 0 2668 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1636968456
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_41
timestamp 1
transform 1 0 4324 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_49
timestamp 1
transform 1 0 5060 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 1
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_91
timestamp 1636968456
transform 1 0 8924 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_103
timestamp 1
transform 1 0 10028 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_111
timestamp 1
transform 1 0 10764 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_113
timestamp 1
transform 1 0 10948 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_124
timestamp 1
transform 1 0 11960 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_130
timestamp 1
transform 1 0 12512 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_150
timestamp 1636968456
transform 1 0 14352 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_162
timestamp 1
transform 1 0 15456 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_169
timestamp 1
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_177
timestamp 1
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_181
timestamp 1
transform 1 0 17204 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_187
timestamp 1
transform 1 0 17756 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1
transform 1 0 18308 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1636968456
transform 1 0 18676 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1636968456
transform 1 0 19780 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_221
timestamp 1
transform 1 0 20884 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_225
timestamp 1
transform 1 0 21252 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_229
timestamp 1
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_238
timestamp 1636968456
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1
transform 1 0 23552 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_256
timestamp 1
transform 1 0 24104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_278
timestamp 1
transform 1 0 26128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_287
timestamp 1
transform 1 0 26956 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_292
timestamp 1
transform 1 0 27416 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_298
timestamp 1
transform 1 0 27968 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_304
timestamp 1
transform 1 0 28520 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_325
timestamp 1
transform 1 0 30452 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_333
timestamp 1
transform 1 0 31188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 6532 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 3220 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform 1 0 6716 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 5060 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 3956 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 26036 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 8096 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 11684 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 6624 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform 1 0 4140 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 7820 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 3864 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 2300 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 6348 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 10764 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 17296 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 8004 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 21988 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 4600 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 3956 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 25392 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 19412 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 3864 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 30636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform 1 0 4876 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 7084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 14812 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform 1 0 12696 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 4048 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 25024 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 4692 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform -1 0 3864 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 10212 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 17480 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 22724 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 5520 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 26864 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 28888 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform -1 0 31188 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform -1 0 10764 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 28704 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform 1 0 10120 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 30452 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform 1 0 10948 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 21528 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform 1 0 11040 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 11684 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform -1 0 12512 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 30452 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 8280 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform -1 0 3588 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform -1 0 8188 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform -1 0 9476 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 28520 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 27968 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 27416 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 26956 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 26680 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 25760 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform 1 0 25116 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 24656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform -1 0 24104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform -1 0 22448 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_64
timestamp 1
transform -1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_65
timestamp 1
transform -1 0 8280 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_66
timestamp 1
transform -1 0 8924 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_67
timestamp 1
transform -1 0 13248 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_68
timestamp 1
transform -1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_jimktrains_vslc_69
timestamp 1
transform -1 0 11960 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire17
timestamp 1
transform -1 0 9384 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire18
timestamp 1
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  wire19
timestamp 1
transform 1 0 20332 0 1 11424
box -38 -48 406 592
<< labels >>
flabel metal4 s 4316 496 4636 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12090 496 12410 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19864 496 20184 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27638 496 27958 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11430 496 11750 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19204 496 19524 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26978 496 27298 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 29318 22104 29378 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 28214 22104 28274 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 27662 22104 27722 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 27110 22104 27170 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 26006 22104 26066 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 25454 22104 25514 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 24902 22104 24962 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 23798 22104 23858 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 23246 22104 23306 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 22694 22104 22754 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 21590 22104 21650 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 21038 22104 21098 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 20486 22104 20546 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 19382 22104 19442 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 9998 22104 10058 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal4 s 9446 22104 9506 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal4 s 8342 22104 8402 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal4 s 7790 22104 7850 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal4 s 7238 22104 7298 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal4 s 6134 22104 6194 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal4 s 14414 22104 14474 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal output
flabel metal4 s 13862 22104 13922 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal output
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal output
flabel metal4 s 12758 22104 12818 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal output
flabel metal4 s 12206 22104 12266 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal output
flabel metal4 s 11654 22104 11714 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal output
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal output
flabel metal4 s 10550 22104 10610 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal output
flabel metal4 s 18830 22104 18890 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal output
flabel metal4 s 18278 22104 18338 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal output
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal output
flabel metal4 s 17174 22104 17234 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal output
flabel metal4 s 16622 22104 16682 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal output
flabel metal4 s 16070 22104 16130 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal output
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal output
flabel metal4 s 14966 22104 15026 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
