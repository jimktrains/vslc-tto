`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave or surfer.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  tt_um_jimktrains_vslc user_project (

`ifdef GL_TEST
   .VPWR(VPWR),
   .VGND(VGND),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

`ifdef GL_TEST
  wire [7:0]stack = {
    // user_project.\core.exec.stack[15] ,
    // user_project.\core.exec.stack[14] ,
    // user_project.\core.exec.stack[13] ,
    // user_project.\core.exec.stack[12] ,
    // user_project.\core.exec.stack[11] ,
    // user_project.\core.exec.stack[10] ,
    // user_project.\core.exec.stack[9] ,
    // user_project.\core.exec.stack[8] ,
    user_project.\core.exec.stack[7] ,
    user_project.\core.exec.stack[6] ,
    user_project.\core.exec.stack[5] ,
    user_project.\core.exec.stack[4] ,
    user_project.\core.exec.stack[3] ,
    user_project.\core.exec.hos ,
    user_project.\core.exec.nos ,
    user_project.\core.exec.stack[0]
  };
`endif
`ifndef GL_TEST
  wire [7:0]stack = user_project.core.exec.stack ;
`endif
  wire tos = stack[0];


endmodule
